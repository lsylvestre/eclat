-- code generated from the following source code:
--   ../ocaml-vm/vm/mlvalue.ecl
--   ../ocaml-vm/vm/fail.ecl
--   ../ocaml-vm/vm/ram.ecl
--   ../ocaml-vm/vm/runtime.ecl
--   ../ocaml-vm/vm/debug.ecl
--   ../ocaml-vm/vm/alloc.ecl
--   ../ocaml-vm/vm/prims.ecl
--   ../ocaml-vm/bytecode.ecl
--   ../ocaml-vm/vm/vm.ecl
--   ../ocaml-vm/vm/target-specific/intel-max10/IOs.ecl
--   ../ocaml-vm/vm/target-specific/intel-max10/main.ecl
--
-- with the following command:
--
--    ./eclat -arg ((true,true,true,true,true,true,true,true,true,true),(true,false)) ../ocaml-vm/vm/mlvalue.ecl ../ocaml-vm/vm/fail.ecl ../ocaml-vm/vm/ram.ecl ../ocaml-vm/vm/runtime.ecl ../ocaml-vm/vm/debug.ecl ../ocaml-vm/vm/alloc.ecl ../ocaml-vm/vm/prims.ecl ../ocaml-vm/bytecode.ecl ../ocaml-vm/vm/vm.ecl ../ocaml-vm/vm/target-specific/intel-max10/IOs.ecl ../ocaml-vm/vm/target-specific/intel-max10/main.ecl

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.runtime.all;


entity main is
  
  port(signal clk    : in std_logic;
       signal reset  : in std_logic;
       signal run    : in std_logic;
       signal rdy    : out value(0 to 0);
       signal argument : in value(0 to 11);
       signal result : out value(0 to 57));
       
end entity;
architecture rtl of main is

  type t_state is (compute2134);
  signal state: t_state;
  type t_state_var3002 is (compute2140, pause_setI2141, pause_setI2142, pause_setI2143, pause_setI2144, pause_setI2145, pause_setI2146, pause_setI2147, pause_setI2148, pause_setI2149, pause_setI2150, pause_setI2151, pause_setI2152, pause_setI2153, pause_setI2154, pause_setI2155, pause_setI2156, pause_setI2157, pause_setI2158, pause_setI2159, pause_setI2160, pause_setI2161, pause_setI2162, pause_setI2163, pause_setI2164, pause_setI2165, pause_setI2166, pause_setI2167, pause_setI2168, pause_setI2169, pause_setI2170, pause_setI2171, pause_setI2172, pause_setI2173, pause_setI2174, pause_setI2175, pause_setI2176, pause_setI2177, pause_setI2178, pause_setI2179, pause_setI2180, pause_setI2181, pause_setI2182, pause_setI2183, pause_setI2184, pause_setI2185, pause_setI2186, pause_setI2187, pause_setI2188, pause_setI2189, pause_setI2190, pause_setI2191, pause_setI2192, pause_setI2193, pause_setI2194, pause_setI2195, pause_setI2196, pause_setI2197, pause_setI2198, pause_setI2199, pause_setI2200, pause_setI2201, pause_setI2202, pause_setI2203, pause_setI2204, pause_setI2205, pause_setI2206, pause_setI2207, pause_setI2208, pause_setI2209, pause_setI2210, pause_setI2211, pause_setI2212, pause_setI2213, pause_setI2214, pause_setI2215, pause_setI2216, pause_setI2217, pause_setI2218, pause_setI2219, pause_setI2220, pause_setI2221, pause_setI2222, pause_setI2223, pause_setI2224, pause_setI2225, pause_setI2226, pause_setI2227, pause_setI2228, pause_setI2229, pause_setI2230, pause_setI2231, pause_setI2232, pause_setI2233, pause_setI2234, pause_setI2235, pause_setI2236, pause_setI2237, pause_setI2238, pause_setI2239, pause_setI2240, pause_setI2241, pause_setI2242, pause_setI2243, pause_setI2244, pause_setI2245, pause_setI2246, pause_setI2247, pause_setI2248, pause_setI2249, pause_setI2250, pause_setI2251, pause_setI2252, pause_setI2253, pause_setI2254, pause_setI2255, pause_setI2256, pause_setI2257, pause_setI2258, pause_setI2259, pause_setI2260, pause_setI2261, pause_setI2262, pause_setI2263, pause_setI2264, pause_setI2265, pause_setI2266, pause_setI2267, pause_setI2268, pause_setI2269, pause_setI2270, pause_setI2271, pause_setI2272, pause_setI2273, pause_setI2274, pause_setI2275, pause_setI2276, pause_setI2277, pause_setI2278, pause_setI2279, pause_setI2280, pause_setI2281, pause_setI2282, pause_setI2283, pause_setI2284, pause_setI2285, pause_setI2286, pause_setI2287, pause_setI2288, pause_setI2289, pause_setI2290, pause_setI2291, pause_setI2292, pause_setI2293, pause_setI2294, pause_setI2295, pause_setI2296, pause_setI2297, pause_setI2298, pause_setI2299, pause_setI2300, pause_setI2301, pause_setI2302, pause_setI2303, pause_setI2304, pause_setI2305, pause_setI2306, pause_setI2307, pause_setI2308, pause_setI2309, pause_setI2310, pause_setI2311, pause_setI2312, pause_setI2313, pause_setI2314, pause_setI2315, pause_setI2316, pause_setI2317, pause_setI2318, pause_setI2319, pause_setI2320, pause_setI2321, pause_setI2322, pause_setI2323, pause_setI2324, pause_setI2325, pause_setI2326, pause_setI2327, pause_setI2328, pause_setI2329, pause_setI2330, pause_setI2331, pause_setI2332, pause_setI2333, pause_setI2334, pause_setI2335, pause_setI2336, pause_setI2337, pause_setI2338, pause_setI2339, pause_setI2340, pause_setI2341, pause_setI2342, pause_setI2343, pause_setI2344, pause_setI2345, pause_setI2346, pause_setI2347, pause_setI2348, pause_setI2349, pause_setI2350, pause_setI2351, pause_setI2352, pause_setI2353, pause_setI2354, pause_setI2355, pause_setI2356, pause_setI2357, pause_setI2358, pause_setI2359, pause_setI2360, pause_setI2361, pause_setI2362, pause_setI2363, pause_setI2364, pause_setI2365, pause_setI2366, pause_setI2367, pause_setI2368, pause_setI2369, pause_setI2370, pause_setI2371, pause_setI2372, pause_setI2373, pause_setI2374, pause_setI2375, pause_setI2376, pause_setI2377, pause_setI2378, pause_setI2379, pause_setI2380, pause_setI2381, pause_setI2382, pause_setI2383, pause_setI2384, pause_setI2385, pause_setI2386, pause_setI2387, pause_setI2388, pause_setI2389, pause_setI2390, pause_setI2391, pause_setI2392, pause_setI2393, pause_setI2394, pause_setI2395, pause_setI2396, pause_setI2397, pause_setI2398, pause_setI2399, pause_setI2400, pause_setI2401, pause_setI2402, pause_setI2403, pause_setI2404, pause_setI2405, pause_setI2406, pause_setI2407, pause_setI2408, pause_setI2409, pause_setI2410, pause_setI2411, pause_setI2412, pause_setI2413, pause_setI2414, pause_setI2415, pause_setI2416, pause_setI2417, pause_setI2418, pause_setI2419, pause_setI2420, pause_setI2421, pause_setI2422, pause_setI2423, pause_setI2424, pause_setI2425, pause_setI2426, pause_setI2427, pause_setI2428, pause_setI2429, pause_setI2430, pause_setI2431, pause_setI2432, pause_setI2433, pause_setI2434, pause_setI2435, pause_setI2436, pause_setI2437, pause_setI2438, pause_setI2439, pause_setI2440, pause_setI2441, pause_setI2442, pause_setI2443, pause_setI2444, pause_setI2445, pause_setI2446, pause_setI2447, pause_setI2448, pause_setI2449, pause_setI2450, pause_setI2451, pause_setI2452, pause_setI2453, pause_setI2454, pause_setI2455, pause_setI2456, pause_setI2457, pause_setI2458, pause_setI2459, pause_setI2460, pause_setI2461, pause_setI2462, pause_setI2463, pause_setI2464, pause_setI2465, pause_setI2466, pause_setI2467, pause_setI2468, pause_setI2469, pause_setI2470, pause_setI2471, pause_setI2472, pause_setI2473, pause_setI2474, pause_setI2475, pause_setI2476, pause_setI2477, pause_setI2478, pause_setI2479, pause_setI2480, pause_setI2481, pause_setI2482, pause_setI2483, pause_setI2484, pause_setI2485, pause_setI2486, pause_setI2487, pause_setI2488, pause_setI2489, pause_setI2490, pause_setI2491, pause_setI2492, pause_setI2493, pause_setI2494, pause_setI2495, pause_setI2496, pause_setI2497, pause_setI2498, pause_setI2499, pause_setI2500, pause_setI2501, pause_setI2502, pause_setI2503, pause_setI2504, pause_setI2505, pause_setI2506, pause_setI2507, pause_setI2508, pause_setI2509, pause_setI2510, pause_setI2511, pause_setI2512, pause_setI2513, pause_setI2514, pause_setI2515, pause_setI2516, pause_setI2517, pause_setI2518, pause_setI2519, pause_setI2520, pause_setI2521, pause_setI2522, pause_setI2523, pause_setI2524, pause_setI2525, pause_setI2526, pause_setI2527, pause_setI2528, pause_setI2529, pause_setI2530, pause_setI2531, pause_setI2532, pause_setI2533, pause_setI2534, pause_setI2535, pause_setI2536, pause_setI2537, pause_setI2538, pause_setI2539, pause_setI2540, pause_setI2541, pause_setI2542, pause_setI2543, pause_setI2544, pause_setI2545, pause_setI2546, pause_setI2547, pause_setI2548, pause_setI2549, pause_setI2550, pause_setI2551, pause_setI2552, pause_setI2553, pause_setI2554, pause_setI2555, pause_setI2556, pause_setI2557, pause_setI2558, pause_setI2559, pause_setI2560, pause_setI2561, pause_setI2562, pause_setI2563, pause_setI2564, pause_setI2565, pause_setI2566, pause_setI2567, pause_setI2568, pause_setI2569, pause_setI2570, pause_setI2571, pause_setI2572, pause_setI2573, pause_setI2574, pause_setI2575, pause_setI2576, pause_setI2577, pause_setI2578, pause_setI2579);
  signal state_var3002: t_state_var3002;
  type t_state_var3001 is (compute2589, \$1410_forever\, \$1452_loop\, \$1489_loop\, \$1526_loop\, \$581_loop\, aux, copy_root_in_ram, \loop\, pause_getI2592, pause_getI2598, pause_getI2601, pause_getI2604, pause_getI2609, pause_getI2615, pause_getI2618, pause_getI2621, pause_getI2624, pause_getI2628, pause_getI2631, pause_getI2637, pause_getI2640, pause_getI2644, pause_getI2650, pause_getI2653, pause_getII2593, pause_getII2599, pause_getII2602, pause_getII2605, pause_getII2610, pause_getII2616, pause_getII2619, pause_getII2622, pause_getII2625, pause_getII2629, pause_getII2632, pause_getII2638, pause_getII2641, pause_getII2645, pause_getII2651, pause_getII2654, pause_setI2590, pause_setI2591, pause_setI2595, pause_setI2596, pause_setI2597, pause_setI2607, pause_setI2608, pause_setI2612, pause_setI2613, pause_setI2614, pause_setI2630, pause_setI2634, pause_setI2635, pause_setI2636, pause_setI2643, pause_setI2647, pause_setI2648, pause_setI2649);
  signal state_var3001: t_state_var3001;
  type t_state_var3000 is (compute2584, \$103_w\, \$1278_forever\, \$1281_forever\, \$1284_forever\, \$1342_modulo\, \$74_fill\, \$855_forever\, \$921_forever\, apply, binop_compare, binop_int, branch_if, compare, compbranch, fill, forever, loop_push, make_block, make_block_n, modulo, offsetclosure_n, pause_getI2660, pause_getI2672, pause_getI2675, pause_getI2678, pause_getI2687, pause_getI2690, pause_getI2693, pause_getI2697, pause_getI2702, pause_getI2705, pause_getI2707, pause_getI2709, pause_getI2711, pause_getI2713, pause_getI2715, pause_getI2717, pause_getI2719, pause_getI2723, pause_getI2726, pause_getI2729, pause_getI2732, pause_getI2735, pause_getI2738, pause_getI2741, pause_getI2744, pause_getI2746, pause_getI2748, pause_getI2750, pause_getI2752, pause_getI2755, pause_getI2758, pause_getI2761, pause_getI2765, pause_getI2768, pause_getI2770, pause_getI2776, pause_getI2778, pause_getI2780, pause_getI2782, pause_getI2785, pause_getI2788, pause_getI2791, pause_getI2794, pause_getI2796, pause_getI2798, pause_getI2800, pause_getI2803, pause_getI2805, pause_getI2807, pause_getI2809, pause_getI2812, pause_getI2814, pause_getI2816, pause_getI2818, pause_getI2820, pause_getI2822, pause_getI2824, pause_getI2830, pause_getI2832, pause_getI2836, pause_getI2838, pause_getI2844, pause_getI2846, pause_getI2848, pause_getI2850, pause_getI2852, pause_getI2856, pause_getI2859, pause_getI2861, pause_getI2863, pause_getI2869, pause_getI2871, pause_getI2876, pause_getI2879, pause_getI2881, pause_getI2883, pause_getI2890, pause_getI2894, pause_getI2898, pause_getI2900, pause_getI2904, pause_getI2906, pause_getI2908, pause_getI2912, pause_getI2914, pause_getI2916, pause_getI2918, pause_getI2922, pause_getI2924, pause_getI2926, pause_getI2928, pause_getI2932, pause_getI2935, pause_getI2938, pause_getI2941, pause_getI2947, pause_getI2949, pause_getI2951, pause_getI2953, pause_getI2957, pause_getI2962, pause_getI2966, pause_getI2976, pause_getI2979, pause_getI2982, pause_getI2985, pause_getI2988, pause_getII2661, pause_getII2673, pause_getII2676, pause_getII2679, pause_getII2688, pause_getII2691, pause_getII2694, pause_getII2698, pause_getII2703, pause_getII2706, pause_getII2708, pause_getII2710, pause_getII2712, pause_getII2714, pause_getII2716, pause_getII2718, pause_getII2720, pause_getII2724, pause_getII2727, pause_getII2730, pause_getII2733, pause_getII2736, pause_getII2739, pause_getII2742, pause_getII2745, pause_getII2747, pause_getII2749, pause_getII2751, pause_getII2753, pause_getII2756, pause_getII2759, pause_getII2762, pause_getII2766, pause_getII2769, pause_getII2771, pause_getII2777, pause_getII2779, pause_getII2781, pause_getII2783, pause_getII2786, pause_getII2789, pause_getII2792, pause_getII2795, pause_getII2797, pause_getII2799, pause_getII2801, pause_getII2804, pause_getII2806, pause_getII2808, pause_getII2810, pause_getII2813, pause_getII2815, pause_getII2817, pause_getII2819, pause_getII2821, pause_getII2823, pause_getII2825, pause_getII2831, pause_getII2833, pause_getII2837, pause_getII2839, pause_getII2845, pause_getII2847, pause_getII2849, pause_getII2851, pause_getII2853, pause_getII2857, pause_getII2860, pause_getII2862, pause_getII2864, pause_getII2870, pause_getII2872, pause_getII2877, pause_getII2880, pause_getII2882, pause_getII2884, pause_getII2891, pause_getII2895, pause_getII2899, pause_getII2901, pause_getII2905, pause_getII2907, pause_getII2909, pause_getII2913, pause_getII2915, pause_getII2917, pause_getII2919, pause_getII2923, pause_getII2925, pause_getII2927, pause_getII2929, pause_getII2933, pause_getII2936, pause_getII2939, pause_getII2942, pause_getII2948, pause_getII2950, pause_getII2952, pause_getII2954, pause_getII2958, pause_getII2963, pause_getII2967, pause_getII2977, pause_getII2980, pause_getII2983, pause_getII2986, pause_getII2989, pause_setI2585, pause_setI2662, pause_setI2664, pause_setI2666, pause_setI2668, pause_setI2669, pause_setI2670, pause_setI2692, pause_setI2696, pause_setI2700, pause_setI2721, pause_setI2722, pause_setI2725, pause_setI2728, pause_setI2731, pause_setI2734, pause_setI2737, pause_setI2740, pause_setI2743, pause_setI2754, pause_setI2757, pause_setI2760, pause_setI2763, pause_setI2764, pause_setI2772, pause_setI2773, pause_setI2774, pause_setI2775, pause_setI2784, pause_setI2787, pause_setI2790, pause_setI2793, pause_setI2802, pause_setI2811, pause_setI2826, pause_setI2827, pause_setI2828, pause_setI2829, pause_setI2834, pause_setI2835, pause_setI2840, pause_setI2841, pause_setI2842, pause_setI2843, pause_setI2855, pause_setI2865, pause_setI2866, pause_setI2868, pause_setI2873, pause_setI2874, pause_setI2875, pause_setI2878, pause_setI2886, pause_setI2887, pause_setI2888, pause_setI2889, pause_setI2893, pause_setI2897, pause_setI2903, pause_setI2911, pause_setI2921, pause_setI2930, pause_setI2931, pause_setI2934, pause_setI2940, pause_setI2944, pause_setI2945, pause_setI2955, pause_setI2956, pause_setI2960, pause_setI2961, pause_setI2965, pause_setI2968, pause_setI2970, pause_setI2972, pause_setI2973, pause_setI2974, w, w0, w1, w3, \wait\);
  signal state_var3000: t_state_var3000;
  type array_value_16 is array (natural range <>) of value(0 to 15);
  type array_value_31 is array (natural range <>) of value(0 to 30);
  type array_value_32 is array (natural range <>) of value(0 to 31);
  signal ram : array_value_32(0 to 16383) := (others => "000"& X"000000" & X"0" & eclat_true); 
  signal \$ram_value\ : value(0 to 31);
  signal \$ram_ptr\ : natural range 0 to 16383;
  signal \$ram_ptr_write\ : natural range 0 to 16383;
  signal \$ram_write\ : value(0 to 31);
  signal \$ram_write_request\ : std_logic := '0';
  signal global_end : array_value_16(0 to 0) := (others => X"000" & X"0"); 
  signal \$global_end_value\ : value(0 to 15);
  signal \$global_end_ptr\ : natural range 0 to 0;
  signal \$global_end_ptr_write\ : natural range 0 to 0;
  signal \$global_end_write\ : value(0 to 15);
  signal \$global_end_write_request\ : std_logic := '0';
  signal code : array_value_31(0 to 423) := (others => "000"& X"000000" & X"0"); 
  signal \$code_value\ : value(0 to 30);
  signal \$code_ptr\ : natural range 0 to 423;
  signal \$code_ptr_write\ : natural range 0 to 423;
  signal \$code_write\ : value(0 to 30);
  signal \$code_write_request\ : std_logic := '0';
  
  begin
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$ram_write_request\ = '1' then
                    ram(\$ram_ptr_write\) <= \$ram_write\;
                  else
                   \$ram_value\ <= ram(\$ram_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$global_end_write_request\ = '1' then
                    global_end(\$global_end_ptr_write\) <= \$global_end_write\;
                  else
                   \$global_end_value\ <= global_end(\$global_end_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$code_write_request\ = '1' then
                    code(\$code_ptr_write\) <= \$code_write\;
                  else
                   \$code_value\ <= code(\$code_ptr\);
                  end if;
            end if;
        end process;
    
    process(clk)
      variable \$v932\ : value(0 to 1) := (others => '0');
      variable loop_arg, \$v584\, make_block_result, \$v576\, \$v866\, 
               \$v593\, w0_arg, \$v620\, \$v540\ : value(0 to 95) := (others => '0');
      variable compare_arg : value(0 to 93) := (others => '0');
      variable \$v814\, \$v908\, \$v624\, \$v810\, \$v830\, \$v1433\, 
               \$v625\, \$v615\, \$v701\, \$v1409\, \$v707\, \$v827\, 
               \$v871\, \$v599\, \$v563\, \$v668\, \$v87\, \$v796\, \$v649\, 
               \$v722\, \$v632\, \$v623\, \$v886\, \$v718\, \$v813\, \$v906\, 
               \$v676\, \$v703\, \$v715\, \$v581\, \$v805\, \$v822\, \$v829\, 
               \$v868\, \$v689\, \$v688\, \$v878\, \$v1468\, \$v818\, 
               \$v717\, \$v832\, \$v799\, \$v680\, \$v702\, \$v821\, \$v831\, 
               \$v802\, \$v614\, \$v613\, \$v907\, \$v1408\, \$v693\, \$v716\ : value(0 to 47) := (others => '0');
      variable \$1526_loop_arg\, aux_arg, loop_push_arg, \$103_w_arg\, 
               \$1452_loop_arg\, \$581_loop_arg\, w_arg, \$1489_loop_arg\ : value(0 to 63) := (others => '0');
      variable branch_if_arg, \$v524\, \$v518\, \$v522\ : value(0 to 122) := (others => '0');
      variable \$v2981\, \$v2978\, \$v2987\, \$v2984\ : value(0 to 7) := (others => '0');
      variable \$235_sp\, \$1008_sp\, \$210_sp\, \$35_sp\, fill_result, 
               \$558_next\, \$33_sp\, \$1100_sp\, \$342_sp\, \$1048_sp\, 
               \$84_sp\, copy_root_in_ram_result, \$1271_sp\, \$1267_sp\, 
               \$1057_sp\, \$341_sp\, \$v407\, \$983_sp\, \$354_sp\, 
               \$1103_sp\, \$1263_sp\, \$59_sp\, \$133_sp\, \$562_next\, 
               \$557_next\, loop_push_result, \$241_sp\, idx, \$324_sp\, 
               \$123_sp\, \$166_sp\, \$83_sp\, \$1075_sp\, \$988_sp\, 
               \$125_ofs\, \$104_sp\, \$289_sp\, \$148_sp\, \$75_sp\, 
               \$74_fill_result\, \$128_sp\, \$1003_sp\, \$993_sp\, 
               \$242_sp\, \$351_sp\, \$187_sp\, \$131_sp\, \$127_sp\, 
               \$556_next\, \$30_sp\, \$339_sp\, \$55_sp\, \$1106_sp\, 
               \$1066_sp\, \$1275_sp\, w0_result, \$981_sp\, \$1013_sp\, 
               \$347_sp\, \$364_sp\, \$81_sp\, \$998_sp\, \$39_sp\, 
               \$288_sp\, \$v234\, aux_result, w3_result, \$345_sp\, 
               \$130_sp\, \$346_sp\, \$340_sp\, \$34_sp\, \$357_sp\, 
               \$103_w_result\, loop_result, \$v227\ : value(0 to 15) := (others => '0');
      variable \$v509\ : value(0 to 2) := (others => '0');
      variable \$1342_modulo_arg\, modulo_arg : value(0 to 61) := (others => '0');
      variable wait_arg : value(0 to 96) := (others => '0');
      variable result2132 : value(0 to 57) := (others => '0');
      variable copy_root_in_ram_id, make_block_id, compare_id : value(0 to 11) := (others => '0');
      variable compbranch_arg : value(0 to 215) := (others => '0');
      variable \$v515\, \$v516\ : value(0 to 3) := (others => '0');
      variable \$1342_modulo_result\, modulo_result, \$v179\, \$v2910\, 
               \$313_res\, \$v2920\, \$1343_r\, \$v29\, arg, \$v44\, r, 
               \$v2896\, \$v2892\, \$v259\, argument3, argument1, \$v2902\, 
               argument2 : value(0 to 30) := (others => '0');
      variable offsetclosure_n_arg : value(0 to 137) := (others => '0');
      variable result2587 : value(0 to 127) := (others => '0');
      variable make_block_arg : value(0 to 103) := (others => '0');
      variable \$233_b\, \$v2652\, \$v2998\, \$v2136\, \$v2854\, \$v2617\, 
               \$v2990\, rdy2588, \$v2646\, \$v2997\, \$581_loop_result\, 
               \$v2627\, \$v2999\, \$v1397_init_done\, \$v2581\, \$v2656\, 
               \$v2964\, \$v516_init_done\, \$v2704\, \$v2971\, \$v2680\, 
               \$v2135\, \$v2674\, \$v2993\, \$v2699\, \$v2594\, \$v2937\, 
               \$v2701\, \$1452_loop_result\, result2138, \$v2684\, rdy2583, 
               \$v2975\, \$v2626\, \$v2991\, \$v2969\, \$v2683\, \$v2867\, 
               \$v2586\, \$v2681\, \$v2767\, \$v522_init_done\, \$v2620\, 
               \$300_res\, \$v2642\, \$1489_loop_result\, \$v2606\, \$v2600\, 
               \$v2667\, \$1526_loop_result\, \$v2659\, \$v2943\, \$v2137\, 
               \$v2677\, \$v934\, \$v2663\, \$v2682\, \$v2623\, \$v2685\, 
               \$v2665\, \$v2671\, \$v2996\, \$v2611\, \$v511_init_done\, 
               \$v2695\, \$v1377_init_done\, \$v2603\, \$v2959\, \$v2633\, 
               \$v2639\, \$v2858\, \$v2658\, rdy2139, \$v2995\, \$v2994\, 
               \$12_rdy\, \$v2655\, b, rdy2133, w1_result, \$v934_init_done\, 
               w_result, \$v2946\, compare_result, \$v2885\ : value(0 to 0) := (others => '0');
      variable apply_arg : value(0 to 165) := (others => '0');
      variable make_block_n_arg : value(0 to 171) := (others => '0');
      variable fill_arg, \$v51\, \$74_fill_arg\, w3_arg, wait_result, 
               \$v1400\, w1_arg, copy_root_in_ram_arg, \$v1380\ : value(0 to 79) := (others => '0');
      variable \$v1397\, \$v1395\ : value(0 to 128) := (others => '0');
      variable \$236_next_env\, \$66_v\, \$967_v\, \$1315_v\, \$955_v\, 
               \$1200_v\, \$v86\, \$1218_v\, \$989_v\, \$v18\, \$v146\, 
               \$902_v\, \$1501\, \$1464\, \$1067\, \$1208_v\, \$1014_v\, 
               \$916_v\, \$1041\, \$1353_v\, \$817_v\, \$660_v\, \$1308_v\, 
               \$v287\, \$368_v\, \$971_v\, \$1226_v\, \$1033\, \$918_v\, 
               \$1449_hd\, cy, \$800_v\, \$1383_v\, \$1183_v\, \$878_v\, 
               \$v402\, \$1025\, \$1241_v\, \$826_v\, \$770_v\, \$898_v\, 
               \$1058\, \$1249_v\, \$v2686\, \$1153_v\, \$912_v\, \$1538\, 
               \$864_v\, \$1228_v\, \$1049\, \$578_w\, \$1004_v\, \$v274\, 
               \$975_v\, \$120_v\, \$900_v\, \$979_v\, \$1379_v\, \$914_v\, 
               \$890_v\, \$1523_hd\, \$876_v\, \$1330_v\, \$v412\, \$888_v\, 
               \$v225\, \$579_hd\, \$959_v\, \$1239_v\, \$592_hd\, \$v80\, 
               \$1076\, \$1139_v\, \$904_v\, \$1163_v\, \$70_v\, \$1009_v\, 
               \$886_v\, \$1447_w\, \$1235_v\, f0, \$852_v\, \$984_v\, 
               \$778\, \$v400\, \$321_v\, \$v134\, \$1245_v\, \$1129_v\, 
               \$963_v\, \$v426\, \$1486_hd\, \$735_v\, \$796_v\, \$1484_w\, 
               \$794_v\, \$v100\, \$951_v\, \$v1377\, \$1109_v\, \$1210_v\, 
               \$1186_hd\, \$245_v\, \$811_v\, \$813_v\, \$253_next_acc\, 
               \$868_v\, \$1119_v\, \$v104\, \$762_v\, \$1173_v\, \$1521_w\, 
               \$122_v\, \$v2689\, \$590_hd\, \$1017\, \$1381_v\, \$999_v\, 
               \$994_v\, \$v511\ : value(0 to 31) := (others => '0');
      variable \$v677\, \$v704\, binop_int_arg, \$v690\, \$v665\, 
               binop_compare_arg, \$v719\ : value(0 to 153) := (others => '0');
      variable binop_compare_result, apply_result, result2582, 
               make_block_n_result, branch_if_result, offsetclosure_n_result, 
               compbranch_result, binop_int_result : value(0 to 121) := (others => '0');
      
    begin
      
      if rising_edge(clk) then
        if (reset = '1') then
          default_zero(\$v1380\); default_zero(\$v227\); 
          default_zero(loop_result); default_zero(\$v719\); 
          default_zero(binop_compare_arg); default_zero(\$v511\); 
          default_zero(\$v2885\); default_zero(\$1489_loop_arg\); 
          default_zero(compare_result); default_zero(\$103_w_result\); 
          default_zero(\$357_sp\); default_zero(\$v2946\); 
          default_zero(\$994_v\); default_zero(w_result); 
          default_zero(\$34_sp\); default_zero(\$340_sp\); 
          default_zero(\$999_v\); default_zero(\$1381_v\); 
          default_zero(\$v934_init_done\); default_zero(\$346_sp\); 
          default_zero(\$130_sp\); default_zero(\$1017\); 
          default_zero(w1_result); default_zero(w_arg); 
          default_zero(\$590_hd\); default_zero(modulo_arg); 
          default_zero(rdy2133); default_zero(\$345_sp\); 
          default_zero(w3_result); default_zero(\$v2984\); 
          default_zero(\$v2689\); default_zero(\$122_v\); 
          default_zero(\$v540\); default_zero(b); default_zero(\$1521_w\); 
          default_zero(\$v716\); default_zero(\$1173_v\); 
          default_zero(aux_result); default_zero(\$v2655\); 
          default_zero(\$762_v\); default_zero(\$v693\); 
          default_zero(\$v234\); default_zero(compare_arg); 
          default_zero(\$v104\); default_zero(\$1119_v\); 
          default_zero(\$868_v\); default_zero(\$v1408\); 
          default_zero(\$253_next_acc\); default_zero(\$581_loop_arg\); 
          default_zero(\$288_sp\); default_zero(\$v932\); 
          default_zero(\$39_sp\); default_zero(\$813_v\); 
          default_zero(\$v620\); default_zero(\$811_v\); 
          default_zero(\$998_sp\); default_zero(\$81_sp\); 
          default_zero(\$v665\); default_zero(\$v907\); 
          default_zero(\$12_rdy\); default_zero(copy_root_in_ram_arg); 
          default_zero(\$364_sp\); default_zero(\$347_sp\); 
          default_zero(\$245_v\); default_zero(\$1186_hd\); 
          default_zero(w0_arg); default_zero(\$v2994\); 
          default_zero(\$v2995\); default_zero(\$1013_sp\); 
          default_zero(rdy2139); default_zero(binop_int_result); 
          default_zero(\$1210_v\); default_zero(\$1109_v\); 
          default_zero(\$v1377\); default_zero(\$v690\); 
          default_zero(\$v516\); default_zero(\$981_sp\); 
          default_zero(\$v2658\); default_zero(\$951_v\); 
          default_zero(\$v593\); default_zero(w0_result); 
          default_zero(\$1275_sp\); default_zero(\$v100\); 
          default_zero(\$v2858\); default_zero(w1_arg); 
          default_zero(\$794_v\); default_zero(\$1342_modulo_arg\); 
          default_zero(\$1484_w\); default_zero(\$v613\); 
          default_zero(\$796_v\); default_zero(\$v2639\); 
          default_zero(\$v614\); default_zero(\$1066_sp\); 
          default_zero(\$v2633\); default_zero(\$v2959\); 
          default_zero(\$v2603\); default_zero(\$735_v\); 
          default_zero(\$1106_sp\); default_zero(\$v802\); 
          default_zero(\$55_sp\); default_zero(\$339_sp\); 
          default_zero(\$v831\); default_zero(\$v1377_init_done\); 
          default_zero(\$30_sp\); default_zero(\$1486_hd\); 
          default_zero(\$v2695\); default_zero(\$v426\); 
          default_zero(\$556_next\); default_zero(compbranch_result); 
          default_zero(make_block_arg); default_zero(\$v511_init_done\); 
          default_zero(\$v2611\); default_zero(\$v1400\); 
          default_zero(\$127_sp\); default_zero(\$v2996\); 
          default_zero(\$131_sp\); default_zero(\$963_v\); 
          default_zero(\$v866\); default_zero(\$v821\); 
          default_zero(\$1129_v\); default_zero(\$1245_v\); 
          default_zero(\$v2671\); default_zero(argument2); 
          default_zero(\$v576\); default_zero(\$v1395\); 
          default_zero(\$187_sp\); default_zero(\$v702\); 
          default_zero(\$351_sp\); default_zero(\$242_sp\); 
          default_zero(\$993_sp\); default_zero(make_block_result); 
          default_zero(\$v2665\); default_zero(\$v2902\); 
          default_zero(\$v134\); default_zero(\$321_v\); 
          default_zero(\$v400\); default_zero(\$1003_sp\); 
          default_zero(\$v680\); default_zero(\$778\); 
          default_zero(\$128_sp\); default_zero(\$984_v\); 
          default_zero(wait_result); default_zero(\$74_fill_result\); 
          default_zero(\$75_sp\); default_zero(\$148_sp\); 
          default_zero(\$852_v\); default_zero(f0); default_zero(\$289_sp\); 
          default_zero(wait_arg); default_zero(\$v2685\); 
          default_zero(argument1); default_zero(\$1235_v\); 
          default_zero(\$1447_w\); default_zero(\$886_v\); 
          default_zero(\$v2623\); default_zero(\$1009_v\); 
          default_zero(make_block_n_arg); default_zero(\$v799\); 
          default_zero(\$v832\); default_zero(\$70_v\); 
          default_zero(\$1163_v\); default_zero(\$v584\); 
          default_zero(\$904_v\); default_zero(\$v2682\); 
          default_zero(\$v522\); default_zero(\$104_sp\); 
          default_zero(\$1452_loop_arg\); default_zero(\$1139_v\); 
          default_zero(\$1076\); default_zero(offsetclosure_n_result); 
          default_zero(\$v2663\); default_zero(\$103_w_arg\); 
          default_zero(\$v717\); default_zero(\$v80\); 
          default_zero(\$125_ofs\); default_zero(\$592_hd\); 
          default_zero(\$v934\); default_zero(\$988_sp\); 
          default_zero(loop_push_arg); default_zero(\$v2677\); 
          default_zero(\$v2137\); default_zero(\$v2943\); 
          default_zero(\$v818\); default_zero(\$1075_sp\); 
          default_zero(result2587); default_zero(compbranch_arg); 
          default_zero(compare_id); default_zero(\$1239_v\); 
          default_zero(apply_arg); default_zero(\$959_v\); 
          default_zero(\$83_sp\); default_zero(\$579_hd\); 
          default_zero(\$166_sp\); default_zero(\$v225\); 
          default_zero(branch_if_result); default_zero(\$v518\); 
          default_zero(\$v1468\); default_zero(\$v2659\); 
          default_zero(\$1526_loop_result\); default_zero(\$888_v\); 
          default_zero(\$v2667\); default_zero(\$v412\); 
          default_zero(\$1330_v\); default_zero(loop_arg); 
          default_zero(\$876_v\); default_zero(\$v2600\); 
          default_zero(\$123_sp\); default_zero(\$v878\); 
          default_zero(\$v2606\); default_zero(\$v1397\); 
          default_zero(\$324_sp\); default_zero(\$1489_loop_result\); 
          default_zero(\$v688\); default_zero(\$1523_hd\); 
          default_zero(\$890_v\); default_zero(\$v689\); 
          default_zero(\$914_v\); default_zero(\$v2642\); default_zero(idx); 
          default_zero(\$1379_v\); default_zero(\$v868\); 
          default_zero(\$v829\); default_zero(\$979_v\); 
          default_zero(\$300_res\); default_zero(\$900_v\); 
          default_zero(binop_int_arg); default_zero(\$241_sp\); 
          default_zero(argument3); default_zero(loop_push_result); 
          default_zero(\$v2620\); default_zero(\$v822\); 
          default_zero(\$v805\); default_zero(\$v2987\); 
          default_zero(\$557_next\); default_zero(\$v259\); 
          default_zero(\$v522_init_done\); default_zero(\$v2767\); 
          default_zero(\$v2892\); default_zero(\$120_v\); 
          default_zero(\$v2896\); default_zero(\$975_v\); 
          default_zero(\$v581\); default_zero(aux_arg); 
          default_zero(make_block_n_result); default_zero(\$v274\); 
          default_zero(\$1004_v\); default_zero(result2582); 
          default_zero(\$v2978\); default_zero(\$v2681\); 
          default_zero(\$562_next\); default_zero(\$v2981\); 
          default_zero(\$v2586\); default_zero(\$v2867\); default_zero(r); 
          default_zero(\$133_sp\); default_zero(\$578_w\); 
          default_zero(\$59_sp\); default_zero(\$v2683\); 
          default_zero(\$v2969\); default_zero(\$v44\); 
          default_zero(\$1263_sp\); default_zero(\$1103_sp\); 
          default_zero(arg); default_zero(\$v715\); default_zero(\$354_sp\); 
          default_zero(\$1049\); default_zero(\$v29\); 
          default_zero(\$1228_v\); default_zero(\$v703\); 
          default_zero(\$864_v\); default_zero(\$v2991\); 
          default_zero(\$1538\); default_zero(\$v2626\); 
          default_zero(\$912_v\); default_zero(\$v676\); 
          default_zero(\$983_sp\); default_zero(\$v407\); 
          default_zero(result2132); default_zero(\$v906\); 
          default_zero(\$341_sp\); default_zero(\$1153_v\); 
          default_zero(\$1057_sp\); default_zero(\$v2686\); 
          default_zero(\$v813\); default_zero(make_block_id); 
          default_zero(\$v704\); default_zero(\$1249_v\); 
          default_zero(\$v2975\); default_zero(\$1267_sp\); 
          default_zero(\$v718\); default_zero(\$1271_sp\); 
          default_zero(\$1058\); default_zero(\$1343_r\); 
          default_zero(\$898_v\); default_zero(\$770_v\); 
          default_zero(rdy2583); default_zero(copy_root_in_ram_result); 
          default_zero(\$v886\); default_zero(\$826_v\); 
          default_zero(\$v2684\); default_zero(\$v2920\); 
          default_zero(result2138); default_zero(\$1452_loop_result\); 
          default_zero(\$v509\); default_zero(\$v623\); 
          default_zero(\$1241_v\); default_zero(\$1025\); 
          default_zero(\$v632\); default_zero(\$v402\); 
          default_zero(\$878_v\); default_zero(\$1183_v\); 
          default_zero(\$v2701\); default_zero(\$v2937\); 
          default_zero(\$v2594\); default_zero(\$v2699\); 
          default_zero(\$1383_v\); default_zero(\$v722\); 
          default_zero(\$313_res\); default_zero(\$800_v\); default_zero(cy); 
          default_zero(\$1449_hd\); default_zero(\$918_v\); 
          default_zero(\$1033\); default_zero(\$v2993\); 
          default_zero(\$v2674\); default_zero(\$1226_v\); 
          default_zero(\$v2135\); default_zero(\$971_v\); 
          default_zero(\$v649\); default_zero(\$368_v\); 
          default_zero(\$v287\); default_zero(\$1308_v\); 
          default_zero(\$84_sp\); default_zero(\$v2680\); 
          default_zero(\$v2971\); default_zero(\$v2910\); 
          default_zero(\$660_v\); default_zero(\$v796\); 
          default_zero(\$1048_sp\); default_zero(w3_arg); 
          default_zero(\$v87\); default_zero(\$817_v\); 
          default_zero(\$v668\); default_zero(\$1353_v\); 
          default_zero(\$v563\); default_zero(\$v599\); 
          default_zero(\$342_sp\); default_zero(\$1041\); 
          default_zero(\$v524\); default_zero(copy_root_in_ram_id); 
          default_zero(\$74_fill_arg\); default_zero(\$v2704\); 
          default_zero(\$v677\); default_zero(\$916_v\); 
          default_zero(\$v871\); default_zero(\$v516_init_done\); 
          default_zero(\$v827\); default_zero(\$1014_v\); 
          default_zero(\$v515\); default_zero(\$1208_v\); 
          default_zero(\$1067\); default_zero(\$v179\); 
          default_zero(\$1464\); default_zero(\$v2964\); 
          default_zero(\$1501\); default_zero(modulo_result); 
          default_zero(\$902_v\); default_zero(\$v2656\); 
          default_zero(\$v2581\); default_zero(\$v146\); 
          default_zero(apply_result); default_zero(offsetclosure_n_arg); 
          default_zero(\$v18\); default_zero(\$v707\); 
          default_zero(\$1100_sp\); default_zero(\$989_v\); 
          default_zero(\$v1397_init_done\); default_zero(\$v2999\); 
          default_zero(\$v2627\); default_zero(binop_compare_result); 
          default_zero(\$581_loop_result\); default_zero(\$v2997\); 
          default_zero(\$1218_v\); default_zero(\$v1409\); 
          default_zero(\$33_sp\); default_zero(\$v701\); 
          default_zero(\$1526_loop_arg\); 
          default_zero(\$1342_modulo_result\); default_zero(\$v51\); 
          default_zero(\$v2646\); default_zero(\$v615\); 
          default_zero(\$v86\); default_zero(\$558_next\); 
          default_zero(rdy2588); default_zero(\$1200_v\); 
          default_zero(\$v625\); default_zero(\$955_v\); 
          default_zero(\$1315_v\); default_zero(\$v1433\); 
          default_zero(\$v2990\); default_zero(fill_result); 
          default_zero(\$35_sp\); default_zero(\$210_sp\); 
          default_zero(\$967_v\); default_zero(\$v2617\); 
          default_zero(\$v2854\); default_zero(\$v830\); 
          default_zero(\$v810\); default_zero(branch_if_arg); 
          default_zero(\$66_v\); default_zero(\$v624\); 
          default_zero(\$1008_sp\); default_zero(\$235_sp\); 
          default_zero(\$236_next_env\); default_zero(fill_arg); 
          default_zero(\$v908\); default_zero(\$v2136\); 
          default_zero(\$v814\); default_zero(\$v2998\); 
          default_zero(\$v2652\); default_zero(\$233_b\); 
          rdy <= "1";
          rdy2133 := "0";
          state <= compute2134;
          state_var3002 <= compute2140;
          state_var3001 <= compute2589;
          state_var3000 <= compute2584;
          
        else if run = '1' then
          case state is
          when compute2134 =>
            rdy2133 := eclat_false;
            \$v2999\ := eclat_not(""&argument(10));
            if \$v2999\(0) = '1' then
              result2132 := ""&argument(11) & ""&argument(11) & ""&argument(11) & ""&argument(11) & ""&argument(11) & ""&argument(11) & ""&argument(11) & ""&argument(11) & ""&argument(11) & ""&argument(11) & X"63" & X"0" & X"3" & X"71" & X"71" & X"61" & X"61";
              rdy2133 := eclat_true;
              state <= compute2134;
            else
              \$v2998\ := eclat_not(\$v1377_init_done\);
              if \$v2998\(0) = '1' then
                \$v1377\ := X"0000000" & X"0";
                \$v1377_init_done\ := eclat_true;
              end if;
              \$v1377\ := eclat_if(""&argument(11) & X"0000000" & X"0" & eclat_add(\$v1377\ & X"0000000" & X"1"));
              cy := \$v1377\;
              \$v2997\ := eclat_not(\$v516_init_done\);
              if \$v2997\(0) = '1' then
                \$v516\ := eclat_false & eclat_false & eclat_false & eclat_false;
                \$v516_init_done\ := eclat_true;
              end if;
              \$v2996\ := eclat_not(""&\$v516\(2));
              if \$v2996\(0) = '1' then
                case state_var3002 is
                when pause_setI2141 =>
                  \$code_write_request\ <= '0';
                  result2138 := eclat_unit;
                  rdy2139 := eclat_true;
                  state_var3002 <= compute2140;
                when pause_setI2142 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 423;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"8f";
                  state_var3002 <= pause_setI2141;
                when pause_setI2143 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 422;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"5";
                  state_var3002 <= pause_setI2142;
                when pause_setI2144 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 421;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"13";
                  state_var3002 <= pause_setI2143;
                when pause_setI2145 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 420;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"2";
                  state_var3002 <= pause_setI2144;
                when pause_setI2146 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 419;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"13";
                  state_var3002 <= pause_setI2145;
                when pause_setI2147 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 418;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"00000" & X"10");
                  state_var3002 <= pause_setI2146;
                when pause_setI2148 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 417;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"55";
                  state_var3002 <= pause_setI2147;
                when pause_setI2149 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 416;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"7a";
                  state_var3002 <= pause_setI2148;
                when pause_setI2150 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 415;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2149;
                when pause_setI2151 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 414;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"2";
                  state_var3002 <= pause_setI2150;
                when pause_setI2152 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 413;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"14";
                  state_var3002 <= pause_setI2151;
                when pause_setI2153 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 412;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2152;
                when pause_setI2154 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 411;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"7f";
                  state_var3002 <= pause_setI2153;
                when pause_setI2155 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 410;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"9";
                  state_var3002 <= pause_setI2154;
                when pause_setI2156 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 409;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2155;
                when pause_setI2157 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 408;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2156;
                when pause_setI2158 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 407;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"5d";
                  state_var3002 <= pause_setI2157;
                when pause_setI2159 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 406;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"21";
                  state_var3002 <= pause_setI2158;
                when pause_setI2160 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 405;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"e";
                  state_var3002 <= pause_setI2159;
                when pause_setI2161 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 404;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"7";
                  state_var3002 <= pause_setI2160;
                when pause_setI2162 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 403;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"67";
                  state_var3002 <= pause_setI2161;
                when pause_setI2163 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 402;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"5c";
                  state_var3002 <= pause_setI2162;
                when pause_setI2164 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 401;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"12";
                  state_var3002 <= pause_setI2163;
                when pause_setI2165 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 400;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"55";
                  state_var3002 <= pause_setI2164;
                when pause_setI2166 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 399;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"7d";
                  state_var3002 <= pause_setI2165;
                when pause_setI2167 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 398;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"c";
                  state_var3002 <= pause_setI2166;
                when pause_setI2168 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 397;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"9";
                  state_var3002 <= pause_setI2167;
                when pause_setI2169 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 396;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"b";
                  state_var3002 <= pause_setI2168;
                when pause_setI2170 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 395;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"69";
                  state_var3002 <= pause_setI2169;
                when pause_setI2171 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 394;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"69";
                  state_var3002 <= pause_setI2170;
                when pause_setI2172 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 393;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"00000" & X"76");
                  state_var3002 <= pause_setI2171;
                when pause_setI2173 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 392;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2172;
                when pause_setI2174 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 391;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"2b";
                  state_var3002 <= pause_setI2173;
                when pause_setI2175 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 390;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"12";
                  state_var3002 <= pause_setI2174;
                when pause_setI2176 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 389;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"39";
                  state_var3002 <= pause_setI2175;
                when pause_setI2177 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 388;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"00000" & X"57");
                  state_var3002 <= pause_setI2176;
                when pause_setI2178 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 387;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2177;
                when pause_setI2179 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 386;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"2b";
                  state_var3002 <= pause_setI2178;
                when pause_setI2180 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 385;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"16";
                  state_var3002 <= pause_setI2179;
                when pause_setI2181 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 384;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"39";
                  state_var3002 <= pause_setI2180;
                when pause_setI2182 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 383;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2181;
                when pause_setI2183 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 382;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"00000" & X"b9");
                  state_var3002 <= pause_setI2182;
                when pause_setI2184 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 381;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2183;
                when pause_setI2185 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 380;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2184;
                when pause_setI2186 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 379;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"2c";
                  state_var3002 <= pause_setI2185;
                when pause_setI2187 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 378;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"13";
                  state_var3002 <= pause_setI2186;
                when pause_setI2188 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 377;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"39";
                  state_var3002 <= pause_setI2187;
                when pause_setI2189 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 376;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"00000" & X"20");
                  state_var3002 <= pause_setI2188;
                when pause_setI2190 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 375;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2189;
                when pause_setI2191 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 374;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"2b";
                  state_var3002 <= pause_setI2190;
                when pause_setI2192 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 373;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"11";
                  state_var3002 <= pause_setI2191;
                when pause_setI2193 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 372;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"39";
                  state_var3002 <= pause_setI2192;
                when pause_setI2194 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 371;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"21";
                  state_var3002 <= pause_setI2193;
                when pause_setI2195 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 370;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"c";
                  state_var3002 <= pause_setI2194;
                when pause_setI2196 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 369;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"64";
                  state_var3002 <= pause_setI2195;
                when pause_setI2197 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 368;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"14";
                  state_var3002 <= pause_setI2196;
                when pause_setI2198 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 367;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"39";
                  state_var3002 <= pause_setI2197;
                when pause_setI2199 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 366;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2198;
                when pause_setI2200 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 365;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"00000" & X"bd");
                  state_var3002 <= pause_setI2199;
                when pause_setI2201 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 364;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2200;
                when pause_setI2202 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 363;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2201;
                when pause_setI2203 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 362;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"2c";
                  state_var3002 <= pause_setI2202;
                when pause_setI2204 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 361;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"00000" & X"cf");
                  state_var3002 <= pause_setI2203;
                when pause_setI2205 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 360;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2204;
                when pause_setI2206 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 359;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2205;
                when pause_setI2207 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 358;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"2c";
                  state_var3002 <= pause_setI2206;
                when pause_setI2208 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 357;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"4";
                  state_var3002 <= pause_setI2207;
                when pause_setI2209 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 356;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"25";
                  state_var3002 <= pause_setI2208;
                when pause_setI2210 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 355;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"b";
                  state_var3002 <= pause_setI2209;
                when pause_setI2211 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 354;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2210;
                when pause_setI2212 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 353;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"40";
                  state_var3002 <= pause_setI2211;
                when pause_setI2213 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 352;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"d";
                  state_var3002 <= pause_setI2212;
                when pause_setI2214 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 351;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"63";
                  state_var3002 <= pause_setI2213;
                when pause_setI2215 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 350;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"00000" & X"22");
                  state_var3002 <= pause_setI2214;
                when pause_setI2216 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 349;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2215;
                when pause_setI2217 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 348;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2216;
                when pause_setI2218 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 347;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"2c";
                  state_var3002 <= pause_setI2217;
                when pause_setI2219 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 346;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2218;
                when pause_setI2220 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 345;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2219;
                when pause_setI2221 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 344;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"2a";
                  state_var3002 <= pause_setI2220;
                when pause_setI2222 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 343;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"29";
                  state_var3002 <= pause_setI2221;
                when pause_setI2223 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 342;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"4";
                  state_var3002 <= pause_setI2222;
                when pause_setI2224 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 341;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"25";
                  state_var3002 <= pause_setI2223;
                when pause_setI2225 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 340;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"c";
                  state_var3002 <= pause_setI2224;
                when pause_setI2226 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 339;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"36";
                  state_var3002 <= pause_setI2225;
                when pause_setI2227 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 338;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2226;
                when pause_setI2228 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 337;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"5";
                  state_var3002 <= pause_setI2227;
                when pause_setI2229 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 336;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"25";
                  state_var3002 <= pause_setI2228;
                when pause_setI2230 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 335;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"32";
                  state_var3002 <= pause_setI2229;
                when pause_setI2231 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 334;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2230;
                when pause_setI2232 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 333;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"40";
                  state_var3002 <= pause_setI2231;
                when pause_setI2233 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 332;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"44";
                  state_var3002 <= pause_setI2232;
                when pause_setI2234 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 331;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"c";
                  state_var3002 <= pause_setI2233;
                when pause_setI2235 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 330;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2234;
                when pause_setI2236 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 329;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"40";
                  state_var3002 <= pause_setI2235;
                when pause_setI2237 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 328;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"b";
                  state_var3002 <= pause_setI2236;
                when pause_setI2238 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 327;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"c";
                  state_var3002 <= pause_setI2237;
                when pause_setI2239 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 326;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"21";
                  state_var3002 <= pause_setI2238;
                when pause_setI2240 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 325;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"1b";
                  state_var3002 <= pause_setI2239;
                when pause_setI2241 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 324;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"43";
                  state_var3002 <= pause_setI2240;
                when pause_setI2242 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 323;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2241;
                when pause_setI2243 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 322;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"10";
                  state_var3002 <= pause_setI2242;
                when pause_setI2244 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 321;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"56";
                  state_var3002 <= pause_setI2243;
                when pause_setI2245 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 320;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"a";
                  state_var3002 <= pause_setI2244;
                when pause_setI2246 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 319;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"43";
                  state_var3002 <= pause_setI2245;
                when pause_setI2247 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 318;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"b";
                  state_var3002 <= pause_setI2246;
                when pause_setI2248 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 317;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"44";
                  state_var3002 <= pause_setI2247;
                when pause_setI2249 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 316;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2248;
                when pause_setI2250 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 315;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2249;
                when pause_setI2251 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 314;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"28";
                  state_var3002 <= pause_setI2250;
                when pause_setI2252 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 313;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"64";
                  state_var3002 <= pause_setI2251;
                when pause_setI2253 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 312;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"4";
                  state_var3002 <= pause_setI2252;
                when pause_setI2254 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 311;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"27";
                  state_var3002 <= pause_setI2253;
                when pause_setI2255 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 310;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"16";
                  state_var3002 <= pause_setI2254;
                when pause_setI2256 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 309;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"36";
                  state_var3002 <= pause_setI2255;
                when pause_setI2257 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 308;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"69";
                  state_var3002 <= pause_setI2256;
                when pause_setI2258 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 307;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"43";
                  state_var3002 <= pause_setI2257;
                when pause_setI2259 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 306;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"b";
                  state_var3002 <= pause_setI2258;
                when pause_setI2260 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 305;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"44";
                  state_var3002 <= pause_setI2259;
                when pause_setI2261 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 304;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2260;
                when pause_setI2262 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 303;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"a";
                  state_var3002 <= pause_setI2261;
                when pause_setI2263 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 302;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"56";
                  state_var3002 <= pause_setI2262;
                when pause_setI2264 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 301;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2263;
                when pause_setI2265 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 300;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"5";
                  state_var3002 <= pause_setI2264;
                when pause_setI2266 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 299;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"25";
                  state_var3002 <= pause_setI2265;
                when pause_setI2267 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 298;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"15";
                  state_var3002 <= pause_setI2266;
                when pause_setI2268 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 297;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"36";
                  state_var3002 <= pause_setI2267;
                when pause_setI2269 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 296;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"21";
                  state_var3002 <= pause_setI2268;
                when pause_setI2270 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 295;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"b";
                  state_var3002 <= pause_setI2269;
                when pause_setI2271 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 294;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"3";
                  state_var3002 <= pause_setI2270;
                when pause_setI2272 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 293;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"00000" & X"35");
                  state_var3002 <= pause_setI2271;
                when pause_setI2273 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 292;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"2";
                  state_var3002 <= pause_setI2272;
                when pause_setI2274 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 291;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2273;
                when pause_setI2275 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 290;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"2c";
                  state_var3002 <= pause_setI2274;
                when pause_setI2276 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 289;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"14";
                  state_var3002 <= pause_setI2275;
                when pause_setI2277 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 288;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"36";
                  state_var3002 <= pause_setI2276;
                when pause_setI2278 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 287;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"a";
                  state_var3002 <= pause_setI2277;
                when pause_setI2279 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 286;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"00000" & X"17");
                  state_var3002 <= pause_setI2278;
                when pause_setI2280 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 285;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"3";
                  state_var3002 <= pause_setI2279;
                when pause_setI2281 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 284;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"2b";
                  state_var3002 <= pause_setI2280;
                when pause_setI2282 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 283;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"13";
                  state_var3002 <= pause_setI2281;
                when pause_setI2283 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 282;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"36";
                  state_var3002 <= pause_setI2282;
                when pause_setI2284 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 281;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"12";
                  state_var3002 <= pause_setI2283;
                when pause_setI2285 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 280;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"36";
                  state_var3002 <= pause_setI2284;
                when pause_setI2286 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 279;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"a";
                  state_var3002 <= pause_setI2285;
                when pause_setI2287 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 278;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"21";
                  state_var3002 <= pause_setI2286;
                when pause_setI2288 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 277;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"11";
                  state_var3002 <= pause_setI2287;
                when pause_setI2289 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 276;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"36";
                  state_var3002 <= pause_setI2288;
                when pause_setI2290 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 275;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2289;
                when pause_setI2291 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 274;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"3";
                  state_var3002 <= pause_setI2290;
                when pause_setI2292 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 273;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"26";
                  state_var3002 <= pause_setI2291;
                when pause_setI2293 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 272;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"10";
                  state_var3002 <= pause_setI2292;
                when pause_setI2294 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 271;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"36";
                  state_var3002 <= pause_setI2293;
                when pause_setI2295 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 270;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"1c";
                  state_var3002 <= pause_setI2294;
                when pause_setI2296 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 269;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"22";
                  state_var3002 <= pause_setI2295;
                when pause_setI2297 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 268;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"1b";
                  state_var3002 <= pause_setI2296;
                when pause_setI2298 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 267;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"000000" & X"a");
                  state_var3002 <= pause_setI2297;
                when pause_setI2299 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 266;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2298;
                when pause_setI2300 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 265;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"2b";
                  state_var3002 <= pause_setI2299;
                when pause_setI2301 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 264;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"b";
                  state_var3002 <= pause_setI2300;
                when pause_setI2302 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 263;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"18";
                  state_var3002 <= pause_setI2301;
                when pause_setI2303 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 262;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2302;
                when pause_setI2304 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 261;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"28";
                  state_var3002 <= pause_setI2303;
                when pause_setI2305 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 260;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2304;
                when pause_setI2306 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 259;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"40";
                  state_var3002 <= pause_setI2305;
                when pause_setI2307 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 258;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"b";
                  state_var3002 <= pause_setI2306;
                when pause_setI2308 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 257;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"16";
                  state_var3002 <= pause_setI2307;
                when pause_setI2309 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 256;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2308;
                when pause_setI2310 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 255;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"28";
                  state_var3002 <= pause_setI2309;
                when pause_setI2311 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 254;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"f";
                  state_var3002 <= pause_setI2310;
                when pause_setI2312 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 253;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"35";
                  state_var3002 <= pause_setI2311;
                when pause_setI2313 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 252;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"3";
                  state_var3002 <= pause_setI2312;
                when pause_setI2314 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 251;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"26";
                  state_var3002 <= pause_setI2313;
                when pause_setI2315 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 250;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"1b";
                  state_var3002 <= pause_setI2314;
                when pause_setI2316 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 249;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"1c";
                  state_var3002 <= pause_setI2315;
                when pause_setI2317 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 248;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"21";
                  state_var3002 <= pause_setI2316;
                when pause_setI2318 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 247;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"32";
                  state_var3002 <= pause_setI2317;
                when pause_setI2319 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 246;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"000000" & X"1");
                  state_var3002 <= pause_setI2318;
                when pause_setI2320 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 245;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"7f";
                  state_var3002 <= pause_setI2319;
                when pause_setI2321 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 244;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2320;
                when pause_setI2322 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 243;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"a";
                  state_var3002 <= pause_setI2321;
                when pause_setI2323 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 242;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2322;
                when pause_setI2324 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 241;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"83";
                  state_var3002 <= pause_setI2323;
                when pause_setI2325 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 240;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2324;
                when pause_setI2326 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 239;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"3";
                  state_var3002 <= pause_setI2325;
                when pause_setI2327 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 238;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"28";
                  state_var3002 <= pause_setI2326;
                when pause_setI2328 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 237;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"64";
                  state_var3002 <= pause_setI2327;
                when pause_setI2329 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 236;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"4";
                  state_var3002 <= pause_setI2328;
                when pause_setI2330 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 235;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"28";
                  state_var3002 <= pause_setI2329;
                when pause_setI2331 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 234;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"7";
                  state_var3002 <= pause_setI2330;
                when pause_setI2332 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 233;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"27";
                  state_var3002 <= pause_setI2331;
                when pause_setI2333 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 232;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"32";
                  state_var3002 <= pause_setI2332;
                when pause_setI2334 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 231;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2333;
                when pause_setI2335 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 230;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"7f";
                  state_var3002 <= pause_setI2334;
                when pause_setI2336 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 229;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"d";
                  state_var3002 <= pause_setI2335;
                when pause_setI2337 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 228;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"d";
                  state_var3002 <= pause_setI2336;
                when pause_setI2338 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 227;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"44";
                  state_var3002 <= pause_setI2337;
                when pause_setI2339 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 226;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"3";
                  state_var3002 <= pause_setI2338;
                when pause_setI2340 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 225;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"a";
                  state_var3002 <= pause_setI2339;
                when pause_setI2341 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 224;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"56";
                  state_var3002 <= pause_setI2340;
                when pause_setI2342 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 223;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"58";
                  state_var3002 <= pause_setI2341;
                when pause_setI2343 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 222;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"79";
                  state_var3002 <= pause_setI2342;
                when pause_setI2344 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 221;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"d";
                  state_var3002 <= pause_setI2343;
                when pause_setI2345 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 220;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"6f";
                  state_var3002 <= pause_setI2344;
                when pause_setI2346 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 219;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"b";
                  state_var3002 <= pause_setI2345;
                when pause_setI2347 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 218;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2346;
                when pause_setI2348 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 217;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"12";
                  state_var3002 <= pause_setI2347;
                when pause_setI2349 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 216;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"56";
                  state_var3002 <= pause_setI2348;
                when pause_setI2350 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 215;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"58";
                  state_var3002 <= pause_setI2349;
                when pause_setI2351 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 214;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"79";
                  state_var3002 <= pause_setI2350;
                when pause_setI2352 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 213;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"d";
                  state_var3002 <= pause_setI2351;
                when pause_setI2353 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 212;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"6e";
                  state_var3002 <= pause_setI2352;
                when pause_setI2354 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 211;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"b";
                  state_var3002 <= pause_setI2353;
                when pause_setI2355 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 210;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2354;
                when pause_setI2356 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 209;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"1a";
                  state_var3002 <= pause_setI2355;
                when pause_setI2357 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 208;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"56";
                  state_var3002 <= pause_setI2356;
                when pause_setI2358 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 207;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"58";
                  state_var3002 <= pause_setI2357;
                when pause_setI2359 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 206;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"79";
                  state_var3002 <= pause_setI2358;
                when pause_setI2360 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 205;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"d";
                  state_var3002 <= pause_setI2359;
                when pause_setI2361 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 204;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"a";
                  state_var3002 <= pause_setI2360;
                when pause_setI2362 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 203;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"43";
                  state_var3002 <= pause_setI2361;
                when pause_setI2363 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 202;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"2";
                  state_var3002 <= pause_setI2362;
                when pause_setI2364 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 201;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"24";
                  state_var3002 <= pause_setI2363;
                when pause_setI2365 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 200;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"56";
                  state_var3002 <= pause_setI2364;
                when pause_setI2366 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 199;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"2";
                  state_var3002 <= pause_setI2365;
                when pause_setI2367 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 198;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"2";
                  state_var3002 <= pause_setI2366;
                when pause_setI2368 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 197;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"2a";
                  state_var3002 <= pause_setI2367;
                when pause_setI2369 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 196;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"29";
                  state_var3002 <= pause_setI2368;
                when pause_setI2370 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 195;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"2";
                  state_var3002 <= pause_setI2369;
                when pause_setI2371 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 194;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"28";
                  state_var3002 <= pause_setI2370;
                when pause_setI2372 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 193;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"4";
                  state_var3002 <= pause_setI2371;
                when pause_setI2373 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 192;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"26";
                  state_var3002 <= pause_setI2372;
                when pause_setI2374 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 191;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"e";
                  state_var3002 <= pause_setI2373;
                when pause_setI2375 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 190;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"36";
                  state_var3002 <= pause_setI2374;
                when pause_setI2376 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 189;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"21";
                  state_var3002 <= pause_setI2375;
                when pause_setI2377 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 188;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"c";
                  state_var3002 <= pause_setI2376;
                when pause_setI2378 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 187;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"43";
                  state_var3002 <= pause_setI2377;
                when pause_setI2379 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 186;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"c";
                  state_var3002 <= pause_setI2378;
                when pause_setI2380 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 185;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"22";
                  state_var3002 <= pause_setI2379;
                when pause_setI2381 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 184;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"32";
                  state_var3002 <= pause_setI2380;
                when pause_setI2382 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 183;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"b";
                  state_var3002 <= pause_setI2381;
                when pause_setI2383 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 182;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"44";
                  state_var3002 <= pause_setI2382;
                when pause_setI2384 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 181;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2383;
                when pause_setI2385 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 180;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"e";
                  state_var3002 <= pause_setI2384;
                when pause_setI2386 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 179;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"56";
                  state_var3002 <= pause_setI2385;
                when pause_setI2387 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 178;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2386;
                when pause_setI2388 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 177;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2387;
                when pause_setI2389 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 176;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"2a";
                  state_var3002 <= pause_setI2388;
                when pause_setI2390 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 175;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"29";
                  state_var3002 <= pause_setI2389;
                when pause_setI2391 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 174;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"2";
                  state_var3002 <= pause_setI2390;
                when pause_setI2392 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 173;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"28";
                  state_var3002 <= pause_setI2391;
                when pause_setI2393 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 172;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2392;
                when pause_setI2394 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 171;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"40";
                  state_var3002 <= pause_setI2393;
                when pause_setI2395 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 170;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"b";
                  state_var3002 <= pause_setI2394;
                when pause_setI2396 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 169;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"22";
                  state_var3002 <= pause_setI2395;
                when pause_setI2397 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 168;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"32";
                  state_var3002 <= pause_setI2396;
                when pause_setI2398 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 167;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2397;
                when pause_setI2399 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 166;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"7f";
                  state_var3002 <= pause_setI2398;
                when pause_setI2400 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 165;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"b";
                  state_var3002 <= pause_setI2399;
                when pause_setI2401 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 164;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2400;
                when pause_setI2402 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 163;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"2";
                  state_var3002 <= pause_setI2401;
                when pause_setI2403 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 162;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"28";
                  state_var3002 <= pause_setI2402;
                when pause_setI2404 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 161;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"63";
                  state_var3002 <= pause_setI2403;
                when pause_setI2405 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 160;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"4";
                  state_var3002 <= pause_setI2404;
                when pause_setI2406 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 159;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"56";
                  state_var3002 <= pause_setI2405;
                when pause_setI2407 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 158;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"7d";
                  state_var3002 <= pause_setI2406;
                when pause_setI2408 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 157;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"b";
                  state_var3002 <= pause_setI2407;
                when pause_setI2409 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 156;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2408;
                when pause_setI2410 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 155;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2409;
                when pause_setI2411 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 154;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"2a";
                  state_var3002 <= pause_setI2410;
                when pause_setI2412 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 153;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"29";
                  state_var3002 <= pause_setI2411;
                when pause_setI2413 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 152;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"ce";
                  state_var3002 <= pause_setI2412;
                when pause_setI2414 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 151;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"54";
                  state_var3002 <= pause_setI2413;
                when pause_setI2415 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 150;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"10";
                  state_var3002 <= pause_setI2414;
                when pause_setI2416 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 149;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"39";
                  state_var3002 <= pause_setI2415;
                when pause_setI2417 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 148;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"00000" & X"41");
                  state_var3002 <= pause_setI2416;
                when pause_setI2418 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 147;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2417;
                when pause_setI2419 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 146;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"2b";
                  state_var3002 <= pause_setI2418;
                when pause_setI2420 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 145;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"15";
                  state_var3002 <= pause_setI2419;
                when pause_setI2421 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 144;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"39";
                  state_var3002 <= pause_setI2420;
                when pause_setI2422 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 143;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"00000" & X"1d");
                  state_var3002 <= pause_setI2421;
                when pause_setI2423 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 142;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2422;
                when pause_setI2424 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 141;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"2b";
                  state_var3002 <= pause_setI2423;
                when pause_setI2425 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 140;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"c";
                  state_var3002 <= pause_setI2424;
                when pause_setI2426 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 139;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"39";
                  state_var3002 <= pause_setI2425;
                when pause_setI2427 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 138;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"000000" & X"f");
                  state_var3002 <= pause_setI2426;
                when pause_setI2428 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 137;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2427;
                when pause_setI2429 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 136;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"2b";
                  state_var3002 <= pause_setI2428;
                when pause_setI2430 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 135;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"d";
                  state_var3002 <= pause_setI2429;
                when pause_setI2431 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 134;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"39";
                  state_var3002 <= pause_setI2430;
                when pause_setI2432 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 133;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2431;
                when pause_setI2433 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 132;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"00000" & X"64");
                  state_var3002 <= pause_setI2432;
                when pause_setI2434 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 131;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2433;
                when pause_setI2435 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 130;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2434;
                when pause_setI2436 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 129;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"2c";
                  state_var3002 <= pause_setI2435;
                when pause_setI2437 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 128;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"3";
                  state_var3002 <= pause_setI2436;
                when pause_setI2438 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 127;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"26";
                  state_var3002 <= pause_setI2437;
                when pause_setI2439 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 126;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"d";
                  state_var3002 <= pause_setI2438;
                when pause_setI2440 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 125;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"36";
                  state_var3002 <= pause_setI2439;
                when pause_setI2441 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 124;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"b";
                  state_var3002 <= pause_setI2440;
                when pause_setI2442 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 123;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"63";
                  state_var3002 <= pause_setI2441;
                when pause_setI2443 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 122;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"4";
                  state_var3002 <= pause_setI2442;
                when pause_setI2444 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 121;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"26";
                  state_var3002 <= pause_setI2443;
                when pause_setI2445 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 120;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"c";
                  state_var3002 <= pause_setI2444;
                when pause_setI2446 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 119;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"c";
                  state_var3002 <= pause_setI2445;
                when pause_setI2447 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 118;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"63";
                  state_var3002 <= pause_setI2446;
                when pause_setI2448 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 117;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"00000" & X"13");
                  state_var3002 <= pause_setI2447;
                when pause_setI2449 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 116;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2448;
                when pause_setI2450 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 115;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2449;
                when pause_setI2451 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 114;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"2c";
                  state_var3002 <= pause_setI2450;
                when pause_setI2452 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 113;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"2";
                  state_var3002 <= pause_setI2451;
                when pause_setI2453 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 112;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"28";
                  state_var3002 <= pause_setI2452;
                when pause_setI2454 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 111;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2453;
                when pause_setI2455 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 110;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"4";
                  state_var3002 <= pause_setI2454;
                when pause_setI2456 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 109;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"26";
                  state_var3002 <= pause_setI2455;
                when pause_setI2457 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 108;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"32";
                  state_var3002 <= pause_setI2456;
                when pause_setI2458 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 107;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"44";
                  state_var3002 <= pause_setI2457;
                when pause_setI2459 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 106;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"b";
                  state_var3002 <= pause_setI2458;
                when pause_setI2460 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 105;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2459;
                when pause_setI2461 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 104;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"7f";
                  state_var3002 <= pause_setI2460;
                when pause_setI2462 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 103;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2461;
                when pause_setI2463 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 102;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"9";
                  state_var3002 <= pause_setI2462;
                when pause_setI2464 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 101;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"56";
                  state_var3002 <= pause_setI2463;
                when pause_setI2465 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 100;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2464;
                when pause_setI2466 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 99;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2465;
                when pause_setI2467 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 98;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"2a";
                  state_var3002 <= pause_setI2466;
                when pause_setI2468 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 97;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"29";
                  state_var3002 <= pause_setI2467;
                when pause_setI2469 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 96;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"5";
                  state_var3002 <= pause_setI2468;
                when pause_setI2470 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 95;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"26";
                  state_var3002 <= pause_setI2469;
                when pause_setI2471 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 94;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"c";
                  state_var3002 <= pause_setI2470;
                when pause_setI2472 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 93;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"d";
                  state_var3002 <= pause_setI2471;
                when pause_setI2473 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 92;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"63";
                  state_var3002 <= pause_setI2472;
                when pause_setI2474 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 91;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"00000" & X"28");
                  state_var3002 <= pause_setI2473;
                when pause_setI2475 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 90;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"2";
                  state_var3002 <= pause_setI2474;
                when pause_setI2476 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 89;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2475;
                when pause_setI2477 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 88;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"2c";
                  state_var3002 <= pause_setI2476;
                when pause_setI2478 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 87;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"c";
                  state_var3002 <= pause_setI2477;
                when pause_setI2479 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 86;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"36";
                  state_var3002 <= pause_setI2478;
                when pause_setI2480 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 85;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2479;
                when pause_setI2481 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 84;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2480;
                when pause_setI2482 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 83;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"2a";
                  state_var3002 <= pause_setI2481;
                when pause_setI2483 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 82;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"29";
                  state_var3002 <= pause_setI2482;
                when pause_setI2484 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 81;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"3";
                  state_var3002 <= pause_setI2483;
                when pause_setI2485 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 80;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"25";
                  state_var3002 <= pause_setI2484;
                when pause_setI2486 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 79;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"1b";
                  state_var3002 <= pause_setI2485;
                when pause_setI2487 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 78;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2486;
                when pause_setI2488 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 77;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"6";
                  state_var3002 <= pause_setI2487;
                when pause_setI2489 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 76;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"26";
                  state_var3002 <= pause_setI2488;
                when pause_setI2490 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 75;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"32";
                  state_var3002 <= pause_setI2489;
                when pause_setI2491 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 74;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"c";
                  state_var3002 <= pause_setI2490;
                when pause_setI2492 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 73;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"3";
                  state_var3002 <= pause_setI2491;
                when pause_setI2493 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 72;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"6";
                  state_var3002 <= pause_setI2492;
                when pause_setI2494 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 71;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"26";
                  state_var3002 <= pause_setI2493;
                when pause_setI2495 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 70;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"32";
                  state_var3002 <= pause_setI2494;
                when pause_setI2496 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 69;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"c";
                  state_var3002 <= pause_setI2495;
                when pause_setI2497 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 68;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2496;
                when pause_setI2498 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 67;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"40";
                  state_var3002 <= pause_setI2497;
                when pause_setI2499 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 66;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"b";
                  state_var3002 <= pause_setI2498;
                when pause_setI2500 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 65;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"3";
                  state_var3002 <= pause_setI2499;
                when pause_setI2501 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 64;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"9";
                  state_var3002 <= pause_setI2500;
                when pause_setI2502 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 63;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"56";
                  state_var3002 <= pause_setI2501;
                when pause_setI2503 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 62;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"21";
                  state_var3002 <= pause_setI2502;
                when pause_setI2504 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 61;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"1c";
                  state_var3002 <= pause_setI2503;
                when pause_setI2505 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 60;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"a";
                  state_var3002 <= pause_setI2504;
                when pause_setI2506 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 59;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"43";
                  state_var3002 <= pause_setI2505;
                when pause_setI2507 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 58;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"b";
                  state_var3002 <= pause_setI2506;
                when pause_setI2508 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 57;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"44";
                  state_var3002 <= pause_setI2507;
                when pause_setI2509 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 56;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2508;
                when pause_setI2510 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 55;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"17";
                  state_var3002 <= pause_setI2509;
                when pause_setI2511 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 54;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"56";
                  state_var3002 <= pause_setI2510;
                when pause_setI2512 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 53;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2511;
                when pause_setI2513 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 52;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2512;
                when pause_setI2514 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 51;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"2a";
                  state_var3002 <= pause_setI2513;
                when pause_setI2515 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 50;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"29";
                  state_var3002 <= pause_setI2514;
                when pause_setI2516 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 49;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"2";
                  state_var3002 <= pause_setI2515;
                when pause_setI2517 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 48;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"28";
                  state_var3002 <= pause_setI2516;
                when pause_setI2518 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 47;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2517;
                when pause_setI2519 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 46;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"4";
                  state_var3002 <= pause_setI2518;
                when pause_setI2520 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 45;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"26";
                  state_var3002 <= pause_setI2519;
                when pause_setI2521 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 44;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"32";
                  state_var3002 <= pause_setI2520;
                when pause_setI2522 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 43;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"44";
                  state_var3002 <= pause_setI2521;
                when pause_setI2523 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 42;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"b";
                  state_var3002 <= pause_setI2522;
                when pause_setI2524 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 41;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2523;
                when pause_setI2525 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 40;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"40";
                  state_var3002 <= pause_setI2524;
                when pause_setI2526 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 39;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"43";
                  state_var3002 <= pause_setI2525;
                when pause_setI2527 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 38;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"b";
                  state_var3002 <= pause_setI2526;
                when pause_setI2528 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 37;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2527;
                when pause_setI2529 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 36;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"b";
                  state_var3002 <= pause_setI2528;
                when pause_setI2530 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 35;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"56";
                  state_var3002 <= pause_setI2529;
                when pause_setI2531 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 34;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2530;
                when pause_setI2532 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 33;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2531;
                when pause_setI2533 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 32;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"2a";
                  state_var3002 <= pause_setI2532;
                when pause_setI2534 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 31;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"29";
                  state_var3002 <= pause_setI2533;
                when pause_setI2535 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 30;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"63";
                  state_var3002 <= pause_setI2534;
                when pause_setI2536 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 29;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"54";
                  state_var3002 <= pause_setI2535;
                when pause_setI2537 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 28;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"e";
                  state_var3002 <= pause_setI2536;
                when pause_setI2538 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 27;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"39";
                  state_var3002 <= pause_setI2537;
                when pause_setI2539 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 26;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2538;
                when pause_setI2540 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 25;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"00000" & X"16");
                  state_var3002 <= pause_setI2539;
                when pause_setI2541 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 24;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2540;
                when pause_setI2542 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 23;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2541;
                when pause_setI2543 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 22;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"2c";
                  state_var3002 <= pause_setI2542;
                when pause_setI2544 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 21;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"2";
                  state_var3002 <= pause_setI2543;
                when pause_setI2545 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 20;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"28";
                  state_var3002 <= pause_setI2544;
                when pause_setI2546 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 19;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2545;
                when pause_setI2547 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 18;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"2";
                  state_var3002 <= pause_setI2546;
                when pause_setI2548 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 17;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"28";
                  state_var3002 <= pause_setI2547;
                when pause_setI2549 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 16;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2548;
                when pause_setI2550 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 15;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"40";
                  state_var3002 <= pause_setI2549;
                when pause_setI2551 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 14;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"43";
                  state_var3002 <= pause_setI2550;
                when pause_setI2552 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 13;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"b";
                  state_var3002 <= pause_setI2551;
                when pause_setI2553 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 12;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"22";
                  state_var3002 <= pause_setI2552;
                when pause_setI2554 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 11;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"32";
                  state_var3002 <= pause_setI2553;
                when pause_setI2555 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 10;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"44";
                  state_var3002 <= pause_setI2554;
                when pause_setI2556 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 9;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"b";
                  state_var3002 <= pause_setI2555;
                when pause_setI2557 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 8;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2556;
                when pause_setI2558 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 7;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"c";
                  state_var3002 <= pause_setI2557;
                when pause_setI2559 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 6;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"56";
                  state_var3002 <= pause_setI2558;
                when pause_setI2560 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 5;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"0";
                  state_var3002 <= pause_setI2559;
                when pause_setI2561 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 4;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"000000" & X"1";
                  state_var3002 <= pause_setI2560;
                when pause_setI2562 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 3;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"2a";
                  state_var3002 <= pause_setI2561;
                when pause_setI2563 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 2;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"29";
                  state_var3002 <= pause_setI2562;
                when pause_setI2564 =>
                  \$code_write_request\ <= '0';
                  \$code_ptr_write\ <= 1;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"15";
                  state_var3002 <= pause_setI2563;
                when pause_setI2565 =>
                  \$global_end_write_request\ <= '0';
                  \$code_ptr_write\ <= 0;
                  \$code_write_request\ <= '1';
                  \$code_write\ <= "000"& X"00000" & X"54";
                  state_var3002 <= pause_setI2564;
                when pause_setI2566 =>
                  \$ram_write_request\ <= '0';
                  \$global_end_ptr_write\ <= 0;
                  \$global_end_write_request\ <= '1';
                  \$global_end_write\ <= eclat_add(X"3e80" & X"00" & X"17");
                  state_var3002 <= pause_setI2565;
                when pause_setI2567 =>
                  \$ram_write_request\ <= '0';
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(X"3e80" & X"00" & X"16")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= "000"& X"000000" & X"0" & eclat_true;
                  state_var3002 <= pause_setI2566;
                when pause_setI2568 =>
                  \$ram_write_request\ <= '0';
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(X"3e80" & X"00" & X"15")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= "000"& X"000000" & X"0" & eclat_true;
                  state_var3002 <= pause_setI2567;
                when pause_setI2569 =>
                  \$ram_write_request\ <= '0';
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(X"3e80" & X"00" & X"14")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= "000"& X"000000" & X"0" & eclat_true;
                  state_var3002 <= pause_setI2568;
                when pause_setI2570 =>
                  \$ram_write_request\ <= '0';
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(X"3e80" & X"00" & X"13")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= "000"& X"000000" & X"0" & eclat_true;
                  state_var3002 <= pause_setI2569;
                when pause_setI2571 =>
                  \$ram_write_request\ <= '0';
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(X"3e80" & X"00" & X"12")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= "000"& X"000000" & X"0" & eclat_true;
                  state_var3002 <= pause_setI2570;
                when pause_setI2572 =>
                  \$ram_write_request\ <= '0';
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(X"3e80" & X"00" & X"11")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= "000"& X"000000" & X"0" & eclat_true;
                  state_var3002 <= pause_setI2571;
                when pause_setI2573 =>
                  \$ram_write_request\ <= '0';
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(X"3e80" & X"00" & X"10")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= "000"& X"000000" & X"0" & eclat_true;
                  state_var3002 <= pause_setI2572;
                when pause_setI2574 =>
                  \$ram_write_request\ <= '0';
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(X"3e80" & X"000" & X"f")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= eclat_resize(X"3e80",31) & eclat_false;
                  state_var3002 <= pause_setI2573;
                when pause_setI2575 =>
                  \$ram_write_request\ <= '0';
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(X"3e80" & X"000" & X"2")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= "000"& X"000000" & X"0" & eclat_true;
                  state_var3002 <= pause_setI2574;
                when pause_setI2576 =>
                  \$ram_write_request\ <= '0';
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(X"3e80" & X"000" & X"1")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= "000"& X"000000" & X"0" & eclat_true;
                  state_var3002 <= pause_setI2575;
                when pause_setI2577 =>
                  \$ram_write_request\ <= '0';
                  \$ram_ptr_write\ <= 16000;
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= eclat_lor(eclat_lsl(eclat_resize(X"0" & X"0",31) & "000"& X"00000" & X"18") & eclat_lsl(eclat_resize(X"000" & X"2",31) & "000"& X"000000" & X"2")) & eclat_true;
                  state_var3002 <= pause_setI2576;
                when pause_setI2578 =>
                  \$ram_write_request\ <= '0';
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(X"3e80" & X"000" & X"e")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= "000"& X"000000" & X"0" & eclat_true;
                  state_var3002 <= pause_setI2577;
                when pause_setI2579 =>
                  \$ram_write_request\ <= '0';
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(X"3e80" & X"000" & X"d")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= "000"& X"000000" & X"0" & eclat_true;
                  state_var3002 <= pause_setI2578;
                when compute2140 =>
                  rdy2139 := eclat_false;
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(X"3e80" & X"000" & X"c")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= "000"& X"000000" & X"0" & eclat_true;
                  state_var3002 <= pause_setI2579;
                end case;
                \$v2581\ := eclat_not(rdy2139);
                if \$v2581\(0) = '1' then
                  result2138 := eclat_unit;
                end if;
                \$v932\ := result2138 & rdy2139;
                \$v2137\ := eclat_not(\$v934_init_done\);
                if \$v2137\(0) = '1' then
                  \$v934\ := eclat_false;
                  \$v934_init_done\ := eclat_true;
                end if;
                \$v934\ := eclat_and(eclat_if(\$v934\ & eclat_true & ""&\$v932\(1)) & eclat_not(eclat_false));
                \$12_rdy\ := \$v934\;
                \$v516\ := eclat_false & eclat_true & \$12_rdy\ & ""&\$v516\(3);
              else
                \$v2995\ := eclat_not(\$v522_init_done\);
                if \$v2995\(0) = '1' then
                  \$v522\ := X"000" & X"0" & "000"& X"000000" & X"1" & eclat_true & X"0" & X"3e8" & "000"& X"000000" & X"1" & eclat_true & X"0" & X"0" & X"000" & X"0" & eclat_false & eclat_false & eclat_true;
                  \$v522_init_done\ := eclat_true;
                end if;
                \$v2994\ := eclat_not(""&\$v516\(2));
                if \$v2994\(0) = '1' then
                  \$v522\ := \$v522\(0 to 121) & eclat_true;
                else
                  case state_var3000 is
                  when \$103_w\ =>
                    \$v2858\ := eclat_gt(\$103_w_arg\(0 to 7) & \$103_w_arg\(56 to 63));
                    if \$v2858\(0) = '1' then
                      \$103_w_result\ := \$103_w_arg\(8 to 23);
                      \$104_sp\ := \$103_w_result\;
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$104_sp\ & X"000" & X"1")));
                      state_var3000 <= pause_getI2863;
                    else
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$103_w_arg\(8 to 23) & X"000" & X"1")));
                      state_var3000 <= pause_getI2856;
                    end if;
                  when \$1278_forever\ =>
                    state_var3000 <= \$1278_forever\;
                  when \$1281_forever\ =>
                    state_var3000 <= \$1281_forever\;
                  when \$1284_forever\ =>
                    state_var3000 <= \$1284_forever\;
                  when \$1342_modulo\ =>
                    \$v2684\ := eclat_lt(\$1342_modulo_arg\(0 to 30) & \$1342_modulo_arg\(31 to 61));
                    if \$v2684\(0) = '1' then
                      \$1342_modulo_result\ := \$1342_modulo_arg\(0 to 30);
                      \$1343_r\ := \$1342_modulo_result\;
                      \$313_res\ := eclat_if(eclat_lt(binop_int_arg(48 to 78) & "000"& X"000000" & X"0") & eclat_sub("000"& X"000000" & X"0" & \$1343_r\) & \$1343_r\);
                      binop_int_result := eclat_add(binop_int_arg(32 to 47) & X"000" & X"1") & \$313_res\ & eclat_true & \$v886\(32 to 47) & binop_int_arg(96 to 151) & binop_int_arg(152 to 153);
                      result2582 := binop_int_result;
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    else
                      \$1342_modulo_arg\ := eclat_sub(\$1342_modulo_arg\(0 to 30) & \$1342_modulo_arg\(31 to 61)) & \$1342_modulo_arg\(31 to 61);
                      state_var3000 <= \$1342_modulo\;
                    end if;
                  when \$74_fill\ =>
                    \$v2959\ := eclat_ge(\$74_fill_arg\(0 to 15) & \$74_fill_arg\(64 to 79));
                    if \$v2959\(0) = '1' then
                      \$74_fill_result\ := \$74_fill_arg\(16 to 31);
                      \$75_sp\ := \$74_fill_result\;
                      result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"3") & \$v593\(64 to 95) & \$75_sp\ & \$v593\(32 to 63) & \$v522\(96 to 103) & \$v522\(104 to 119) & \$v522\(120 to 121);
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    else
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$74_fill_arg\(16 to 31) & X"000" & X"1")));
                      state_var3000 <= pause_getI2957;
                    end if;
                  when \$855_forever\ =>
                    state_var3000 <= \$855_forever\;
                  when \$921_forever\ =>
                    state_var3000 <= \$921_forever\;
                  when apply =>
                    eclat_print_string(of_string("ENV:"));
                    
                    eclat_print_int(apply_arg(108 to 138));
                    
                    eclat_print_string(of_string("<"));
                    
                    \$v2681\ := ""&apply_arg(139);
                    if \$v2681\(0) = '1' then
                      eclat_print_string(of_string("int"));
                      
                      eclat_print_string(of_string(">"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$v2680\ := ""&apply_arg(0);
                      if \$v2680\(0) = '1' then
                        \$ram_ptr\ <= to_integer(unsigned(eclat_sub(apply_arg(92 to 107) & X"000" & X"1")));
                        state_var3000 <= pause_getI2678;
                      else
                        \$v906\ := "000"& X"000000" & X"1" & eclat_true & apply_arg(92 to 107);
                        \$v2677\ := ""&apply_arg(1);
                        if \$v2677\(0) = '1' then
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v906\(32 to 47) & X"000" & X"1")));
                          state_var3000 <= pause_getI2675;
                        else
                          \$v907\ := "000"& X"000000" & X"1" & eclat_true & \$v906\(32 to 47);
                          \$v2674\ := ""&apply_arg(2);
                          if \$v2674\(0) = '1' then
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v907\(32 to 47) & X"000" & X"1")));
                            state_var3000 <= pause_getI2672;
                          else
                            \$v908\ := "000"& X"000000" & X"1" & eclat_true & \$v907\(32 to 47);
                            \$v2671\ := ""&apply_arg(11);
                            if \$v2671\(0) = '1' then
                              \$339_sp\ := eclat_add(eclat_sub(\$v908\(32 to 47) & apply_arg(12 to 27)) & apply_arg(28 to 43));
                              \$v2667\ := ""&apply_arg(2);
                              if \$v2667\(0) = '1' then
                                \$ram_ptr_write\ <= to_integer(unsigned(\$339_sp\));
                                \$ram_write_request\ <= '1';
                                \$ram_write\ <= \$v908\(0 to 31);
                                state_var3000 <= pause_setI2666;
                              else
                                \$340_sp\ := \$339_sp\;
                                \$v2665\ := ""&apply_arg(1);
                                if \$v2665\(0) = '1' then
                                  \$ram_ptr_write\ <= to_integer(unsigned(\$340_sp\));
                                  \$ram_write_request\ <= '1';
                                  \$ram_write\ <= \$v907\(0 to 31);
                                  state_var3000 <= pause_setI2664;
                                else
                                  \$341_sp\ := \$340_sp\;
                                  \$v2663\ := ""&apply_arg(0);
                                  if \$v2663\(0) = '1' then
                                    \$ram_ptr_write\ <= to_integer(unsigned(\$341_sp\));
                                    \$ram_write_request\ <= '1';
                                    \$ram_write\ <= \$v906\(0 to 31);
                                    state_var3000 <= pause_setI2662;
                                  else
                                    \$342_sp\ := \$341_sp\;
                                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(apply_arg(60 to 90),16) & X"000" & X"0") & X"000" & X"1")));
                                    state_var3000 <= pause_getI2660;
                                  end if;
                                end if;
                              end if;
                            else
                              \$ram_ptr_write\ <= to_integer(unsigned(\$v908\(32 to 47)));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= eclat_resize(apply_arg(140 to 147),31) & eclat_true;
                              state_var3000 <= pause_setI2670;
                            end if;
                          end if;
                        end if;
                      end if;
                    else
                      eclat_print_string(of_string("ptr"));
                      
                      eclat_print_string(of_string(">"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$v2680\ := ""&apply_arg(0);
                      if \$v2680\(0) = '1' then
                        \$ram_ptr\ <= to_integer(unsigned(eclat_sub(apply_arg(92 to 107) & X"000" & X"1")));
                        state_var3000 <= pause_getI2678;
                      else
                        \$v906\ := "000"& X"000000" & X"1" & eclat_true & apply_arg(92 to 107);
                        \$v2677\ := ""&apply_arg(1);
                        if \$v2677\(0) = '1' then
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v906\(32 to 47) & X"000" & X"1")));
                          state_var3000 <= pause_getI2675;
                        else
                          \$v907\ := "000"& X"000000" & X"1" & eclat_true & \$v906\(32 to 47);
                          \$v2674\ := ""&apply_arg(2);
                          if \$v2674\(0) = '1' then
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v907\(32 to 47) & X"000" & X"1")));
                            state_var3000 <= pause_getI2672;
                          else
                            \$v908\ := "000"& X"000000" & X"1" & eclat_true & \$v907\(32 to 47);
                            \$v2671\ := ""&apply_arg(11);
                            if \$v2671\(0) = '1' then
                              \$339_sp\ := eclat_add(eclat_sub(\$v908\(32 to 47) & apply_arg(12 to 27)) & apply_arg(28 to 43));
                              \$v2667\ := ""&apply_arg(2);
                              if \$v2667\(0) = '1' then
                                \$ram_ptr_write\ <= to_integer(unsigned(\$339_sp\));
                                \$ram_write_request\ <= '1';
                                \$ram_write\ <= \$v908\(0 to 31);
                                state_var3000 <= pause_setI2666;
                              else
                                \$340_sp\ := \$339_sp\;
                                \$v2665\ := ""&apply_arg(1);
                                if \$v2665\(0) = '1' then
                                  \$ram_ptr_write\ <= to_integer(unsigned(\$340_sp\));
                                  \$ram_write_request\ <= '1';
                                  \$ram_write\ <= \$v907\(0 to 31);
                                  state_var3000 <= pause_setI2664;
                                else
                                  \$341_sp\ := \$340_sp\;
                                  \$v2663\ := ""&apply_arg(0);
                                  if \$v2663\(0) = '1' then
                                    \$ram_ptr_write\ <= to_integer(unsigned(\$341_sp\));
                                    \$ram_write_request\ <= '1';
                                    \$ram_write\ <= \$v906\(0 to 31);
                                    state_var3000 <= pause_setI2662;
                                  else
                                    \$342_sp\ := \$341_sp\;
                                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(apply_arg(60 to 90),16) & X"000" & X"0") & X"000" & X"1")));
                                    state_var3000 <= pause_getI2660;
                                  end if;
                                end if;
                              end if;
                            else
                              \$ram_ptr_write\ <= to_integer(unsigned(\$v908\(32 to 47)));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= eclat_resize(apply_arg(140 to 147),31) & eclat_true;
                              state_var3000 <= pause_setI2670;
                            end if;
                          end if;
                        end if;
                      end if;
                    end if;
                  when binop_compare =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(binop_compare_arg(80 to 95) & X"000" & X"1")));
                    state_var3000 <= pause_getI2690;
                  when binop_int =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(binop_int_arg(80 to 95) & X"000" & X"1")));
                    state_var3000 <= pause_getI2687;
                  when branch_if =>
                    \$v2704\ := eclat_if(""&branch_if_arg(0) & eclat_not(eclat_neq(branch_if_arg(17 to 47) & "000"& X"000000" & X"0")) & eclat_neq(branch_if_arg(17 to 47) & "000"& X"000000" & X"0"));
                    if \$v2704\(0) = '1' then
                      \$code_ptr\ <= to_integer(unsigned(eclat_add(branch_if_arg(1 to 16) & X"000" & X"1")));
                      state_var3000 <= pause_getI2702;
                    else
                      branch_if_result := eclat_add(branch_if_arg(1 to 16) & X"000" & X"2") & branch_if_arg(17 to 48) & branch_if_arg(49 to 64) & branch_if_arg(65 to 120) & branch_if_arg(121 to 122);
                      result2582 := branch_if_result;
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    end if;
                  when compare =>
                    \$v2689\ := compare_arg(0 to 31);
                    case \$v2689\ is
                    when X"0000000" & X"0" =>
                      compare_result := eclat_eq(compare_arg(32 to 62) & compare_arg(63 to 93));
                      case compare_id is
                      when X"00" & X"d" =>
                        \$300_res\ := compare_result;
                        binop_compare_result := eclat_add(binop_compare_arg(32 to 47) & X"000" & X"1") & 
                        eclat_if(\$300_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & \$v878\(32 to 47) & binop_compare_arg(96 to 151) & binop_compare_arg(152 to 153);
                        result2582 := binop_compare_result;
                        rdy2583 := eclat_true;
                        state_var3000 <= compute2584;
                      when X"0" & X"33" =>
                        \$233_b\ := compare_result;
                        compbranch_result := eclat_if(\$233_b\ & eclat_add(eclat_add(compbranch_arg(94 to 109) & X"000" & X"2") & eclat_resize(compbranch_arg(63 to 93),16)) & compbranch_arg(110 to 141) & compbranch_arg(142 to 157) & compbranch_arg(158 to 213) & compbranch_arg(214 to 215) & eclat_add(compbranch_arg(94 to 109) & X"000" & X"3") & compbranch_arg(110 to 141) & compbranch_arg(142 to 157) & compbranch_arg(158 to 213) & compbranch_arg(214 to 215));
                        result2582 := compbranch_result;
                        rdy2583 := eclat_true;
                        state_var3000 <= compute2584;
                      when others =>
                        
                      end case;
                    when X"0000000" & X"1" =>
                      compare_result := eclat_not(eclat_eq(compare_arg(32 to 62) & compare_arg(63 to 93)));
                      case compare_id is
                      when X"00" & X"d" =>
                        \$300_res\ := compare_result;
                        binop_compare_result := eclat_add(binop_compare_arg(32 to 47) & X"000" & X"1") & 
                        eclat_if(\$300_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & \$v878\(32 to 47) & binop_compare_arg(96 to 151) & binop_compare_arg(152 to 153);
                        result2582 := binop_compare_result;
                        rdy2583 := eclat_true;
                        state_var3000 <= compute2584;
                      when X"0" & X"33" =>
                        \$233_b\ := compare_result;
                        compbranch_result := eclat_if(\$233_b\ & eclat_add(eclat_add(compbranch_arg(94 to 109) & X"000" & X"2") & eclat_resize(compbranch_arg(63 to 93),16)) & compbranch_arg(110 to 141) & compbranch_arg(142 to 157) & compbranch_arg(158 to 213) & compbranch_arg(214 to 215) & eclat_add(compbranch_arg(94 to 109) & X"000" & X"3") & compbranch_arg(110 to 141) & compbranch_arg(142 to 157) & compbranch_arg(158 to 213) & compbranch_arg(214 to 215));
                        result2582 := compbranch_result;
                        rdy2583 := eclat_true;
                        state_var3000 <= compute2584;
                      when others =>
                        
                      end case;
                    when X"0000000" & X"2" =>
                      compare_result := eclat_lt(compare_arg(32 to 62) & compare_arg(63 to 93));
                      case compare_id is
                      when X"00" & X"d" =>
                        \$300_res\ := compare_result;
                        binop_compare_result := eclat_add(binop_compare_arg(32 to 47) & X"000" & X"1") & 
                        eclat_if(\$300_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & \$v878\(32 to 47) & binop_compare_arg(96 to 151) & binop_compare_arg(152 to 153);
                        result2582 := binop_compare_result;
                        rdy2583 := eclat_true;
                        state_var3000 <= compute2584;
                      when X"0" & X"33" =>
                        \$233_b\ := compare_result;
                        compbranch_result := eclat_if(\$233_b\ & eclat_add(eclat_add(compbranch_arg(94 to 109) & X"000" & X"2") & eclat_resize(compbranch_arg(63 to 93),16)) & compbranch_arg(110 to 141) & compbranch_arg(142 to 157) & compbranch_arg(158 to 213) & compbranch_arg(214 to 215) & eclat_add(compbranch_arg(94 to 109) & X"000" & X"3") & compbranch_arg(110 to 141) & compbranch_arg(142 to 157) & compbranch_arg(158 to 213) & compbranch_arg(214 to 215));
                        result2582 := compbranch_result;
                        rdy2583 := eclat_true;
                        state_var3000 <= compute2584;
                      when others =>
                        
                      end case;
                    when X"0000000" & X"3" =>
                      compare_result := eclat_if(eclat_lt(compare_arg(32 to 62) & compare_arg(63 to 93)) & eclat_true & eclat_eq(compare_arg(32 to 62) & compare_arg(63 to 93)));
                      case compare_id is
                      when X"00" & X"d" =>
                        \$300_res\ := compare_result;
                        binop_compare_result := eclat_add(binop_compare_arg(32 to 47) & X"000" & X"1") & 
                        eclat_if(\$300_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & \$v878\(32 to 47) & binop_compare_arg(96 to 151) & binop_compare_arg(152 to 153);
                        result2582 := binop_compare_result;
                        rdy2583 := eclat_true;
                        state_var3000 <= compute2584;
                      when X"0" & X"33" =>
                        \$233_b\ := compare_result;
                        compbranch_result := eclat_if(\$233_b\ & eclat_add(eclat_add(compbranch_arg(94 to 109) & X"000" & X"2") & eclat_resize(compbranch_arg(63 to 93),16)) & compbranch_arg(110 to 141) & compbranch_arg(142 to 157) & compbranch_arg(158 to 213) & compbranch_arg(214 to 215) & eclat_add(compbranch_arg(94 to 109) & X"000" & X"3") & compbranch_arg(110 to 141) & compbranch_arg(142 to 157) & compbranch_arg(158 to 213) & compbranch_arg(214 to 215));
                        result2582 := compbranch_result;
                        rdy2583 := eclat_true;
                        state_var3000 <= compute2584;
                      when others =>
                        
                      end case;
                    when X"0000000" & X"4" =>
                      compare_result := eclat_not(eclat_if(eclat_lt(compare_arg(32 to 62) & compare_arg(63 to 93)) & eclat_true & eclat_eq(compare_arg(32 to 62) & compare_arg(63 to 93))));
                      case compare_id is
                      when X"00" & X"d" =>
                        \$300_res\ := compare_result;
                        binop_compare_result := eclat_add(binop_compare_arg(32 to 47) & X"000" & X"1") & 
                        eclat_if(\$300_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & \$v878\(32 to 47) & binop_compare_arg(96 to 151) & binop_compare_arg(152 to 153);
                        result2582 := binop_compare_result;
                        rdy2583 := eclat_true;
                        state_var3000 <= compute2584;
                      when X"0" & X"33" =>
                        \$233_b\ := compare_result;
                        compbranch_result := eclat_if(\$233_b\ & eclat_add(eclat_add(compbranch_arg(94 to 109) & X"000" & X"2") & eclat_resize(compbranch_arg(63 to 93),16)) & compbranch_arg(110 to 141) & compbranch_arg(142 to 157) & compbranch_arg(158 to 213) & compbranch_arg(214 to 215) & eclat_add(compbranch_arg(94 to 109) & X"000" & X"3") & compbranch_arg(110 to 141) & compbranch_arg(142 to 157) & compbranch_arg(158 to 213) & compbranch_arg(214 to 215));
                        result2582 := compbranch_result;
                        rdy2583 := eclat_true;
                        state_var3000 <= compute2584;
                      when others =>
                        
                      end case;
                    when X"0000000" & X"5" =>
                      compare_result := eclat_not(eclat_lt(compare_arg(32 to 62) & compare_arg(63 to 93)));
                      case compare_id is
                      when X"00" & X"d" =>
                        \$300_res\ := compare_result;
                        binop_compare_result := eclat_add(binop_compare_arg(32 to 47) & X"000" & X"1") & 
                        eclat_if(\$300_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & \$v878\(32 to 47) & binop_compare_arg(96 to 151) & binop_compare_arg(152 to 153);
                        result2582 := binop_compare_result;
                        rdy2583 := eclat_true;
                        state_var3000 <= compute2584;
                      when X"0" & X"33" =>
                        \$233_b\ := compare_result;
                        compbranch_result := eclat_if(\$233_b\ & eclat_add(eclat_add(compbranch_arg(94 to 109) & X"000" & X"2") & eclat_resize(compbranch_arg(63 to 93),16)) & compbranch_arg(110 to 141) & compbranch_arg(142 to 157) & compbranch_arg(158 to 213) & compbranch_arg(214 to 215) & eclat_add(compbranch_arg(94 to 109) & X"000" & X"3") & compbranch_arg(110 to 141) & compbranch_arg(142 to 157) & compbranch_arg(158 to 213) & compbranch_arg(214 to 215));
                        result2582 := compbranch_result;
                        rdy2583 := eclat_true;
                        state_var3000 <= compute2584;
                      when others =>
                        
                      end case;
                    when others =>
                      compare_result := eclat_false;
                      case compare_id is
                      when X"00" & X"d" =>
                        \$300_res\ := compare_result;
                        binop_compare_result := eclat_add(binop_compare_arg(32 to 47) & X"000" & X"1") & 
                        eclat_if(\$300_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & \$v878\(32 to 47) & binop_compare_arg(96 to 151) & binop_compare_arg(152 to 153);
                        result2582 := binop_compare_result;
                        rdy2583 := eclat_true;
                        state_var3000 <= compute2584;
                      when X"0" & X"33" =>
                        \$233_b\ := compare_result;
                        compbranch_result := eclat_if(\$233_b\ & eclat_add(eclat_add(compbranch_arg(94 to 109) & X"000" & X"2") & eclat_resize(compbranch_arg(63 to 93),16)) & compbranch_arg(110 to 141) & compbranch_arg(142 to 157) & compbranch_arg(158 to 213) & compbranch_arg(214 to 215) & eclat_add(compbranch_arg(94 to 109) & X"000" & X"3") & compbranch_arg(110 to 141) & compbranch_arg(142 to 157) & compbranch_arg(158 to 213) & compbranch_arg(214 to 215));
                        result2582 := compbranch_result;
                        rdy2583 := eclat_true;
                        state_var3000 <= compute2584;
                      when others =>
                        
                      end case;
                    end case;
                  when compbranch =>
                    compare_id := X"0" & X"33";
                    compare_arg := compbranch_arg(0 to 31) & compbranch_arg(32 to 62) & compbranch_arg(110 to 140);
                    state_var3000 <= compare;
                  when fill =>
                    \$v2943\ := eclat_gt(fill_arg(0 to 15) & fill_arg(32 to 47));
                    if \$v2943\(0) = '1' then
                      fill_result := fill_arg(16 to 31);
                      \$59_sp\ := fill_result;
                      result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"3") & \$v576\(64 to 95) & \$59_sp\ & \$v576\(32 to 63) & \$v522\(96 to 103) & \$v522\(104 to 119) & \$v522\(120 to 121);
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    else
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(fill_arg(16 to 31) & X"000" & X"1")));
                      state_var3000 <= pause_getI2941;
                    end if;
                  when forever =>
                    state_var3000 <= forever;
                  when loop_push =>
                    \$v2767\ := eclat_ge(loop_push_arg(16 to 23) & eclat_sub(loop_push_arg(56 to 63) & X"0" & X"2"));
                    if \$v2767\(0) = '1' then
                      loop_push_result := loop_push_arg(0 to 15);
                      \$235_sp\ := loop_push_result;
                      \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v522\(64 to 94),16) & X"000" & X"1") & X"000" & X"1")));
                      state_var3000 <= pause_getI2768;
                    else
                      \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(loop_push_arg(24 to 54),16) & eclat_resize(eclat_add(loop_push_arg(16 to 23) & X"0" & X"2"),16)) & X"000" & X"1")));
                      state_var3000 <= pause_getI2765;
                    end if;
                  when make_block =>
                    eclat_print_string(of_string("GC-ALLOC:(size="));
                    
                    eclat_print_int(eclat_add(eclat_if(eclat_eq(make_block_arg(88 to 103) & X"000" & X"0") & X"000" & X"1" & make_block_arg(88 to 103)) & X"000" & X"1"));
                    
                    eclat_print_string(of_string(")"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    wait_arg := eclat_unit & make_block_arg(16 to 47) & make_block_arg(48 to 79) & make_block_arg(0 to 15) & eclat_add(
                    eclat_if(eclat_eq(make_block_arg(88 to 103) & X"000" & X"0") & X"000" & X"1" & make_block_arg(88 to 103)) & X"000" & X"1");
                    state_var3000 <= \wait\;
                  when make_block_n =>
                    make_block_id := X"00" & X"e";
                    make_block_arg := make_block_n_arg(16 to 31) & make_block_n_arg(82 to 113) & make_block_n_arg(114 to 145) & eclat_resize(make_block_n_arg(35 to 65),8) & make_block_n_arg(66 to 81);
                    state_var3000 <= make_block;
                  when modulo =>
                    \$v2682\ := eclat_lt(modulo_arg(0 to 30) & modulo_arg(31 to 61));
                    if \$v2682\(0) = '1' then
                      modulo_result := modulo_arg(0 to 30);
                      r := modulo_result;
                      \$313_res\ := eclat_if(eclat_lt(binop_int_arg(48 to 78) & "000"& X"000000" & X"0") & eclat_sub("000"& X"000000" & X"0" & r) & r);
                      binop_int_result := eclat_add(binop_int_arg(32 to 47) & X"000" & X"1") & \$313_res\ & eclat_true & \$v886\(32 to 47) & binop_int_arg(96 to 151) & binop_int_arg(152 to 153);
                      result2582 := binop_int_result;
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    else
                      modulo_arg := eclat_sub(modulo_arg(0 to 30) & modulo_arg(31 to 61)) & modulo_arg(31 to 61);
                      state_var3000 <= modulo;
                    end if;
                  when offsetclosure_n =>
                    offsetclosure_n_result := offsetclosure_n_arg(0 to 15) & eclat_resize(eclat_add(eclat_resize(offsetclosure_n_arg(48 to 78),16) & offsetclosure_n_arg(32 to 47)),31) & eclat_false & offsetclosure_n_arg(16 to 31) & offsetclosure_n_arg(80 to 135) & offsetclosure_n_arg(136 to 137);
                    result2582 := offsetclosure_n_result;
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getI2660 =>
                    state_var3000 <= pause_getII2661;
                  when pause_getI2672 =>
                    state_var3000 <= pause_getII2673;
                  when pause_getI2675 =>
                    state_var3000 <= pause_getII2676;
                  when pause_getI2678 =>
                    state_var3000 <= pause_getII2679;
                  when pause_getI2687 =>
                    state_var3000 <= pause_getII2688;
                  when pause_getI2690 =>
                    state_var3000 <= pause_getII2691;
                  when pause_getI2693 =>
                    state_var3000 <= pause_getII2694;
                  when pause_getI2697 =>
                    state_var3000 <= pause_getII2698;
                  when pause_getI2702 =>
                    state_var3000 <= pause_getII2703;
                  when pause_getI2705 =>
                    state_var3000 <= pause_getII2706;
                  when pause_getI2707 =>
                    state_var3000 <= pause_getII2708;
                  when pause_getI2709 =>
                    state_var3000 <= pause_getII2710;
                  when pause_getI2711 =>
                    state_var3000 <= pause_getII2712;
                  when pause_getI2713 =>
                    state_var3000 <= pause_getII2714;
                  when pause_getI2715 =>
                    state_var3000 <= pause_getII2716;
                  when pause_getI2717 =>
                    state_var3000 <= pause_getII2718;
                  when pause_getI2719 =>
                    state_var3000 <= pause_getII2720;
                  when pause_getI2723 =>
                    state_var3000 <= pause_getII2724;
                  when pause_getI2726 =>
                    state_var3000 <= pause_getII2727;
                  when pause_getI2729 =>
                    state_var3000 <= pause_getII2730;
                  when pause_getI2732 =>
                    state_var3000 <= pause_getII2733;
                  when pause_getI2735 =>
                    state_var3000 <= pause_getII2736;
                  when pause_getI2738 =>
                    state_var3000 <= pause_getII2739;
                  when pause_getI2741 =>
                    state_var3000 <= pause_getII2742;
                  when pause_getI2744 =>
                    state_var3000 <= pause_getII2745;
                  when pause_getI2746 =>
                    state_var3000 <= pause_getII2747;
                  when pause_getI2748 =>
                    state_var3000 <= pause_getII2749;
                  when pause_getI2750 =>
                    state_var3000 <= pause_getII2751;
                  when pause_getI2752 =>
                    state_var3000 <= pause_getII2753;
                  when pause_getI2755 =>
                    state_var3000 <= pause_getII2756;
                  when pause_getI2758 =>
                    state_var3000 <= pause_getII2759;
                  when pause_getI2761 =>
                    state_var3000 <= pause_getII2762;
                  when pause_getI2765 =>
                    state_var3000 <= pause_getII2766;
                  when pause_getI2768 =>
                    state_var3000 <= pause_getII2769;
                  when pause_getI2770 =>
                    state_var3000 <= pause_getII2771;
                  when pause_getI2776 =>
                    state_var3000 <= pause_getII2777;
                  when pause_getI2778 =>
                    state_var3000 <= pause_getII2779;
                  when pause_getI2780 =>
                    state_var3000 <= pause_getII2781;
                  when pause_getI2782 =>
                    state_var3000 <= pause_getII2783;
                  when pause_getI2785 =>
                    state_var3000 <= pause_getII2786;
                  when pause_getI2788 =>
                    state_var3000 <= pause_getII2789;
                  when pause_getI2791 =>
                    state_var3000 <= pause_getII2792;
                  when pause_getI2794 =>
                    state_var3000 <= pause_getII2795;
                  when pause_getI2796 =>
                    state_var3000 <= pause_getII2797;
                  when pause_getI2798 =>
                    state_var3000 <= pause_getII2799;
                  when pause_getI2800 =>
                    state_var3000 <= pause_getII2801;
                  when pause_getI2803 =>
                    state_var3000 <= pause_getII2804;
                  when pause_getI2805 =>
                    state_var3000 <= pause_getII2806;
                  when pause_getI2807 =>
                    state_var3000 <= pause_getII2808;
                  when pause_getI2809 =>
                    state_var3000 <= pause_getII2810;
                  when pause_getI2812 =>
                    state_var3000 <= pause_getII2813;
                  when pause_getI2814 =>
                    state_var3000 <= pause_getII2815;
                  when pause_getI2816 =>
                    state_var3000 <= pause_getII2817;
                  when pause_getI2818 =>
                    state_var3000 <= pause_getII2819;
                  when pause_getI2820 =>
                    state_var3000 <= pause_getII2821;
                  when pause_getI2822 =>
                    state_var3000 <= pause_getII2823;
                  when pause_getI2824 =>
                    state_var3000 <= pause_getII2825;
                  when pause_getI2830 =>
                    state_var3000 <= pause_getII2831;
                  when pause_getI2832 =>
                    state_var3000 <= pause_getII2833;
                  when pause_getI2836 =>
                    state_var3000 <= pause_getII2837;
                  when pause_getI2838 =>
                    state_var3000 <= pause_getII2839;
                  when pause_getI2844 =>
                    state_var3000 <= pause_getII2845;
                  when pause_getI2846 =>
                    state_var3000 <= pause_getII2847;
                  when pause_getI2848 =>
                    state_var3000 <= pause_getII2849;
                  when pause_getI2850 =>
                    state_var3000 <= pause_getII2851;
                  when pause_getI2852 =>
                    state_var3000 <= pause_getII2853;
                  when pause_getI2856 =>
                    state_var3000 <= pause_getII2857;
                  when pause_getI2859 =>
                    state_var3000 <= pause_getII2860;
                  when pause_getI2861 =>
                    state_var3000 <= pause_getII2862;
                  when pause_getI2863 =>
                    state_var3000 <= pause_getII2864;
                  when pause_getI2869 =>
                    state_var3000 <= pause_getII2870;
                  when pause_getI2871 =>
                    state_var3000 <= pause_getII2872;
                  when pause_getI2876 =>
                    state_var3000 <= pause_getII2877;
                  when pause_getI2879 =>
                    state_var3000 <= pause_getII2880;
                  when pause_getI2881 =>
                    state_var3000 <= pause_getII2882;
                  when pause_getI2883 =>
                    state_var3000 <= pause_getII2884;
                  when pause_getI2890 =>
                    state_var3000 <= pause_getII2891;
                  when pause_getI2894 =>
                    state_var3000 <= pause_getII2895;
                  when pause_getI2898 =>
                    state_var3000 <= pause_getII2899;
                  when pause_getI2900 =>
                    state_var3000 <= pause_getII2901;
                  when pause_getI2904 =>
                    state_var3000 <= pause_getII2905;
                  when pause_getI2906 =>
                    state_var3000 <= pause_getII2907;
                  when pause_getI2908 =>
                    state_var3000 <= pause_getII2909;
                  when pause_getI2912 =>
                    state_var3000 <= pause_getII2913;
                  when pause_getI2914 =>
                    state_var3000 <= pause_getII2915;
                  when pause_getI2916 =>
                    state_var3000 <= pause_getII2917;
                  when pause_getI2918 =>
                    state_var3000 <= pause_getII2919;
                  when pause_getI2922 =>
                    state_var3000 <= pause_getII2923;
                  when pause_getI2924 =>
                    state_var3000 <= pause_getII2925;
                  when pause_getI2926 =>
                    state_var3000 <= pause_getII2927;
                  when pause_getI2928 =>
                    state_var3000 <= pause_getII2929;
                  when pause_getI2932 =>
                    state_var3000 <= pause_getII2933;
                  when pause_getI2935 =>
                    state_var3000 <= pause_getII2936;
                  when pause_getI2938 =>
                    state_var3000 <= pause_getII2939;
                  when pause_getI2941 =>
                    state_var3000 <= pause_getII2942;
                  when pause_getI2947 =>
                    state_var3000 <= pause_getII2948;
                  when pause_getI2949 =>
                    state_var3000 <= pause_getII2950;
                  when pause_getI2951 =>
                    state_var3000 <= pause_getII2952;
                  when pause_getI2953 =>
                    state_var3000 <= pause_getII2954;
                  when pause_getI2957 =>
                    state_var3000 <= pause_getII2958;
                  when pause_getI2962 =>
                    state_var3000 <= pause_getII2963;
                  when pause_getI2966 =>
                    state_var3000 <= pause_getII2967;
                  when pause_getI2976 =>
                    state_var3000 <= pause_getII2977;
                  when pause_getI2979 =>
                    state_var3000 <= pause_getII2980;
                  when pause_getI2982 =>
                    state_var3000 <= pause_getII2983;
                  when pause_getI2985 =>
                    state_var3000 <= pause_getII2986;
                  when pause_getI2988 =>
                    state_var3000 <= pause_getII2989;
                  when pause_getII2661 =>
                    \$v274\ := \$ram_value\;
                    apply_result := eclat_resize(\$v274\(0 to 30),16) & apply_arg(60 to 91) & \$342_sp\ & apply_arg(60 to 91) & apply_arg(3 to 10) & apply_arg(148 to 163) & apply_arg(164 to 165);
                    result2582 := apply_result;
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2673 =>
                    \$1379_v\ := \$ram_value\;
                    \$v908\ := \$1379_v\ & eclat_sub(\$v907\(32 to 47) & X"000" & X"1");
                    \$v2671\ := ""&apply_arg(11);
                    if \$v2671\(0) = '1' then
                      \$339_sp\ := eclat_add(eclat_sub(\$v908\(32 to 47) & apply_arg(12 to 27)) & apply_arg(28 to 43));
                      \$v2667\ := ""&apply_arg(2);
                      if \$v2667\(0) = '1' then
                        \$ram_ptr_write\ <= to_integer(unsigned(\$339_sp\));
                        \$ram_write_request\ <= '1';
                        \$ram_write\ <= \$v908\(0 to 31);
                        state_var3000 <= pause_setI2666;
                      else
                        \$340_sp\ := \$339_sp\;
                        \$v2665\ := ""&apply_arg(1);
                        if \$v2665\(0) = '1' then
                          \$ram_ptr_write\ <= to_integer(unsigned(\$340_sp\));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$v907\(0 to 31);
                          state_var3000 <= pause_setI2664;
                        else
                          \$341_sp\ := \$340_sp\;
                          \$v2663\ := ""&apply_arg(0);
                          if \$v2663\(0) = '1' then
                            \$ram_ptr_write\ <= to_integer(unsigned(\$341_sp\));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$v906\(0 to 31);
                            state_var3000 <= pause_setI2662;
                          else
                            \$342_sp\ := \$341_sp\;
                            \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(apply_arg(60 to 90),16) & X"000" & X"0") & X"000" & X"1")));
                            state_var3000 <= pause_getI2660;
                          end if;
                        end if;
                      end if;
                    else
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v908\(32 to 47)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= eclat_resize(apply_arg(140 to 147),31) & eclat_true;
                      state_var3000 <= pause_setI2670;
                    end if;
                  when pause_getII2676 =>
                    \$1381_v\ := \$ram_value\;
                    \$v907\ := \$1381_v\ & eclat_sub(\$v906\(32 to 47) & X"000" & X"1");
                    \$v2674\ := ""&apply_arg(2);
                    if \$v2674\(0) = '1' then
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v907\(32 to 47) & X"000" & X"1")));
                      state_var3000 <= pause_getI2672;
                    else
                      \$v908\ := "000"& X"000000" & X"1" & eclat_true & \$v907\(32 to 47);
                      \$v2671\ := ""&apply_arg(11);
                      if \$v2671\(0) = '1' then
                        \$339_sp\ := eclat_add(eclat_sub(\$v908\(32 to 47) & apply_arg(12 to 27)) & apply_arg(28 to 43));
                        \$v2667\ := ""&apply_arg(2);
                        if \$v2667\(0) = '1' then
                          \$ram_ptr_write\ <= to_integer(unsigned(\$339_sp\));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$v908\(0 to 31);
                          state_var3000 <= pause_setI2666;
                        else
                          \$340_sp\ := \$339_sp\;
                          \$v2665\ := ""&apply_arg(1);
                          if \$v2665\(0) = '1' then
                            \$ram_ptr_write\ <= to_integer(unsigned(\$340_sp\));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$v907\(0 to 31);
                            state_var3000 <= pause_setI2664;
                          else
                            \$341_sp\ := \$340_sp\;
                            \$v2663\ := ""&apply_arg(0);
                            if \$v2663\(0) = '1' then
                              \$ram_ptr_write\ <= to_integer(unsigned(\$341_sp\));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$v906\(0 to 31);
                              state_var3000 <= pause_setI2662;
                            else
                              \$342_sp\ := \$341_sp\;
                              \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(apply_arg(60 to 90),16) & X"000" & X"0") & X"000" & X"1")));
                              state_var3000 <= pause_getI2660;
                            end if;
                          end if;
                        end if;
                      else
                        \$ram_ptr_write\ <= to_integer(unsigned(\$v908\(32 to 47)));
                        \$ram_write_request\ <= '1';
                        \$ram_write\ <= eclat_resize(apply_arg(140 to 147),31) & eclat_true;
                        state_var3000 <= pause_setI2670;
                      end if;
                    end if;
                  when pause_getII2679 =>
                    \$1383_v\ := \$ram_value\;
                    \$v906\ := \$1383_v\ & eclat_sub(apply_arg(92 to 107) & X"000" & X"1");
                    \$v2677\ := ""&apply_arg(1);
                    if \$v2677\(0) = '1' then
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v906\(32 to 47) & X"000" & X"1")));
                      state_var3000 <= pause_getI2675;
                    else
                      \$v907\ := "000"& X"000000" & X"1" & eclat_true & \$v906\(32 to 47);
                      \$v2674\ := ""&apply_arg(2);
                      if \$v2674\(0) = '1' then
                        \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v907\(32 to 47) & X"000" & X"1")));
                        state_var3000 <= pause_getI2672;
                      else
                        \$v908\ := "000"& X"000000" & X"1" & eclat_true & \$v907\(32 to 47);
                        \$v2671\ := ""&apply_arg(11);
                        if \$v2671\(0) = '1' then
                          \$339_sp\ := eclat_add(eclat_sub(\$v908\(32 to 47) & apply_arg(12 to 27)) & apply_arg(28 to 43));
                          \$v2667\ := ""&apply_arg(2);
                          if \$v2667\(0) = '1' then
                            \$ram_ptr_write\ <= to_integer(unsigned(\$339_sp\));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$v908\(0 to 31);
                            state_var3000 <= pause_setI2666;
                          else
                            \$340_sp\ := \$339_sp\;
                            \$v2665\ := ""&apply_arg(1);
                            if \$v2665\(0) = '1' then
                              \$ram_ptr_write\ <= to_integer(unsigned(\$340_sp\));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$v907\(0 to 31);
                              state_var3000 <= pause_setI2664;
                            else
                              \$341_sp\ := \$340_sp\;
                              \$v2663\ := ""&apply_arg(0);
                              if \$v2663\(0) = '1' then
                                \$ram_ptr_write\ <= to_integer(unsigned(\$341_sp\));
                                \$ram_write_request\ <= '1';
                                \$ram_write\ <= \$v906\(0 to 31);
                                state_var3000 <= pause_setI2662;
                              else
                                \$342_sp\ := \$341_sp\;
                                \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(apply_arg(60 to 90),16) & X"000" & X"0") & X"000" & X"1")));
                                state_var3000 <= pause_getI2660;
                              end if;
                            end if;
                          end if;
                        else
                          \$ram_ptr_write\ <= to_integer(unsigned(\$v908\(32 to 47)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= eclat_resize(apply_arg(140 to 147),31) & eclat_true;
                          state_var3000 <= pause_setI2670;
                        end if;
                      end if;
                    end if;
                  when pause_getII2688 =>
                    \$1353_v\ := \$ram_value\;
                    \$v886\ := \$1353_v\ & eclat_sub(binop_int_arg(80 to 95) & X"000" & X"1");
                    \$v2686\ := binop_int_arg(0 to 31);
                    case \$v2686\ is
                    when X"0000000" & X"0" =>
                      \$313_res\ := eclat_add(binop_int_arg(48 to 78) & \$v886\(0 to 30));
                      binop_int_result := eclat_add(binop_int_arg(32 to 47) & X"000" & X"1") & \$313_res\ & eclat_true & \$v886\(32 to 47) & binop_int_arg(96 to 151) & binop_int_arg(152 to 153);
                      result2582 := binop_int_result;
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    when X"0000000" & X"1" =>
                      \$313_res\ := eclat_sub(binop_int_arg(48 to 78) & \$v886\(0 to 30));
                      binop_int_result := eclat_add(binop_int_arg(32 to 47) & X"000" & X"1") & \$313_res\ & eclat_true & \$v886\(32 to 47) & binop_int_arg(96 to 151) & binop_int_arg(152 to 153);
                      result2582 := binop_int_result;
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    when X"0000000" & X"2" =>
                      \$313_res\ := eclat_mult(binop_int_arg(48 to 78) & \$v886\(0 to 30));
                      binop_int_result := eclat_add(binop_int_arg(32 to 47) & X"000" & X"1") & \$313_res\ & eclat_true & \$v886\(32 to 47) & binop_int_arg(96 to 151) & binop_int_arg(152 to 153);
                      result2582 := binop_int_result;
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    when X"0000000" & X"3" =>
                      \$v2683\ := eclat_eq(\$v886\(0 to 30) & "000"& X"000000" & X"0");
                      if \$v2683\(0) = '1' then
                        \$313_res\ := "000"& X"000000" & X"0";
                        binop_int_result := eclat_add(binop_int_arg(32 to 47) & X"000" & X"1") & \$313_res\ & eclat_true & \$v886\(32 to 47) & binop_int_arg(96 to 151) & binop_int_arg(152 to 153);
                        result2582 := binop_int_result;
                        rdy2583 := eclat_true;
                        state_var3000 <= compute2584;
                      else
                        modulo_arg := eclat_abs(binop_int_arg(48 to 78)) & eclat_abs(\$v886\(0 to 30));
                        state_var3000 <= modulo;
                      end if;
                    when X"0000000" & X"4" =>
                      \$v2685\ := eclat_eq(\$v886\(0 to 30) & "000"& X"000000" & X"0");
                      if \$v2685\(0) = '1' then
                        \$313_res\ := "000"& X"000000" & X"0";
                        binop_int_result := eclat_add(binop_int_arg(32 to 47) & X"000" & X"1") & \$313_res\ & eclat_true & \$v886\(32 to 47) & binop_int_arg(96 to 151) & binop_int_arg(152 to 153);
                        result2582 := binop_int_result;
                        rdy2583 := eclat_true;
                        state_var3000 <= compute2584;
                      else
                        \$1342_modulo_arg\ := eclat_abs(binop_int_arg(48 to 78)) & eclat_abs(\$v886\(0 to 30));
                        state_var3000 <= \$1342_modulo\;
                      end if;
                    when X"0000000" & X"5" =>
                      \$313_res\ := eclat_land(binop_int_arg(48 to 78) & \$v886\(0 to 30));
                      binop_int_result := eclat_add(binop_int_arg(32 to 47) & X"000" & X"1") & \$313_res\ & eclat_true & \$v886\(32 to 47) & binop_int_arg(96 to 151) & binop_int_arg(152 to 153);
                      result2582 := binop_int_result;
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    when X"0000000" & X"6" =>
                      \$313_res\ := eclat_lor(binop_int_arg(48 to 78) & \$v886\(0 to 30));
                      binop_int_result := eclat_add(binop_int_arg(32 to 47) & X"000" & X"1") & \$313_res\ & eclat_true & \$v886\(32 to 47) & binop_int_arg(96 to 151) & binop_int_arg(152 to 153);
                      result2582 := binop_int_result;
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    when X"0000000" & X"7" =>
                      \$313_res\ := eclat_lxor(binop_int_arg(48 to 78) & \$v886\(0 to 30));
                      binop_int_result := eclat_add(binop_int_arg(32 to 47) & X"000" & X"1") & \$313_res\ & eclat_true & \$v886\(32 to 47) & binop_int_arg(96 to 151) & binop_int_arg(152 to 153);
                      result2582 := binop_int_result;
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    when X"0000000" & X"8" =>
                      \$313_res\ := eclat_lsl(binop_int_arg(48 to 78) & \$v886\(0 to 30));
                      binop_int_result := eclat_add(binop_int_arg(32 to 47) & X"000" & X"1") & \$313_res\ & eclat_true & \$v886\(32 to 47) & binop_int_arg(96 to 151) & binop_int_arg(152 to 153);
                      result2582 := binop_int_result;
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    when X"0000000" & X"9" =>
                      \$313_res\ := eclat_lsr(binop_int_arg(48 to 78) & \$v886\(0 to 30));
                      binop_int_result := eclat_add(binop_int_arg(32 to 47) & X"000" & X"1") & \$313_res\ & eclat_true & \$v886\(32 to 47) & binop_int_arg(96 to 151) & binop_int_arg(152 to 153);
                      result2582 := binop_int_result;
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    when X"0000000" & X"a" =>
                      \$313_res\ := eclat_asr(binop_int_arg(48 to 78) & \$v886\(0 to 30));
                      binop_int_result := eclat_add(binop_int_arg(32 to 47) & X"000" & X"1") & \$313_res\ & eclat_true & \$v886\(32 to 47) & binop_int_arg(96 to 151) & binop_int_arg(152 to 153);
                      result2582 := binop_int_result;
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    when X"0000000" & X"b" =>
                      \$313_res\ := eclat_if(eclat_lt(binop_int_arg(48 to 78) & "000"& X"000000" & X"0") & 
                                    eclat_if(eclat_lt(\$v886\(0 to 30) & "000"& X"000000" & X"0") & 
                                    eclat_if(eclat_gt(binop_int_arg(48 to 78) & \$v886\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"0") & 
                                    eclat_if(eclat_lt(\$v886\(0 to 30) & "000"& X"000000" & X"0") & "000"& X"000000" & X"0" & 
                                    eclat_if(eclat_lt(binop_int_arg(48 to 78) & \$v886\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                      binop_int_result := eclat_add(binop_int_arg(32 to 47) & X"000" & X"1") & \$313_res\ & eclat_true & \$v886\(32 to 47) & binop_int_arg(96 to 151) & binop_int_arg(152 to 153);
                      result2582 := binop_int_result;
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    when X"0000000" & X"c" =>
                      \$313_res\ := eclat_if(eclat_lt(binop_int_arg(48 to 78) & "000"& X"000000" & X"0") & 
                                    eclat_if(eclat_lt(\$v886\(0 to 30) & "000"& X"000000" & X"0") & 
                                    eclat_if(eclat_le(binop_int_arg(48 to 78) & \$v886\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"1") & 
                                    eclat_if(eclat_lt(\$v886\(0 to 30) & "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & 
                                    eclat_if(eclat_ge(binop_int_arg(48 to 78) & \$v886\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                      binop_int_result := eclat_add(binop_int_arg(32 to 47) & X"000" & X"1") & \$313_res\ & eclat_true & \$v886\(32 to 47) & binop_int_arg(96 to 151) & binop_int_arg(152 to 153);
                      result2582 := binop_int_result;
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    when others =>
                      \$313_res\ := "000"& X"000000" & X"0";
                      binop_int_result := eclat_add(binop_int_arg(32 to 47) & X"000" & X"1") & \$313_res\ & eclat_true & \$v886\(32 to 47) & binop_int_arg(96 to 151) & binop_int_arg(152 to 153);
                      result2582 := binop_int_result;
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    end case;
                  when pause_getII2691 =>
                    \$1330_v\ := \$ram_value\;
                    \$v878\ := \$1330_v\ & eclat_sub(binop_compare_arg(80 to 95) & X"000" & X"1");
                    compare_id := X"00" & X"d";
                    compare_arg := binop_compare_arg(0 to 31) & binop_compare_arg(48 to 78) & \$v878\(0 to 30);
                    state_var3000 <= compare;
                  when pause_getII2694 =>
                    \$1308_v\ := \$ram_value\;
                    \$v868\ := \$1308_v\ & eclat_sub(\$288_sp\ & X"000" & X"1");
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v866\(64 to 94),16) & X"000" & X"2") & X"000" & X"1")));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v868\(0 to 31);
                    state_var3000 <= pause_setI2692;
                  when pause_getII2698 =>
                    \$1315_v\ := \$ram_value\;
                    \$v871\ := \$1315_v\ & eclat_sub(make_block_n_arg(16 to 31) & X"000" & X"1");
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v866\(64 to 94),16) & X"000" & X"1") & X"000" & X"1")));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v871\(0 to 31);
                    state_var3000 <= pause_setI2696;
                  when pause_getII2703 =>
                    arg := \$code_value\;
                    branch_if_result := eclat_add(eclat_add(branch_if_arg(1 to 16) & X"000" & X"1") & eclat_resize(arg,16)) & branch_if_arg(17 to 48) & branch_if_arg(49 to 64) & branch_if_arg(65 to 120) & branch_if_arg(121 to 122);
                    result2582 := branch_if_result;
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2706 =>
                    \$951_v\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$951_v\ & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2708 =>
                    \$955_v\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$955_v\ & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2710 =>
                    \$959_v\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$959_v\ & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2712 =>
                    \$963_v\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$963_v\ & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2714 =>
                    \$967_v\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$967_v\ & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2716 =>
                    \$971_v\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$971_v\ & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2718 =>
                    \$975_v\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$975_v\ & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2720 =>
                    \$979_v\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$979_v\ & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2724 =>
                    \$984_v\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$984_v\ & \$983_sp\ & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2727 =>
                    \$989_v\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$989_v\ & \$988_sp\ & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2730 =>
                    \$994_v\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$994_v\ & \$993_sp\ & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2733 =>
                    \$999_v\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$999_v\ & \$998_sp\ & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2736 =>
                    \$1004_v\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$1004_v\ & \$1003_sp\ & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2739 =>
                    \$1009_v\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$1009_v\ & \$1008_sp\ & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2742 =>
                    \$1014_v\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$1014_v\ & \$1013_sp\ & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2745 =>
                    \$1017\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$1017\ & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2747 =>
                    \$1025\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$1025\ & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2749 =>
                    \$1033\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$1033\ & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2751 =>
                    \$1041\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$1041\ & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2753 =>
                    \$1049\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$1049\ & \$1048_sp\ & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2756 =>
                    \$1058\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$1058\ & \$1057_sp\ & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2759 =>
                    \$1067\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$1067\ & \$1066_sp\ & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2762 =>
                    \$1076\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$1076\ & \$1075_sp\ & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2766 =>
                    \$v225\ := \$ram_value\;
                    \$ram_ptr_write\ <= to_integer(unsigned(loop_push_arg(0 to 15)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v225\;
                    state_var3000 <= pause_setI2764;
                  when pause_getII2769 =>
                    \$236_next_env\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$v522\(16 to 47) & \$235_sp\ & \$236_next_env\ & eclat_add(\$v522\(96 to 103) & eclat_sub(eclat_resize(\$v227\,8) & X"0" & X"2")) & \$v522\(104 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2771 =>
                    \$592_hd\ := \$ram_value\;
                    \$v227\ := eclat_resize(eclat_lsr(eclat_resize(eclat_resize(\$592_hd\(0 to 30),16),31) & "000"& X"000000" & X"2"),16);
                    loop_push_arg := \$v522\(48 to 63) & X"0" & X"0" & \$v522\(64 to 95) & eclat_resize(\$v227\,8);
                    state_var3000 <= loop_push;
                  when pause_getII2777 =>
                    \$1109_v\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$1109_v\ & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2779 =>
                    \$1119_v\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$1119_v\ & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2781 =>
                    \$1129_v\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$1129_v\ & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2783 =>
                    \$1139_v\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$1139_v\ & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2786 =>
                    \$1153_v\ := \$ram_value\;
                    \$v796\ := \$1153_v\ & eclat_sub(\$v522\(48 to 63) & X"000" & X"1");
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v522\(16 to 46),16) & X"000" & X"0") & X"000" & X"1")));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v796\(0 to 31);
                    state_var3000 <= pause_setI2784;
                  when pause_getII2789 =>
                    \$1163_v\ := \$ram_value\;
                    \$v799\ := \$1163_v\ & eclat_sub(\$v522\(48 to 63) & X"000" & X"1");
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v522\(16 to 46),16) & X"000" & X"1") & X"000" & X"1")));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v799\(0 to 31);
                    state_var3000 <= pause_setI2787;
                  when pause_getII2792 =>
                    \$1173_v\ := \$ram_value\;
                    \$v802\ := \$1173_v\ & eclat_sub(\$v522\(48 to 63) & X"000" & X"1");
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v522\(16 to 46),16) & X"000" & X"2") & X"000" & X"1")));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v802\(0 to 31);
                    state_var3000 <= pause_setI2790;
                  when pause_getII2795 =>
                    \$1183_v\ := \$ram_value\;
                    \$v805\ := \$1183_v\ & eclat_sub(\$v522\(48 to 63) & X"000" & X"1");
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v522\(16 to 46),16) & X"000" & X"3") & X"000" & X"1")));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v805\(0 to 31);
                    state_var3000 <= pause_setI2793;
                  when pause_getII2797 =>
                    \$1186_hd\ := \$ram_value\;
                    \$v234\ := eclat_resize(eclat_lsr(eclat_resize(eclat_resize(\$1186_hd\(0 to 30),16),31) & "000"& X"000000" & X"2"),16);
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & eclat_resize(\$v234\,31) & eclat_true & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2799 =>
                    \$245_v\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$245_v\ & \$v810\(32 to 47) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2801 =>
                    \$1200_v\ := \$ram_value\;
                    \$v810\ := \$1200_v\ & eclat_sub(\$v522\(48 to 63) & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v522\(16 to 46),16) & eclat_resize(\$v810\(0 to 30),16)) & X"000" & X"1")));
                    state_var3000 <= pause_getI2798;
                  when pause_getII2804 =>
                    \$1208_v\ := \$ram_value\;
                    \$v814\ := \$1208_v\ & eclat_sub(\$v813\(32 to 47) & X"000" & X"1");
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v522\(16 to 46),16) & eclat_resize(\$v813\(0 to 30),16)) & X"000" & X"1")));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v814\(0 to 31);
                    state_var3000 <= pause_setI2802;
                  when pause_getII2806 =>
                    \$1210_v\ := \$ram_value\;
                    \$v813\ := \$1210_v\ & eclat_sub(\$v522\(48 to 63) & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v813\(32 to 47) & X"000" & X"1")));
                    state_var3000 <= pause_getI2803;
                  when pause_getII2808 =>
                    \$253_next_acc\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$253_next_acc\ & \$v818\(32 to 47) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2810 =>
                    \$1218_v\ := \$ram_value\;
                    \$v818\ := \$1218_v\ & eclat_sub(\$v522\(48 to 63) & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v522\(16 to 46),16) & eclat_resize(\$v818\(0 to 30),16)) & X"000" & X"1")));
                    state_var3000 <= pause_getI2807;
                  when pause_getII2813 =>
                    \$1226_v\ := \$ram_value\;
                    \$v822\ := \$1226_v\ & eclat_sub(\$v821\(32 to 47) & X"000" & X"1");
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v522\(16 to 46),16) & eclat_resize(\$v821\(0 to 30),16)) & X"000" & X"1")));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v822\(0 to 31);
                    state_var3000 <= pause_setI2811;
                  when pause_getII2815 =>
                    \$1228_v\ := \$ram_value\;
                    \$v821\ := \$1228_v\ & eclat_sub(\$v522\(48 to 63) & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v821\(32 to 47) & X"000" & X"1")));
                    state_var3000 <= pause_getI2812;
                  when pause_getII2817 =>
                    \$1235_v\ := \$ram_value\;
                    \$v827\ := \$1235_v\ & eclat_sub(eclat_sub(\$v522\(48 to 63) & X"000" & X"1") & X"000" & X"1");
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$v522\(16 to 47) & eclat_sub(\$v827\(32 to 47) & X"000" & X"2") & \$v522\(64 to 95) & \$v522\(96 to 103) & eclat_resize(\$v827\(0 to 30),16) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2819 =>
                    \$1239_v\ := \$ram_value\;
                    \$v832\ := \$1239_v\ & eclat_sub(\$v831\(32 to 47) & X"000" & X"1");
                    result2582 := eclat_resize(\$v829\(0 to 30),16) & \$v522\(16 to 47) & \$v832\(32 to 47) & \$v831\(0 to 31) & eclat_resize(\$v832\(0 to 30),8) & eclat_resize(\$v830\(0 to 30),16) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2821 =>
                    \$1241_v\ := \$ram_value\;
                    \$v831\ := \$1241_v\ & eclat_sub(\$v830\(32 to 47) & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v831\(32 to 47) & X"000" & X"1")));
                    state_var3000 <= pause_getI2818;
                  when pause_getII2823 =>
                    \$1245_v\ := \$ram_value\;
                    \$v830\ := \$1245_v\ & eclat_sub(\$v829\(32 to 47) & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v830\(32 to 47) & X"000" & X"1")));
                    state_var3000 <= pause_getI2820;
                  when pause_getII2825 =>
                    \$1249_v\ := \$ram_value\;
                    \$v829\ := \$1249_v\ & eclat_sub(\$v522\(104 to 119) & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v829\(32 to 47) & X"000" & X"1")));
                    state_var3000 <= pause_getI2822;
                  when pause_getII2831 =>
                    \$368_v\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$368_v\ & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2833 =>
                    \$770_v\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"2") & \$770_v\ & \$357_sp\ & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2837 =>
                    \$v287\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"2") & \$v287\ & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2839 =>
                    \$778\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"2") & \$778\ & \$354_sp\ & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2845 =>
                    \$v134\ := \$ram_value\;
                    result2582 := eclat_resize(\$v134\(0 to 30),16) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(16 to 47) & eclat_sub(eclat_resize(argument1,8) & X"0" & X"1") & \$v522\(104 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2847 =>
                    \$v146\ := \$ram_value\;
                    result2582 := eclat_resize(\$v146\(0 to 30),16) & \$v522\(16 to 47) & eclat_sub(\$v522\(48 to 63) & eclat_resize(argument1,16)) & \$v522\(16 to 47) & eclat_sub(\$v522\(96 to 103) & X"0" & X"1") & \$v522\(104 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2849 =>
                    \$794_v\ := \$ram_value\;
                    \$v615\ := \$794_v\ & eclat_sub(\$v614\(32 to 47) & X"000" & X"1");
                    result2582 := eclat_resize(\$v613\(0 to 30),16) & \$v522\(16 to 47) & \$v615\(32 to 47) & \$v614\(0 to 31) & eclat_resize(\$v615\(0 to 30),8) & \$v522\(104 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2851 =>
                    \$796_v\ := \$ram_value\;
                    \$v614\ := \$796_v\ & eclat_sub(\$v613\(32 to 47) & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v614\(32 to 47) & X"000" & X"1")));
                    state_var3000 <= pause_getI2848;
                  when pause_getII2853 =>
                    \$800_v\ := \$ram_value\;
                    \$v613\ := \$800_v\ & eclat_sub(eclat_sub(\$v522\(48 to 63) & eclat_resize(argument1,16)) & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v613\(32 to 47) & X"000" & X"1")));
                    state_var3000 <= pause_getI2850;
                  when pause_getII2857 =>
                    \$826_v\ := \$ram_value\;
                    \$v632\ := \$826_v\ & eclat_sub(\$103_w_arg\(8 to 23) & X"000" & X"1");
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$103_w_arg\(24 to 54),16) & eclat_resize(eclat_add(\$103_w_arg\(0 to 7) & X"0" & X"2"),16)) & X"000" & X"1")));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v632\(0 to 31);
                    state_var3000 <= pause_setI2855;
                  when pause_getII2860 =>
                    \$811_v\ := \$ram_value\;
                    \$v625\ := \$811_v\ & eclat_sub(\$v624\(32 to 47) & X"000" & X"1");
                    result2582 := eclat_resize(\$v623\(0 to 30),16) & \$v620\(64 to 95) & \$v625\(32 to 47) & \$v624\(0 to 31) & eclat_resize(\$v625\(0 to 30),8) & \$v522\(104 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2862 =>
                    \$813_v\ := \$ram_value\;
                    \$v624\ := \$813_v\ & eclat_sub(\$v623\(32 to 47) & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v624\(32 to 47) & X"000" & X"1")));
                    state_var3000 <= pause_getI2859;
                  when pause_getII2864 =>
                    \$817_v\ := \$ram_value\;
                    \$v623\ := \$817_v\ & eclat_sub(\$104_sp\ & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v623\(32 to 47) & X"000" & X"1")));
                    state_var3000 <= pause_getI2861;
                  when pause_getII2870 =>
                    \$120_v\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"2") & \$120_v\ & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2872 =>
                    \$122_v\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"2") & \$122_v\ & eclat_add(\$v522\(48 to 63) & X"000" & X"1") & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2877 =>
                    \$321_v\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"2") & \$321_v\ & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2880 =>
                    \$852_v\ := \$ram_value\;
                    \$v649\ := \$852_v\ & eclat_sub(\$v522\(48 to 63) & X"000" & X"1");
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v522\(16 to 46),16) & eclat_resize(argument1,16)) & X"000" & X"1")));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v649\(0 to 31);
                    state_var3000 <= pause_setI2878;
                  when pause_getII2882 =>
                    \$v179\ := \$code_value\;
                    result2582 := eclat_add(eclat_add(\$v522\(0 to 15) & X"000" & X"2") & eclat_resize(\$v179\,16)) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2884 =>
                    \$590_hd\ := \$ram_value\;
                    idx := eclat_lsr(eclat_resize(\$590_hd\(0 to 30),16) & X"00" & X"18");
                    \$125_ofs\ := eclat_add(eclat_resize(argument1,16) & idx);
                    \$code_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(\$v522\(0 to 15) & X"000" & X"2") & \$125_ofs\)));
                    state_var3000 <= pause_getI2881;
                  when pause_getII2891 =>
                    \$864_v\ := \$ram_value\;
                    \$v668\ := \$864_v\ & eclat_sub(\$v665\(80 to 95) & X"000" & X"1");
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"2") & \$v665\(0 to 31) & \$v668\(32 to 47) & \$v668\(0 to 31) & \$v665\(128 to 135) & \$v665\(136 to 151) & \$v665\(152 to 153);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2895 =>
                    \$868_v\ := \$ram_value\;
                    \$v680\ := \$868_v\ & eclat_sub(\$v677\(80 to 95) & X"000" & X"1");
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"2") & \$v677\(0 to 31) & \$v680\(32 to 47) & \$v680\(0 to 31) & \$v677\(128 to 135) & \$v677\(136 to 151) & \$v677\(152 to 153);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2899 =>
                    \$876_v\ := \$ram_value\;
                    \$v676\ := \$876_v\ & eclat_sub(\$v522\(48 to 63) & X"000" & X"1");
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v676\(32 to 47)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v522\(64 to 95);
                    state_var3000 <= pause_setI2897;
                  when pause_getII2901 =>
                    \$878_v\ := \$ram_value\;
                    \$v693\ := \$878_v\ & eclat_sub(\$v690\(80 to 95) & X"000" & X"1");
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"2") & \$v690\(0 to 31) & \$v693\(32 to 47) & \$v693\(0 to 31) & \$v690\(128 to 135) & \$v690\(136 to 151) & \$v690\(152 to 153);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2905 =>
                    \$886_v\ := \$ram_value\;
                    \$v689\ := \$886_v\ & eclat_sub(\$v688\(32 to 47) & X"000" & X"1");
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v689\(32 to 47)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v522\(64 to 95);
                    state_var3000 <= pause_setI2903;
                  when pause_getII2907 =>
                    \$888_v\ := \$ram_value\;
                    \$v688\ := \$888_v\ & eclat_sub(\$v522\(48 to 63) & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v688\(32 to 47) & X"000" & X"1")));
                    state_var3000 <= pause_getI2904;
                  when pause_getII2909 =>
                    \$890_v\ := \$ram_value\;
                    \$v707\ := \$890_v\ & eclat_sub(\$v704\(80 to 95) & X"000" & X"1");
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"2") & \$v704\(0 to 31) & \$v707\(32 to 47) & \$v707\(0 to 31) & \$v704\(128 to 135) & \$v704\(136 to 151) & \$v704\(152 to 153);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2913 =>
                    \$898_v\ := \$ram_value\;
                    \$v703\ := \$898_v\ & eclat_sub(\$v702\(32 to 47) & X"000" & X"1");
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v703\(32 to 47)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v522\(64 to 95);
                    state_var3000 <= pause_setI2911;
                  when pause_getII2915 =>
                    \$900_v\ := \$ram_value\;
                    \$v702\ := \$900_v\ & eclat_sub(\$v701\(32 to 47) & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v702\(32 to 47) & X"000" & X"1")));
                    state_var3000 <= pause_getI2912;
                  when pause_getII2917 =>
                    \$902_v\ := \$ram_value\;
                    \$v701\ := \$902_v\ & eclat_sub(\$v522\(48 to 63) & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v701\(32 to 47) & X"000" & X"1")));
                    state_var3000 <= pause_getI2914;
                  when pause_getII2919 =>
                    \$904_v\ := \$ram_value\;
                    \$v722\ := \$904_v\ & eclat_sub(\$v719\(80 to 95) & X"000" & X"1");
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"2") & \$v719\(0 to 31) & \$v722\(32 to 47) & \$v722\(0 to 31) & \$v719\(128 to 135) & \$v719\(136 to 151) & \$v719\(152 to 153);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2923 =>
                    \$912_v\ := \$ram_value\;
                    \$v718\ := \$912_v\ & eclat_sub(\$v717\(32 to 47) & X"000" & X"1");
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v718\(32 to 47)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v522\(64 to 95);
                    state_var3000 <= pause_setI2921;
                  when pause_getII2925 =>
                    \$914_v\ := \$ram_value\;
                    \$v717\ := \$914_v\ & eclat_sub(\$v716\(32 to 47) & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v717\(32 to 47) & X"000" & X"1")));
                    state_var3000 <= pause_getI2922;
                  when pause_getII2927 =>
                    \$916_v\ := \$ram_value\;
                    \$v716\ := \$916_v\ & eclat_sub(\$v715\(32 to 47) & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v716\(32 to 47) & X"000" & X"1")));
                    state_var3000 <= pause_getI2924;
                  when pause_getII2929 =>
                    \$918_v\ := \$ram_value\;
                    \$v715\ := \$918_v\ & eclat_sub(\$v522\(48 to 63) & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v715\(32 to 47) & X"000" & X"1")));
                    state_var3000 <= pause_getI2926;
                  when pause_getII2933 =>
                    f0 := \$ram_value\;
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v522\(16 to 46),16) & X"000" & X"0") & X"000" & X"1")));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= eclat_add(f0(0 to 30) & argument1) & eclat_true;
                    state_var3000 <= pause_setI2931;
                  when pause_getII2936 =>
                    \$v86\ := \$ram_value\;
                    \$v87\ := eclat_sub(eclat_sub(eclat_sub(w_arg(16 to 31) & w_arg(32 to 47)) & w_arg(48 to 63)) & w_arg(0 to 15)) & \$v86\;
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v87\(0 to 15)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v87\(16 to 47);
                    state_var3000 <= pause_setI2934;
                  when pause_getII2939 =>
                    \$v80\ := \$ram_value\;
                    result2582 := eclat_resize(\$v80\(0 to 30),16) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(16 to 47) & eclat_sub(eclat_add(\$v522\(96 to 103) & eclat_resize(argument1,8)) & X"0" & X"1") & \$v522\(104 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2942 =>
                    \$735_v\ := \$ram_value\;
                    \$v581\ := \$735_v\ & eclat_sub(fill_arg(16 to 31) & X"000" & X"1");
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(fill_arg(48 to 78),16) & fill_arg(0 to 15)) & X"000" & X"1")));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v581\(0 to 31);
                    state_var3000 <= pause_setI2940;
                  when pause_getII2948 =>
                    \$66_v\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"3") & \$66_v\ & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2950 =>
                    \$v100\ := \$ram_value\;
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v100\(0 to 30),16) & eclat_resize(argument2,16)) & X"000" & X"1")));
                    state_var3000 <= pause_getI2947;
                  when pause_getII2952 =>
                    \$70_v\ := \$ram_value\;
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"3") & \$70_v\ & eclat_add(\$v522\(48 to 63) & X"000" & X"1") & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2954 =>
                    \$v104\ := \$ram_value\;
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v104\(0 to 30),16) & eclat_resize(argument2,16)) & X"000" & X"1")));
                    state_var3000 <= pause_getI2951;
                  when pause_getII2958 =>
                    \$762_v\ := \$ram_value\;
                    \$v599\ := \$762_v\ & eclat_sub(\$74_fill_arg\(16 to 31) & X"000" & X"1");
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$74_fill_arg\(32 to 62),16) & \$74_fill_arg\(0 to 15)) & X"000" & X"1")));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v599\(0 to 31);
                    state_var3000 <= pause_setI2956;
                  when pause_getII2963 =>
                    \$660_v\ := \$ram_value\;
                    \$v563\ := \$660_v\ & eclat_sub(w0_arg(16 to 31) & X"000" & X"1");
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(w0_arg(48 to 78),16) & eclat_sub(eclat_add(w0_arg(0 to 15) & eclat_mult(X"000" & X"2" & w0_arg(32 to 47))) & X"000" & X"1")) & X"000" & X"1")));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v563\(0 to 31);
                    state_var3000 <= pause_setI2961;
                  when pause_getII2967 =>
                    \$v44\ := \$code_value\;
                    \$v51\ := w1_arg(48 to 79) & eclat_mult(X"000" & X"2" & w1_arg(0 to 15)) & eclat_resize(eclat_add(eclat_add(w1_arg(16 to 31) & X"000" & X"2") & eclat_resize(\$v44\,16)),31) & eclat_true;
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v51\(0 to 30),16) & \$v51\(32 to 47)) & X"000" & X"1")));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v51\(48 to 79);
                    state_var3000 <= pause_setI2965;
                  when pause_getII2977 =>
                    \$v29\ := \$code_value\;
                    eclat_print_int(\$v29\);
                    
                    eclat_print_newline(eclat_unit);
                    
                    result2582 := \$v522\(0 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_getII2980 =>
                    argument3 := \$code_value\;
                    \$v2978\ := eclat_resize(\$v259\,8);
                    case \$v2978\ is
                    when X"2c" =>
                      \$v2975\ := eclat_gt(eclat_resize(argument2,16) & X"000" & X"0");
                      if \$v2975\(0) = '1' then
                        \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                        \$ram_write_request\ <= '1';
                        \$ram_write\ <= \$v522\(16 to 47);
                        state_var3000 <= pause_setI2974;
                      else
                        \$30_sp\ := \$v522\(48 to 63);
                        make_block_id := X"0" & X"53";
                        make_block_arg := \$30_sp\ & \$v522\(16 to 47) & \$v522\(64 to 95) & X"f7" & eclat_add(eclat_sub(eclat_mult(X"000" & X"2" & eclat_resize(argument1,16)) & X"000" & X"1") & eclat_resize(argument2,16));
                        state_var3000 <= make_block;
                      end if;
                    when others =>
                      eclat_print_string(of_string("unknown opcode : "));
                      
                      \$code_ptr\ <= to_integer(unsigned(\$v522\(0 to 15)));
                      state_var3000 <= pause_getI2976;
                    end case;
                  when pause_getII2983 =>
                    argument2 := \$code_value\;
                    \$v2981\ := eclat_resize(\$v259\,8);
                    case \$v2981\ is
                    when X"24" =>
                      w_arg := X"000" & X"1" & \$v522\(48 to 63) & eclat_resize(argument1,16) & eclat_resize(argument2,16);
                      state_var3000 <= w;
                    when X"2b" =>
                      \$v2946\ := eclat_gt(eclat_resize(argument1,16) & X"000" & X"0");
                      if \$v2946\(0) = '1' then
                        \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                        \$ram_write_request\ <= '1';
                        \$ram_write\ <= \$v522\(16 to 47);
                        state_var3000 <= pause_setI2945;
                      else
                        \$55_sp\ := \$v522\(48 to 63);
                        make_block_id := X"0" & X"47";
                        make_block_arg := \$55_sp\ & \$v522\(16 to 47) & \$v522\(64 to 95) & X"f7" & eclat_add(eclat_resize(argument1,16) & X"000" & X"1");
                        state_var3000 <= make_block;
                      end if;
                    when X"37" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_add(X"3e80" & eclat_resize(argument1,16))));
                      state_var3000 <= pause_getI2949;
                    when X"38" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(16 to 47);
                      state_var3000 <= pause_setI2955;
                    when X"3e" =>
                      make_block_id := X"0" & X"49";
                      make_block_arg := \$v522\(48 to 63) & \$v522\(16 to 47) & \$v522\(64 to 95) & eclat_resize(argument2,8) & eclat_resize(argument1,16);
                      state_var3000 <= make_block;
                    when X"83" =>
                      compbranch_arg := X"0000000" & X"0" & argument1 & argument2 & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= compbranch;
                    when X"84" =>
                      compbranch_arg := X"0000000" & X"1" & argument1 & argument2 & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= compbranch;
                    when X"85" =>
                      compbranch_arg := X"0000000" & X"2" & argument1 & argument2 & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= compbranch;
                    when X"86" =>
                      compbranch_arg := X"0000000" & X"3" & argument1 & argument2 & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= compbranch;
                    when X"87" =>
                      compbranch_arg := X"0000000" & X"4" & argument1 & argument2 & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= compbranch;
                    when X"88" =>
                      compbranch_arg := X"0000000" & X"5" & argument1 & argument2 & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= compbranch;
                    when others =>
                      \$code_ptr\ <= to_integer(unsigned(eclat_add(\$v522\(0 to 15) & X"000" & X"3")));
                      state_var3000 <= pause_getI2979;
                    end case;
                  when pause_getII2986 =>
                    argument1 := \$code_value\;
                    \$v2984\ := eclat_resize(\$v259\,8);
                    case \$v2984\ is
                    when X"0" & X"8" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$v522\(48 to 63) & eclat_resize(argument1,16)) & X"000" & X"1")));
                      state_var3000 <= pause_getI2830;
                    when X"12" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(16 to 47);
                      state_var3000 <= pause_setI2834;
                    when X"13" =>
                      result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"2") & \$v522\(16 to 47) & eclat_sub(\$v522\(48 to 63) & eclat_resize(argument1,16)) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    when X"14" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$v522\(48 to 63) & X"000" & X"1") & eclat_resize(argument1,16))));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(16 to 47);
                      state_var3000 <= pause_setI2835;
                    when X"19" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v522\(64 to 94),16) & eclat_sub(eclat_resize(argument1,16) & X"000" & X"1")) & X"000" & X"1")));
                      state_var3000 <= pause_getI2836;
                    when X"1e" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(16 to 47);
                      state_var3000 <= pause_setI2840;
                    when X"1f" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= eclat_resize(\$v522\(96 to 103),31) & eclat_true;
                      state_var3000 <= pause_setI2843;
                    when X"20" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v522\(16 to 46),16) & X"000" & X"0") & X"000" & X"1")));
                      state_var3000 <= pause_getI2844;
                    when X"25" =>
                      apply_arg := eclat_true & eclat_false & eclat_false & \$v522\(96 to 103) & eclat_true & eclat_resize(argument1,16) & X"000" & X"1" & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 95) & \$v522\(96 to 103) & \$v522\(104 to 119) & \$v522\(120 to 121);
                      state_var3000 <= apply;
                    when X"26" =>
                      apply_arg := eclat_true & eclat_true & eclat_false & eclat_add(\$v522\(96 to 103) & X"0" & X"1") & eclat_true & eclat_resize(argument1,16) & X"000" & X"2" & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 95) & \$v522\(96 to 103) & \$v522\(104 to 119) & \$v522\(120 to 121);
                      state_var3000 <= apply;
                    when X"27" =>
                      apply_arg := eclat_true & eclat_true & eclat_true & eclat_add(\$v522\(96 to 103) & X"0" & X"2") & eclat_true & eclat_resize(argument1,16) & X"000" & X"3" & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 95) & \$v522\(96 to 103) & \$v522\(104 to 119) & \$v522\(120 to 121);
                      state_var3000 <= apply;
                    when X"28" =>
                      \$v2854\ := eclat_gt(\$v522\(96 to 103) & X"0" & X"0");
                      if \$v2854\(0) = '1' then
                        \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v522\(16 to 46),16) & X"000" & X"0") & X"000" & X"1")));
                        state_var3000 <= pause_getI2846;
                      else
                        \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$v522\(48 to 63) & eclat_resize(argument1,16)) & X"000" & X"1")));
                        state_var3000 <= pause_getI2852;
                      end if;
                    when X"2a" =>
                      \$v2867\ := eclat_ge(\$v522\(96 to 103) & eclat_resize(argument1,8));
                      if \$v2867\(0) = '1' then
                        result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"2") & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 95) & eclat_sub(\$v522\(96 to 103) & eclat_resize(argument1,8)) & \$v522\(104 to 119) & \$v522\(120 to 121);
                        rdy2583 := eclat_true;
                        state_var3000 <= compute2584;
                      else
                        make_block_id := X"0" & X"38";
                        make_block_arg := \$v522\(48 to 63) & \$v522\(16 to 47) & \$v522\(64 to 95) & X"f7" & eclat_resize(eclat_add(\$v522\(96 to 103) & X"0" & X"3"),16);
                        state_var3000 <= make_block;
                      end if;
                    when X"30" =>
                      offsetclosure_n_arg := eclat_add(\$v522\(0 to 15) & X"000" & X"2") & \$v522\(48 to 63) & eclat_resize(argument1,16) & \$v522\(64 to 95) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= offsetclosure_n;
                    when X"34" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(16 to 47);
                      state_var3000 <= pause_setI2868;
                    when X"35" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_add(X"3e80" & eclat_resize(argument1,16))));
                      state_var3000 <= pause_getI2869;
                    when X"36" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(16 to 47);
                      state_var3000 <= pause_setI2873;
                    when X"39" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(X"3e80" & eclat_resize(argument1,16))));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(16 to 47);
                      state_var3000 <= pause_setI2874;
                    when X"3b" =>
                      make_block_n_arg := eclat_add(\$v522\(0 to 15) & X"000" & X"2") & \$v522\(48 to 63) & eclat_false & eclat_false & eclat_false & argument1 & X"000" & X"0" & \$v522\(16 to 47) & \$v522\(64 to 95) & \$v522\(96 to 103) & \$v522\(104 to 119) & \$v522\(120 to 121);
                      state_var3000 <= make_block_n;
                    when X"3d" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(16 to 47);
                      state_var3000 <= pause_setI2875;
                    when X"3f" =>
                      make_block_n_arg := eclat_add(\$v522\(0 to 15) & X"000" & X"2") & \$v522\(48 to 63) & eclat_true & eclat_false & eclat_false & argument1 & X"000" & X"1" & \$v522\(16 to 47) & \$v522\(64 to 95) & \$v522\(96 to 103) & \$v522\(104 to 119) & \$v522\(120 to 121);
                      state_var3000 <= make_block_n;
                    when X"40" =>
                      make_block_n_arg := eclat_add(\$v522\(0 to 15) & X"000" & X"2") & \$v522\(48 to 63) & eclat_true & eclat_true & eclat_false & argument1 & X"000" & X"2" & \$v522\(16 to 47) & \$v522\(64 to 95) & \$v522\(96 to 103) & \$v522\(104 to 119) & \$v522\(120 to 121);
                      state_var3000 <= make_block_n;
                    when X"41" =>
                      make_block_n_arg := eclat_add(\$v522\(0 to 15) & X"000" & X"2") & \$v522\(48 to 63) & eclat_true & eclat_true & eclat_true & argument1 & X"000" & X"3" & \$v522\(16 to 47) & \$v522\(64 to 95) & \$v522\(96 to 103) & \$v522\(104 to 119) & \$v522\(120 to 121);
                      state_var3000 <= make_block_n;
                    when X"42" =>
                      eclat_print_string(of_string("fatal error: "));
                      
                      eclat_print_string(of_string("unsupported instruction SETFLOATFIELD"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      state_var3000 <= forever;
                    when X"47" =>
                      assert eclat_not(""&\$v522\(47)) = eclat_true report "assertion failed" severity error;
                      
                      \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v522\(16 to 46),16) & eclat_resize(argument1,16)) & X"000" & X"1")));
                      state_var3000 <= pause_getI2876;
                    when X"4d" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v522\(48 to 63) & X"000" & X"1")));
                      state_var3000 <= pause_getI2879;
                    when X"4e" =>
                      eclat_print_string(of_string("fatal error: "));
                      
                      eclat_print_string(of_string("unsupported instruction SETFLOATFIELD"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      state_var3000 <= \$855_forever\;
                    when X"57" =>
                      \$v2885\ := ""&\$v522\(47);
                      if \$v2885\(0) = '1' then
                        \$125_ofs\ := eclat_resize(\$v522\(16 to 46),16);
                        \$code_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(\$v522\(0 to 15) & X"000" & X"2") & \$125_ofs\)));
                        state_var3000 <= pause_getI2881;
                      else
                        \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$v522\(16 to 46),16)));
                        state_var3000 <= pause_getI2883;
                      end if;
                    when X"54" =>
                      result2582 := eclat_add(eclat_add(\$v522\(0 to 15) & X"000" & X"1") & eclat_resize(argument1,16)) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    when X"59" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= eclat_resize(\$v522\(96 to 103),31) & eclat_true;
                      state_var3000 <= pause_setI2889;
                    when X"5c" =>
                      result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 95) & \$v522\(96 to 103) & \$v522\(104 to 119) & \$v522\(120 to 121);
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    when X"5d" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(64 to 95);
                      state_var3000 <= pause_setI2893;
                    when X"5e" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v522\(48 to 63) & X"000" & X"1")));
                      state_var3000 <= pause_getI2898;
                    when X"5f" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v522\(48 to 63) & X"000" & X"1")));
                      state_var3000 <= pause_getI2906;
                    when X"60" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v522\(48 to 63) & X"000" & X"1")));
                      state_var3000 <= pause_getI2916;
                    when X"61" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v522\(48 to 63) & X"000" & X"1")));
                      state_var3000 <= pause_getI2928;
                    when X"62" =>
                      eclat_print_string(of_string("fatal error: "));
                      
                      eclat_print_string(of_string("unsupported instruction CALLN"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      state_var3000 <= \$921_forever\;
                    when X"67" =>
                      result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"2") & argument1 & eclat_true & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    when X"6c" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(16 to 47);
                      state_var3000 <= pause_setI2930;
                    when X"7f" =>
                      result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"2") & eclat_add(\$v522\(16 to 46) & argument1) & eclat_true & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    when X"80" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v522\(16 to 46),16) & X"000" & X"0") & X"000" & X"1")));
                      state_var3000 <= pause_getI2932;
                    when X"8b" =>
                      compbranch_arg := X"0000000" & X"2" & argument1 & \$v522\(16 to 46) & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= compbranch;
                    when X"8c" =>
                      compbranch_arg := X"0000000" & X"5" & argument1 & \$v522\(16 to 46) & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= compbranch;
                    when others =>
                      \$code_ptr\ <= to_integer(unsigned(eclat_add(\$v522\(0 to 15) & X"000" & X"2")));
                      state_var3000 <= pause_getI2982;
                    end case;
                  when pause_getII2989 =>
                    \$v259\ := \$code_value\;
                    \$v2987\ := eclat_resize(\$v259\,8);
                    case \$v2987\ is
                    when X"0" & X"0" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$v522\(48 to 63) & X"000" & X"0") & X"000" & X"1")));
                      state_var3000 <= pause_getI2705;
                    when X"0" & X"1" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$v522\(48 to 63) & X"000" & X"1") & X"000" & X"1")));
                      state_var3000 <= pause_getI2707;
                    when X"0" & X"2" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$v522\(48 to 63) & X"000" & X"2") & X"000" & X"1")));
                      state_var3000 <= pause_getI2709;
                    when X"0" & X"3" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$v522\(48 to 63) & X"000" & X"3") & X"000" & X"1")));
                      state_var3000 <= pause_getI2711;
                    when X"0" & X"4" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$v522\(48 to 63) & X"000" & X"4") & X"000" & X"1")));
                      state_var3000 <= pause_getI2713;
                    when X"0" & X"5" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$v522\(48 to 63) & X"000" & X"5") & X"000" & X"1")));
                      state_var3000 <= pause_getI2715;
                    when X"0" & X"6" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$v522\(48 to 63) & X"000" & X"6") & X"000" & X"1")));
                      state_var3000 <= pause_getI2717;
                    when X"0" & X"7" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$v522\(48 to 63) & X"000" & X"7") & X"000" & X"1")));
                      state_var3000 <= pause_getI2719;
                    when X"0" & X"9" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(16 to 47);
                      state_var3000 <= pause_setI2721;
                    when X"0" & X"a" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(16 to 47);
                      state_var3000 <= pause_setI2722;
                    when X"0" & X"b" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(16 to 47);
                      state_var3000 <= pause_setI2725;
                    when X"0" & X"c" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(16 to 47);
                      state_var3000 <= pause_setI2728;
                    when X"0" & X"d" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(16 to 47);
                      state_var3000 <= pause_setI2731;
                    when X"0" & X"e" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(16 to 47);
                      state_var3000 <= pause_setI2734;
                    when X"0" & X"f" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(16 to 47);
                      state_var3000 <= pause_setI2737;
                    when X"10" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(16 to 47);
                      state_var3000 <= pause_setI2740;
                    when X"11" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(16 to 47);
                      state_var3000 <= pause_setI2743;
                    when X"15" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v522\(64 to 94),16) & eclat_sub(X"000" & X"1" & X"000" & X"1")) & X"000" & X"1")));
                      state_var3000 <= pause_getI2744;
                    when X"16" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v522\(64 to 94),16) & eclat_sub(X"000" & X"2" & X"000" & X"1")) & X"000" & X"1")));
                      state_var3000 <= pause_getI2746;
                    when X"17" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v522\(64 to 94),16) & eclat_sub(X"000" & X"3" & X"000" & X"1")) & X"000" & X"1")));
                      state_var3000 <= pause_getI2748;
                    when X"18" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v522\(64 to 94),16) & eclat_sub(X"000" & X"4" & X"000" & X"1")) & X"000" & X"1")));
                      state_var3000 <= pause_getI2750;
                    when X"1a" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(16 to 47);
                      state_var3000 <= pause_setI2754;
                    when X"1b" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(16 to 47);
                      state_var3000 <= pause_setI2757;
                    when X"1c" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(16 to 47);
                      state_var3000 <= pause_setI2760;
                    when X"1d" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(16 to 47);
                      state_var3000 <= pause_setI2763;
                    when X"21" =>
                      apply_arg := eclat_true & eclat_false & eclat_false & X"0" & X"0" & eclat_false & X"000" & X"0" & X"000" & X"0" & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 95) & \$v522\(96 to 103) & \$v522\(104 to 119) & \$v522\(120 to 121);
                      state_var3000 <= apply;
                    when X"22" =>
                      apply_arg := eclat_true & eclat_true & eclat_false & X"0" & X"1" & eclat_false & X"000" & X"0" & X"000" & X"0" & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 95) & \$v522\(96 to 103) & \$v522\(104 to 119) & \$v522\(120 to 121);
                      state_var3000 <= apply;
                    when X"23" =>
                      apply_arg := eclat_true & eclat_true & eclat_true & X"0" & X"2" & eclat_false & X"000" & X"0" & X"000" & X"0" & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 95) & \$v522\(96 to 103) & \$v522\(104 to 119) & \$v522\(120 to 121);
                      state_var3000 <= apply;
                    when X"29" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$v522\(64 to 94),16)));
                      state_var3000 <= pause_getI2770;
                    when X"2d" =>
                      offsetclosure_n_arg := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$v522\(48 to 63) & eclat_sub(X"000" & X"0" & X"000" & X"2") & \$v522\(64 to 95) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= offsetclosure_n;
                    when X"2e" =>
                      offsetclosure_n_arg := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$v522\(48 to 63) & X"000" & X"0" & \$v522\(64 to 95) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= offsetclosure_n;
                    when X"2f" =>
                      offsetclosure_n_arg := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$v522\(48 to 63) & X"000" & X"2" & \$v522\(64 to 95) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= offsetclosure_n;
                    when X"31" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(16 to 47);
                      state_var3000 <= pause_setI2772;
                    when X"32" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(16 to 47);
                      state_var3000 <= pause_setI2773;
                    when X"33" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(16 to 47);
                      state_var3000 <= pause_setI2774;
                    when X"3a" =>
                      make_block_n_arg := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$v522\(48 to 63) & eclat_false & eclat_false & eclat_false & "000"& X"000000" & X"0" & X"000" & X"0" & \$v522\(16 to 47) & \$v522\(64 to 95) & \$v522\(96 to 103) & \$v522\(104 to 119) & \$v522\(120 to 121);
                      state_var3000 <= make_block_n;
                    when X"3c" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(16 to 47);
                      state_var3000 <= pause_setI2775;
                    when X"43" =>
                      assert eclat_not(""&\$v522\(47)) = eclat_true report "assertion failed" severity error;
                      
                      \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v522\(16 to 46),16) & X"000" & X"0") & X"000" & X"1")));
                      state_var3000 <= pause_getI2776;
                    when X"44" =>
                      assert eclat_not(""&\$v522\(47)) = eclat_true report "assertion failed" severity error;
                      
                      \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v522\(16 to 46),16) & X"000" & X"1") & X"000" & X"1")));
                      state_var3000 <= pause_getI2778;
                    when X"45" =>
                      assert eclat_not(""&\$v522\(47)) = eclat_true report "assertion failed" severity error;
                      
                      \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v522\(16 to 46),16) & X"000" & X"2") & X"000" & X"1")));
                      state_var3000 <= pause_getI2780;
                    when X"46" =>
                      assert eclat_not(""&\$v522\(47)) = eclat_true report "assertion failed" severity error;
                      
                      \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v522\(16 to 46),16) & X"000" & X"3") & X"000" & X"1")));
                      state_var3000 <= pause_getI2782;
                    when X"49" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v522\(48 to 63) & X"000" & X"1")));
                      state_var3000 <= pause_getI2785;
                    when X"4a" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v522\(48 to 63) & X"000" & X"1")));
                      state_var3000 <= pause_getI2788;
                    when X"4b" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v522\(48 to 63) & X"000" & X"1")));
                      state_var3000 <= pause_getI2791;
                    when X"4c" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v522\(48 to 63) & X"000" & X"1")));
                      state_var3000 <= pause_getI2794;
                    when X"4f" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$v522\(16 to 46),16)));
                      state_var3000 <= pause_getI2796;
                    when X"50" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v522\(48 to 63) & X"000" & X"1")));
                      state_var3000 <= pause_getI2800;
                    when X"51" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v522\(48 to 63) & X"000" & X"1")));
                      state_var3000 <= pause_getI2805;
                    when X"52" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v522\(48 to 63) & X"000" & X"1")));
                      state_var3000 <= pause_getI2809;
                    when X"53" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v522\(48 to 63) & X"000" & X"1")));
                      state_var3000 <= pause_getI2814;
                    when X"55" =>
                      branch_if_arg := eclat_false & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= branch_if;
                    when X"56" =>
                      branch_if_arg := eclat_true & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= branch_if;
                    when X"58" =>
                      result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & 
                      eclat_if(eclat_eq(\$v522\(16 to 46) & "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    when X"5a" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$v522\(48 to 63) & X"000" & X"1") & X"000" & X"1")));
                      state_var3000 <= pause_getI2816;
                    when X"5b" =>
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v522\(104 to 119) & X"000" & X"1")));
                      state_var3000 <= pause_getI2824;
                    when X"63" =>
                      result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"0" & eclat_true & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    when X"64" =>
                      result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    when X"65" =>
                      result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"2" & eclat_true & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    when X"66" =>
                      result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"3" & eclat_true & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    when X"68" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(16 to 47);
                      state_var3000 <= pause_setI2826;
                    when X"69" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(16 to 47);
                      state_var3000 <= pause_setI2827;
                    when X"6a" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(16 to 47);
                      state_var3000 <= pause_setI2828;
                    when X"6b" =>
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v522\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v522\(16 to 47);
                      state_var3000 <= pause_setI2829;
                    when X"6e" =>
                      binop_int_arg := X"0000000" & X"0" & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= binop_int;
                    when X"6f" =>
                      binop_int_arg := X"0000000" & X"1" & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= binop_int;
                    when X"70" =>
                      binop_int_arg := X"0000000" & X"2" & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= binop_int;
                    when X"71" =>
                      binop_int_arg := X"0000000" & X"3" & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= binop_int;
                    when X"72" =>
                      binop_int_arg := X"0000000" & X"4" & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= binop_int;
                    when X"73" =>
                      binop_int_arg := X"0000000" & X"5" & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= binop_int;
                    when X"74" =>
                      binop_int_arg := X"0000000" & X"6" & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= binop_int;
                    when X"75" =>
                      binop_int_arg := X"0000000" & X"7" & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= binop_int;
                    when X"76" =>
                      binop_int_arg := X"0000000" & X"8" & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= binop_int;
                    when X"77" =>
                      binop_int_arg := X"0000000" & X"9" & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= binop_int;
                    when X"78" =>
                      binop_int_arg := X"0000000" & X"a" & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= binop_int;
                    when X"82" =>
                      eclat_print_string(of_string("fatal error: "));
                      
                      eclat_print_string(of_string("unsupported instruction GETMETHOD"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      state_var3000 <= \$1278_forever\;
                    when X"89" =>
                      binop_int_arg := X"0000000" & X"b" & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= binop_int;
                    when X"8a" =>
                      binop_int_arg := X"0000000" & X"c" & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= binop_int;
                    when X"8d" =>
                      eclat_print_string(of_string("fatal error: "));
                      
                      eclat_print_string(of_string("unsupported instruction GETPUBMET"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      state_var3000 <= \$1281_forever\;
                    when X"8e" =>
                      eclat_print_string(of_string("fatal error: "));
                      
                      eclat_print_string(of_string("unsupported instruction GETDYNMET"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      state_var3000 <= \$1284_forever\;
                    when X"79" =>
                      binop_compare_arg := X"0000000" & X"0" & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= binop_compare;
                    when X"7a" =>
                      binop_compare_arg := X"0000000" & X"1" & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= binop_compare;
                    when X"7b" =>
                      binop_compare_arg := X"0000000" & X"2" & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= binop_compare;
                    when X"7c" =>
                      binop_compare_arg := X"0000000" & X"3" & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= binop_compare;
                    when X"7d" =>
                      binop_compare_arg := X"0000000" & X"4" & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= binop_compare;
                    when X"7e" =>
                      binop_compare_arg := X"0000000" & X"5" & \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      state_var3000 <= binop_compare;
                    when X"81" =>
                      result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & 
                      eclat_if(""&\$v522\(47) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    when X"8f" =>
                      eclat_print_string(of_string("STOP : "));
                      
                      result2582 := \$v522\(0 to 15) & \$v522\(16 to 47) & \$v522\(48 to 63) & \$v522\(64 to 119) & eclat_true & ""&\$v522\(121);
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    when others =>
                      \$code_ptr\ <= to_integer(unsigned(eclat_add(\$v522\(0 to 15) & X"000" & X"1")));
                      state_var3000 <= pause_getI2985;
                    end case;
                  when pause_setI2585 =>
                    \$ram_write_request\ <= '0';
                    make_block_result := \$v1380\(0 to 31) & \$v1380\(32 to 63) & eclat_resize(\$v1380\(64 to 79),31) & eclat_false;
                    case make_block_id is
                    when X"00" & X"e" =>
                      \$v866\ := make_block_result;
                      \$v2701\ := ""&make_block_n_arg(32);
                      if \$v2701\(0) = '1' then
                        \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v866\(64 to 94),16) & X"000" & X"0") & X"000" & X"1")));
                        \$ram_write_request\ <= '1';
                        \$ram_write\ <= \$v866\(0 to 31);
                        state_var3000 <= pause_setI2700;
                      else
                        \$v2699\ := ""&make_block_n_arg(33);
                        if \$v2699\(0) = '1' then
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(make_block_n_arg(16 to 31) & X"000" & X"1")));
                          state_var3000 <= pause_getI2697;
                        else
                          \$288_sp\ := make_block_n_arg(16 to 31);
                          \$v2695\ := ""&make_block_n_arg(34);
                          if \$v2695\(0) = '1' then
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$288_sp\ & X"000" & X"1")));
                            state_var3000 <= pause_getI2693;
                          else
                            \$289_sp\ := \$288_sp\;
                            make_block_n_result := make_block_n_arg(0 to 15) & \$v866\(64 to 95) & \$289_sp\ & \$v866\(32 to 63) & make_block_n_arg(146 to 153) & make_block_n_arg(154 to 169) & make_block_n_arg(170 to 171);
                            result2582 := make_block_n_result;
                            rdy2583 := eclat_true;
                            state_var3000 <= compute2584;
                          end if;
                        end if;
                      end if;
                    when X"0" & X"38" =>
                      \$v620\ := make_block_result;
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v620\(64 to 94),16) & X"000" & X"0") & X"000" & X"1")));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= eclat_resize(eclat_sub(eclat_add(\$v522\(0 to 15) & X"000" & X"2") & X"000" & X"3"),31) & eclat_true;
                      state_var3000 <= pause_setI2866;
                    when X"0" & X"47" =>
                      \$v584\ := make_block_result;
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v584\(64 to 94),16) & X"000" & X"0") & X"000" & X"1")));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= eclat_resize(eclat_add(eclat_add(\$v522\(0 to 15) & X"000" & X"2") & eclat_resize(argument2,16)),31) & eclat_true;
                      state_var3000 <= pause_setI2944;
                    when X"0" & X"49" =>
                      \$v593\ := make_block_result;
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v593\(64 to 94),16) & X"000" & X"0") & X"000" & X"1")));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v593\(0 to 31);
                      state_var3000 <= pause_setI2960;
                    when X"0" & X"53" =>
                      \$v540\ := make_block_result;
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v540\(64 to 94),16) & X"000" & X"0") & X"000" & X"1")));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= eclat_resize(eclat_add(eclat_add(\$v522\(0 to 15) & X"000" & X"3") & eclat_resize(argument3,16)),31) & eclat_true;
                      state_var3000 <= pause_setI2973;
                    when others =>
                      
                    end case;
                  when pause_setI2662 =>
                    \$ram_write_request\ <= '0';
                    \$342_sp\ := eclat_add(\$341_sp\ & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(apply_arg(60 to 90),16) & X"000" & X"0") & X"000" & X"1")));
                    state_var3000 <= pause_getI2660;
                  when pause_setI2664 =>
                    \$ram_write_request\ <= '0';
                    \$341_sp\ := eclat_add(\$340_sp\ & X"000" & X"1");
                    \$v2663\ := ""&apply_arg(0);
                    if \$v2663\(0) = '1' then
                      \$ram_ptr_write\ <= to_integer(unsigned(\$341_sp\));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v906\(0 to 31);
                      state_var3000 <= pause_setI2662;
                    else
                      \$342_sp\ := \$341_sp\;
                      \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(apply_arg(60 to 90),16) & X"000" & X"0") & X"000" & X"1")));
                      state_var3000 <= pause_getI2660;
                    end if;
                  when pause_setI2666 =>
                    \$ram_write_request\ <= '0';
                    \$340_sp\ := eclat_add(\$339_sp\ & X"000" & X"1");
                    \$v2665\ := ""&apply_arg(1);
                    if \$v2665\(0) = '1' then
                      \$ram_ptr_write\ <= to_integer(unsigned(\$340_sp\));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v907\(0 to 31);
                      state_var3000 <= pause_setI2664;
                    else
                      \$341_sp\ := \$340_sp\;
                      \$v2663\ := ""&apply_arg(0);
                      if \$v2663\(0) = '1' then
                        \$ram_ptr_write\ <= to_integer(unsigned(\$341_sp\));
                        \$ram_write_request\ <= '1';
                        \$ram_write\ <= \$v906\(0 to 31);
                        state_var3000 <= pause_setI2662;
                      else
                        \$342_sp\ := \$341_sp\;
                        \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(apply_arg(60 to 90),16) & X"000" & X"0") & X"000" & X"1")));
                        state_var3000 <= pause_getI2660;
                      end if;
                    end if;
                  when pause_setI2668 =>
                    \$ram_write_request\ <= '0';
                    \$347_sp\ := eclat_add(\$346_sp\ & X"000" & X"1");
                    \$339_sp\ := \$347_sp\;
                    \$v2667\ := ""&apply_arg(2);
                    if \$v2667\(0) = '1' then
                      \$ram_ptr_write\ <= to_integer(unsigned(\$339_sp\));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v908\(0 to 31);
                      state_var3000 <= pause_setI2666;
                    else
                      \$340_sp\ := \$339_sp\;
                      \$v2665\ := ""&apply_arg(1);
                      if \$v2665\(0) = '1' then
                        \$ram_ptr_write\ <= to_integer(unsigned(\$340_sp\));
                        \$ram_write_request\ <= '1';
                        \$ram_write\ <= \$v907\(0 to 31);
                        state_var3000 <= pause_setI2664;
                      else
                        \$341_sp\ := \$340_sp\;
                        \$v2663\ := ""&apply_arg(0);
                        if \$v2663\(0) = '1' then
                          \$ram_ptr_write\ <= to_integer(unsigned(\$341_sp\));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$v906\(0 to 31);
                          state_var3000 <= pause_setI2662;
                        else
                          \$342_sp\ := \$341_sp\;
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(apply_arg(60 to 90),16) & X"000" & X"0") & X"000" & X"1")));
                          state_var3000 <= pause_getI2660;
                        end if;
                      end if;
                    end if;
                  when pause_setI2669 =>
                    \$ram_write_request\ <= '0';
                    \$346_sp\ := eclat_add(\$345_sp\ & X"000" & X"1");
                    \$ram_ptr_write\ <= to_integer(unsigned(\$346_sp\));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= eclat_resize(eclat_add(apply_arg(44 to 59) & X"000" & X"1"),31) & eclat_true;
                    state_var3000 <= pause_setI2668;
                  when pause_setI2670 =>
                    \$ram_write_request\ <= '0';
                    \$345_sp\ := eclat_add(\$v908\(32 to 47) & X"000" & X"1");
                    \$ram_ptr_write\ <= to_integer(unsigned(\$345_sp\));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= apply_arg(108 to 139);
                    state_var3000 <= pause_setI2669;
                  when pause_setI2692 =>
                    \$ram_write_request\ <= '0';
                    \$289_sp\ := \$v868\(32 to 47);
                    make_block_n_result := make_block_n_arg(0 to 15) & \$v866\(64 to 95) & \$289_sp\ & \$v866\(32 to 63) & make_block_n_arg(146 to 153) & make_block_n_arg(154 to 169) & make_block_n_arg(170 to 171);
                    result2582 := make_block_n_result;
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_setI2696 =>
                    \$ram_write_request\ <= '0';
                    \$288_sp\ := \$v871\(32 to 47);
                    \$v2695\ := ""&make_block_n_arg(34);
                    if \$v2695\(0) = '1' then
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$288_sp\ & X"000" & X"1")));
                      state_var3000 <= pause_getI2693;
                    else
                      \$289_sp\ := \$288_sp\;
                      make_block_n_result := make_block_n_arg(0 to 15) & \$v866\(64 to 95) & \$289_sp\ & \$v866\(32 to 63) & make_block_n_arg(146 to 153) & make_block_n_arg(154 to 169) & make_block_n_arg(170 to 171);
                      result2582 := make_block_n_result;
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    end if;
                  when pause_setI2700 =>
                    \$ram_write_request\ <= '0';
                    \$v2699\ := ""&make_block_n_arg(33);
                    if \$v2699\(0) = '1' then
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(make_block_n_arg(16 to 31) & X"000" & X"1")));
                      state_var3000 <= pause_getI2697;
                    else
                      \$288_sp\ := make_block_n_arg(16 to 31);
                      \$v2695\ := ""&make_block_n_arg(34);
                      if \$v2695\(0) = '1' then
                        \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$288_sp\ & X"000" & X"1")));
                        state_var3000 <= pause_getI2693;
                      else
                        \$289_sp\ := \$288_sp\;
                        make_block_n_result := make_block_n_arg(0 to 15) & \$v866\(64 to 95) & \$289_sp\ & \$v866\(32 to 63) & make_block_n_arg(146 to 153) & make_block_n_arg(154 to 169) & make_block_n_arg(170 to 171);
                        result2582 := make_block_n_result;
                        rdy2583 := eclat_true;
                        state_var3000 <= compute2584;
                      end if;
                    end if;
                  when pause_setI2721 =>
                    \$ram_write_request\ <= '0';
                    \$364_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$v522\(16 to 47) & \$364_sp\ & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_setI2722 =>
                    \$ram_write_request\ <= '0';
                    \$981_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$v522\(16 to 47) & \$981_sp\ & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_setI2725 =>
                    \$ram_write_request\ <= '0';
                    \$983_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$983_sp\ & X"000" & X"1") & X"000" & X"1")));
                    state_var3000 <= pause_getI2723;
                  when pause_setI2728 =>
                    \$ram_write_request\ <= '0';
                    \$988_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$988_sp\ & X"000" & X"2") & X"000" & X"1")));
                    state_var3000 <= pause_getI2726;
                  when pause_setI2731 =>
                    \$ram_write_request\ <= '0';
                    \$993_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$993_sp\ & X"000" & X"3") & X"000" & X"1")));
                    state_var3000 <= pause_getI2729;
                  when pause_setI2734 =>
                    \$ram_write_request\ <= '0';
                    \$998_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$998_sp\ & X"000" & X"4") & X"000" & X"1")));
                    state_var3000 <= pause_getI2732;
                  when pause_setI2737 =>
                    \$ram_write_request\ <= '0';
                    \$1003_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$1003_sp\ & X"000" & X"5") & X"000" & X"1")));
                    state_var3000 <= pause_getI2735;
                  when pause_setI2740 =>
                    \$ram_write_request\ <= '0';
                    \$1008_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$1008_sp\ & X"000" & X"6") & X"000" & X"1")));
                    state_var3000 <= pause_getI2738;
                  when pause_setI2743 =>
                    \$ram_write_request\ <= '0';
                    \$1013_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$1013_sp\ & X"000" & X"7") & X"000" & X"1")));
                    state_var3000 <= pause_getI2741;
                  when pause_setI2754 =>
                    \$ram_write_request\ <= '0';
                    \$1048_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v522\(64 to 94),16) & eclat_sub(X"000" & X"1" & X"000" & X"1")) & X"000" & X"1")));
                    state_var3000 <= pause_getI2752;
                  when pause_setI2757 =>
                    \$ram_write_request\ <= '0';
                    \$1057_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v522\(64 to 94),16) & eclat_sub(X"000" & X"2" & X"000" & X"1")) & X"000" & X"1")));
                    state_var3000 <= pause_getI2755;
                  when pause_setI2760 =>
                    \$ram_write_request\ <= '0';
                    \$1066_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v522\(64 to 94),16) & eclat_sub(X"000" & X"3" & X"000" & X"1")) & X"000" & X"1")));
                    state_var3000 <= pause_getI2758;
                  when pause_setI2763 =>
                    \$ram_write_request\ <= '0';
                    \$1075_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v522\(64 to 94),16) & eclat_sub(X"000" & X"4" & X"000" & X"1")) & X"000" & X"1")));
                    state_var3000 <= pause_getI2761;
                  when pause_setI2764 =>
                    \$ram_write_request\ <= '0';
                    \$241_sp\ := eclat_add(loop_push_arg(0 to 15) & X"000" & X"1");
                    loop_push_arg := \$241_sp\ & eclat_add(loop_push_arg(16 to 23) & X"0" & X"1") & loop_push_arg(24 to 55) & loop_push_arg(56 to 63);
                    state_var3000 <= loop_push;
                  when pause_setI2772 =>
                    \$ram_write_request\ <= '0';
                    \$1100_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    offsetclosure_n_arg := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$1100_sp\ & eclat_sub(X"000" & X"0" & X"000" & X"2") & \$v522\(64 to 95) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    state_var3000 <= offsetclosure_n;
                  when pause_setI2773 =>
                    \$ram_write_request\ <= '0';
                    \$1103_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    offsetclosure_n_arg := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$1103_sp\ & X"000" & X"0" & \$v522\(64 to 95) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    state_var3000 <= offsetclosure_n;
                  when pause_setI2774 =>
                    \$ram_write_request\ <= '0';
                    \$1106_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    offsetclosure_n_arg := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$1106_sp\ & X"000" & X"2" & \$v522\(64 to 95) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    state_var3000 <= offsetclosure_n;
                  when pause_setI2775 =>
                    \$ram_write_request\ <= '0';
                    \$242_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    make_block_n_arg := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & \$242_sp\ & eclat_false & eclat_false & eclat_false & "000"& X"000000" & X"0" & X"000" & X"0" & \$v522\(16 to 47) & \$v522\(64 to 95) & \$v522\(96 to 103) & \$v522\(104 to 119) & \$v522\(120 to 121);
                    state_var3000 <= make_block_n;
                  when pause_setI2784 =>
                    \$ram_write_request\ <= '0';
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & \$v796\(32 to 47) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_setI2787 =>
                    \$ram_write_request\ <= '0';
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & \$v799\(32 to 47) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_setI2790 =>
                    \$ram_write_request\ <= '0';
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & \$v802\(32 to 47) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_setI2793 =>
                    \$ram_write_request\ <= '0';
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & \$v805\(32 to 47) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_setI2802 =>
                    \$ram_write_request\ <= '0';
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & \$v814\(32 to 47) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_setI2811 =>
                    \$ram_write_request\ <= '0';
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & \$v822\(32 to 47) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_setI2826 =>
                    \$ram_write_request\ <= '0';
                    \$1263_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"0" & eclat_true & \$1263_sp\ & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_setI2827 =>
                    \$ram_write_request\ <= '0';
                    \$1267_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & \$1267_sp\ & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_setI2828 =>
                    \$ram_write_request\ <= '0';
                    \$1271_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"2" & eclat_true & \$1271_sp\ & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_setI2829 =>
                    \$ram_write_request\ <= '0';
                    \$1275_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"3" & eclat_true & \$1275_sp\ & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_setI2834 =>
                    \$ram_write_request\ <= '0';
                    \$357_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$357_sp\ & eclat_resize(argument1,16)) & X"000" & X"1")));
                    state_var3000 <= pause_getI2832;
                  when pause_setI2835 =>
                    \$ram_write_request\ <= '0';
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"2") & "000"& X"000000" & X"1" & eclat_true & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_setI2840 =>
                    \$ram_write_request\ <= '0';
                    \$354_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v522\(64 to 94),16) & eclat_sub(eclat_resize(argument1,16) & X"000" & X"1")) & X"000" & X"1")));
                    state_var3000 <= pause_getI2838;
                  when pause_setI2841 =>
                    \$ram_write_request\ <= '0';
                    \$84_sp\ := eclat_add(\$83_sp\ & X"000" & X"1");
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"2") & \$v522\(16 to 47) & \$84_sp\ & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_setI2842 =>
                    \$ram_write_request\ <= '0';
                    \$83_sp\ := eclat_add(\$81_sp\ & X"000" & X"1");
                    \$ram_ptr_write\ <= to_integer(unsigned(\$83_sp\));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= eclat_resize(eclat_add(eclat_add(\$v522\(0 to 15) & X"000" & X"1") & eclat_resize(argument1,16)),31) & eclat_true;
                    state_var3000 <= pause_setI2841;
                  when pause_setI2843 =>
                    \$ram_write_request\ <= '0';
                    \$81_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    \$ram_ptr_write\ <= to_integer(unsigned(\$81_sp\));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v522\(64 to 95);
                    state_var3000 <= pause_setI2842;
                  when pause_setI2855 =>
                    \$ram_write_request\ <= '0';
                    \$103_w_arg\ := eclat_add(\$103_w_arg\(0 to 7) & X"0" & X"1") & \$v632\(32 to 47) & \$103_w_arg\(24 to 55) & \$103_w_arg\(56 to 63);
                    state_var3000 <= \$103_w\;
                  when pause_setI2865 =>
                    \$ram_write_request\ <= '0';
                    \$103_w_arg\ := X"0" & X"0" & \$v522\(48 to 63) & \$v620\(64 to 95) & \$v522\(96 to 103);
                    state_var3000 <= \$103_w\;
                  when pause_setI2866 =>
                    \$ram_write_request\ <= '0';
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v620\(64 to 94),16) & X"000" & X"1") & X"000" & X"1")));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v620\(32 to 63);
                    state_var3000 <= pause_setI2865;
                  when pause_setI2868 =>
                    \$ram_write_request\ <= '0';
                    \$324_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    offsetclosure_n_arg := eclat_add(\$v522\(0 to 15) & X"000" & X"2") & \$324_sp\ & eclat_resize(argument1,16) & \$v522\(64 to 95) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    state_var3000 <= offsetclosure_n;
                  when pause_setI2873 =>
                    \$ram_write_request\ <= '0';
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(X"3e80" & eclat_resize(argument1,16))));
                    state_var3000 <= pause_getI2871;
                  when pause_setI2874 =>
                    \$ram_write_request\ <= '0';
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"2") & "000"& X"000000" & X"1" & eclat_true & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_setI2875 =>
                    \$ram_write_request\ <= '0';
                    \$123_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    make_block_n_arg := eclat_add(\$v522\(0 to 15) & X"000" & X"2") & \$123_sp\ & eclat_false & eclat_false & eclat_false & argument1 & X"000" & X"0" & \$v522\(16 to 47) & \$v522\(64 to 95) & \$v522\(96 to 103) & \$v522\(104 to 119) & \$v522\(120 to 121);
                    state_var3000 <= make_block_n;
                  when pause_setI2878 =>
                    \$ram_write_request\ <= '0';
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"2") & "000"& X"000000" & X"1" & eclat_true & \$v649\(32 to 47) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_setI2886 =>
                    \$ram_write_request\ <= '0';
                    \$131_sp\ := eclat_add(\$130_sp\ & X"000" & X"1");
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"2") & \$v522\(16 to 47) & \$131_sp\ & \$v522\(64 to 95) & \$v522\(96 to 103) & \$131_sp\ & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_setI2887 =>
                    \$ram_write_request\ <= '0';
                    \$130_sp\ := eclat_add(\$128_sp\ & X"000" & X"1");
                    \$ram_ptr_write\ <= to_integer(unsigned(\$130_sp\));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= eclat_resize(eclat_add(eclat_add(\$v522\(0 to 15) & X"000" & X"1") & eclat_resize(argument1,16)),31) & eclat_true;
                    state_var3000 <= pause_setI2886;
                  when pause_setI2888 =>
                    \$ram_write_request\ <= '0';
                    \$128_sp\ := eclat_add(\$127_sp\ & X"000" & X"1");
                    \$ram_ptr_write\ <= to_integer(unsigned(\$128_sp\));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= eclat_resize(\$v522\(104 to 119),31) & eclat_true;
                    state_var3000 <= pause_setI2887;
                  when pause_setI2889 =>
                    \$ram_write_request\ <= '0';
                    \$127_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    \$ram_ptr_write\ <= to_integer(unsigned(\$127_sp\));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v522\(64 to 95);
                    state_var3000 <= pause_setI2888;
                  when pause_setI2893 =>
                    \$ram_write_request\ <= '0';
                    \$133_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    \$v2892\ := argument1;
                    case \$v2892\ is
                    when "000"& X"000000" & X"0" =>
                      eclat_print_string(of_string("======> "));
                      
                      eclat_print_int(\$v522\(16 to 46));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$v665\ := "000"& X"000000" & X"1" & eclat_true & \$v522\(0 to 15) & \$v522\(16 to 47) & \$133_sp\ & \$v522\(64 to 95) & \$v522\(96 to 103) & \$v522\(104 to 119) & \$v522\(120 to 121);
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v665\(80 to 95) & X"000" & X"1")));
                      state_var3000 <= pause_getI2890;
                    when others =>
                      eclat_print_string(of_string("unknown primitive"));
                      
                      \$v665\ := "000"& X"000000" & X"1" & eclat_true & \$v522\(0 to 15) & \$v522\(16 to 47) & \$133_sp\ & \$v522\(64 to 95) & \$v522\(96 to 103) & \$v522\(104 to 119) & \$v522\(120 to 121);
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v665\(80 to 95) & X"000" & X"1")));
                      state_var3000 <= pause_getI2890;
                    end case;
                  when pause_setI2897 =>
                    \$ram_write_request\ <= '0';
                    \$148_sp\ := eclat_add(\$v676\(32 to 47) & X"000" & X"1");
                    \$v2896\ := argument1;
                    case \$v2896\ is
                    when "000"& X"000000" & X"0" =>
                      eclat_print_string(of_string("======> "));
                      
                      eclat_print_int(\$v522\(16 to 46));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$v677\ := "000"& X"000000" & X"1" & eclat_true & \$v522\(0 to 15) & \$v522\(16 to 47) & \$148_sp\ & \$v522\(64 to 95) & \$v522\(96 to 103) & \$v522\(104 to 119) & \$v522\(120 to 121);
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v677\(80 to 95) & X"000" & X"1")));
                      state_var3000 <= pause_getI2894;
                    when others =>
                      eclat_print_string(of_string("unknown primitive"));
                      
                      \$v677\ := "000"& X"000000" & X"1" & eclat_true & \$v522\(0 to 15) & \$v522\(16 to 47) & \$148_sp\ & \$v522\(64 to 95) & \$v522\(96 to 103) & \$v522\(104 to 119) & \$v522\(120 to 121);
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v677\(80 to 95) & X"000" & X"1")));
                      state_var3000 <= pause_getI2894;
                    end case;
                  when pause_setI2903 =>
                    \$ram_write_request\ <= '0';
                    \$166_sp\ := eclat_add(\$v689\(32 to 47) & X"000" & X"1");
                    \$v2902\ := argument1;
                    case \$v2902\ is
                    when "000"& X"000000" & X"0" =>
                      eclat_print_string(of_string("======> "));
                      
                      eclat_print_int(\$v522\(16 to 46));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$v690\ := "000"& X"000000" & X"1" & eclat_true & \$v522\(0 to 15) & \$v522\(16 to 47) & \$166_sp\ & \$v522\(64 to 95) & \$v522\(96 to 103) & \$v522\(104 to 119) & \$v522\(120 to 121);
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v690\(80 to 95) & X"000" & X"1")));
                      state_var3000 <= pause_getI2900;
                    when others =>
                      eclat_print_string(of_string("unknown primitive"));
                      
                      \$v690\ := "000"& X"000000" & X"1" & eclat_true & \$v522\(0 to 15) & \$v522\(16 to 47) & \$166_sp\ & \$v522\(64 to 95) & \$v522\(96 to 103) & \$v522\(104 to 119) & \$v522\(120 to 121);
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v690\(80 to 95) & X"000" & X"1")));
                      state_var3000 <= pause_getI2900;
                    end case;
                  when pause_setI2911 =>
                    \$ram_write_request\ <= '0';
                    \$187_sp\ := eclat_add(\$v703\(32 to 47) & X"000" & X"1");
                    \$v2910\ := argument1;
                    case \$v2910\ is
                    when "000"& X"000000" & X"0" =>
                      eclat_print_string(of_string("======> "));
                      
                      eclat_print_int(\$v522\(16 to 46));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$v704\ := "000"& X"000000" & X"1" & eclat_true & \$v522\(0 to 15) & \$v522\(16 to 47) & \$187_sp\ & \$v522\(64 to 95) & \$v522\(96 to 103) & \$v522\(104 to 119) & \$v522\(120 to 121);
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v704\(80 to 95) & X"000" & X"1")));
                      state_var3000 <= pause_getI2908;
                    when others =>
                      eclat_print_string(of_string("unknown primitive"));
                      
                      \$v704\ := "000"& X"000000" & X"1" & eclat_true & \$v522\(0 to 15) & \$v522\(16 to 47) & \$187_sp\ & \$v522\(64 to 95) & \$v522\(96 to 103) & \$v522\(104 to 119) & \$v522\(120 to 121);
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v704\(80 to 95) & X"000" & X"1")));
                      state_var3000 <= pause_getI2908;
                    end case;
                  when pause_setI2921 =>
                    \$ram_write_request\ <= '0';
                    \$210_sp\ := eclat_add(\$v718\(32 to 47) & X"000" & X"1");
                    \$v2920\ := argument1;
                    case \$v2920\ is
                    when "000"& X"000000" & X"0" =>
                      eclat_print_string(of_string("======> "));
                      
                      eclat_print_int(\$v522\(16 to 46));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$v719\ := "000"& X"000000" & X"1" & eclat_true & \$v522\(0 to 15) & \$v522\(16 to 47) & \$210_sp\ & \$v522\(64 to 95) & \$v522\(96 to 103) & \$v522\(104 to 119) & \$v522\(120 to 121);
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v719\(80 to 95) & X"000" & X"1")));
                      state_var3000 <= pause_getI2918;
                    when others =>
                      eclat_print_string(of_string("unknown primitive"));
                      
                      \$v719\ := "000"& X"000000" & X"1" & eclat_true & \$v522\(0 to 15) & \$v522\(16 to 47) & \$210_sp\ & \$v522\(64 to 95) & \$v522\(96 to 103) & \$v522\(104 to 119) & \$v522\(120 to 121);
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v719\(80 to 95) & X"000" & X"1")));
                      state_var3000 <= pause_getI2918;
                    end case;
                  when pause_setI2930 =>
                    \$ram_write_request\ <= '0';
                    \$351_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"2") & argument1 & eclat_true & \$351_sp\ & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_setI2931 =>
                    \$ram_write_request\ <= '0';
                    result2582 := eclat_add(\$v522\(0 to 15) & X"000" & X"2") & "000"& X"000000" & X"1" & eclat_true & \$v522\(48 to 63) & \$v522\(64 to 119) & \$v522\(120 to 121);
                    rdy2583 := eclat_true;
                    state_var3000 <= compute2584;
                  when pause_setI2934 =>
                    \$ram_write_request\ <= '0';
                    w_arg := eclat_add(w_arg(0 to 15) & X"000" & X"1") & w_arg(16 to 31) & w_arg(32 to 47) & w_arg(48 to 63);
                    state_var3000 <= w;
                  when pause_setI2940 =>
                    \$ram_write_request\ <= '0';
                    fill_arg := eclat_add(fill_arg(0 to 15) & X"000" & X"1") & \$v581\(32 to 47) & fill_arg(32 to 47) & fill_arg(48 to 79);
                    state_var3000 <= fill;
                  when pause_setI2944 =>
                    \$ram_write_request\ <= '0';
                    \$v576\ := \$v584\(0 to 31) & \$v584\(32 to 63) & \$v584\(64 to 95);
                    fill_arg := X"000" & X"1" & \$55_sp\ & eclat_resize(argument1,16) & \$v576\(64 to 95);
                    state_var3000 <= fill;
                  when pause_setI2945 =>
                    \$ram_write_request\ <= '0';
                    \$55_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    make_block_id := X"0" & X"47";
                    make_block_arg := \$55_sp\ & \$v522\(16 to 47) & \$v522\(64 to 95) & X"f7" & eclat_add(eclat_resize(argument1,16) & X"000" & X"1");
                    state_var3000 <= make_block;
                  when pause_setI2955 =>
                    \$ram_write_request\ <= '0';
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(X"3e80" & eclat_resize(argument1,16))));
                    state_var3000 <= pause_getI2953;
                  when pause_setI2956 =>
                    \$ram_write_request\ <= '0';
                    \$74_fill_arg\ := eclat_add(\$74_fill_arg\(0 to 15) & X"000" & X"1") & \$v599\(32 to 47) & \$74_fill_arg\(32 to 63) & \$74_fill_arg\(64 to 79);
                    state_var3000 <= \$74_fill\;
                  when pause_setI2960 =>
                    \$ram_write_request\ <= '0';
                    \$74_fill_arg\ := X"000" & X"1" & \$v522\(48 to 63) & \$v593\(64 to 95) & eclat_resize(argument1,16);
                    state_var3000 <= \$74_fill\;
                  when pause_setI2961 =>
                    \$ram_write_request\ <= '0';
                    w0_arg := eclat_add(w0_arg(0 to 15) & X"000" & X"1") & \$v563\(32 to 47) & w0_arg(32 to 47) & w0_arg(48 to 79) & w0_arg(80 to 95);
                    state_var3000 <= w0;
                  when pause_setI2965 =>
                    \$ram_write_request\ <= '0';
                    w1_arg := eclat_add(w1_arg(0 to 15) & X"000" & X"1") & w1_arg(16 to 31) & w1_arg(32 to 47) & w1_arg(48 to 79);
                    state_var3000 <= w1;
                  when pause_setI2968 =>
                    \$ram_write_request\ <= '0';
                    \$code_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(w1_arg(16 to 31) & X"000" & X"3") & w1_arg(0 to 15))));
                    state_var3000 <= pause_getI2966;
                  when pause_setI2970 =>
                    \$ram_write_request\ <= '0';
                    \$39_sp\ := eclat_add(w3_arg(16 to 31) & X"000" & X"1");
                    w3_arg := eclat_add(w3_arg(0 to 15) & X"000" & X"1") & \$39_sp\ & w3_arg(32 to 47) & w3_arg(48 to 79);
                    state_var3000 <= w3;
                  when pause_setI2972 =>
                    \$ram_write_request\ <= '0';
                    \$34_sp\ := eclat_add(\$33_sp\ & X"000" & X"1");
                    w3_arg := X"000" & X"1" & \$34_sp\ & eclat_resize(argument1,16) & \$v540\(64 to 95);
                    state_var3000 <= w3;
                  when pause_setI2973 =>
                    \$ram_write_request\ <= '0';
                    w0_arg := X"000" & X"0" & \$30_sp\ & eclat_resize(argument1,16) & \$v540\(64 to 95) & eclat_resize(argument2,16);
                    state_var3000 <= w0;
                  when pause_setI2974 =>
                    \$ram_write_request\ <= '0';
                    \$30_sp\ := eclat_add(\$v522\(48 to 63) & X"000" & X"1");
                    make_block_id := X"0" & X"53";
                    make_block_arg := \$30_sp\ & \$v522\(16 to 47) & \$v522\(64 to 95) & X"f7" & eclat_add(eclat_sub(eclat_mult(X"000" & X"2" & eclat_resize(argument1,16)) & X"000" & X"1") & eclat_resize(argument2,16));
                    state_var3000 <= make_block;
                  when w =>
                    \$v2937\ := eclat_gt(w_arg(0 to 15) & w_arg(32 to 47));
                    if \$v2937\(0) = '1' then
                      w_result := eclat_unit;
                      \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v522\(16 to 46),16) & X"000" & X"0") & X"000" & X"1")));
                      state_var3000 <= pause_getI2938;
                    else
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(w_arg(16 to 31) & w_arg(0 to 15))));
                      state_var3000 <= pause_getI2935;
                    end if;
                  when w0 =>
                    \$v2964\ := eclat_ge(w0_arg(0 to 15) & w0_arg(80 to 95));
                    if \$v2964\(0) = '1' then
                      w0_result := w0_arg(16 to 31);
                      \$33_sp\ := w0_result;
                      w1_arg := X"000" & X"1" & \$v522\(0 to 15) & eclat_resize(argument1,16) & \$v540\(64 to 95);
                      state_var3000 <= w1;
                    else
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(w0_arg(16 to 31) & X"000" & X"1")));
                      state_var3000 <= pause_getI2962;
                    end if;
                  when w1 =>
                    \$v2969\ := eclat_ge(w1_arg(0 to 15) & w1_arg(32 to 47));
                    if \$v2969\(0) = '1' then
                      w1_result := eclat_unit;
                      \$ram_ptr_write\ <= to_integer(unsigned(\$33_sp\));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v540\(64 to 95);
                      state_var3000 <= pause_setI2972;
                    else
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(w1_arg(48 to 78),16) & eclat_sub(eclat_mult(X"000" & X"2" & w1_arg(0 to 15)) & X"000" & X"1")) & X"000" & X"1")));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= eclat_lor(eclat_lsl(eclat_resize(X"f9",31) & "000"& X"00000" & X"18") & eclat_lsl(eclat_resize(eclat_mult(X"000" & X"2" & w1_arg(0 to 15)),31) & "000"& X"000000" & X"2")) & eclat_true;
                      state_var3000 <= pause_setI2968;
                    end if;
                  when w3 =>
                    \$v2971\ := eclat_ge(w3_arg(0 to 15) & w3_arg(32 to 47));
                    if \$v2971\(0) = '1' then
                      w3_result := w3_arg(16 to 31);
                      \$35_sp\ := w3_result;
                      result2582 := eclat_add(eclat_add(\$v522\(0 to 15) & X"000" & X"3") & eclat_resize(argument1,16)) & \$v540\(64 to 95) & \$35_sp\ & \$v540\(32 to 63) & \$v522\(96 to 103) & \$v522\(104 to 119) & \$v522\(120 to 121);
                      rdy2583 := eclat_true;
                      state_var3000 <= compute2584;
                    else
                      \$ram_ptr_write\ <= to_integer(unsigned(w3_arg(16 to 31)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= eclat_resize(eclat_add(eclat_resize(w3_arg(48 to 78),16) & eclat_mult(X"000" & X"2" & w3_arg(0 to 15))),31) & eclat_true;
                      state_var3000 <= pause_setI2970;
                    end if;
                  when \wait\ =>
                    \$v2659\ := eclat_not(\$v1397_init_done\);
                    if \$v2659\(0) = '1' then
                      \$v1397\ := wait_arg(1 to 32) & wait_arg(33 to 64) & X"0" & X"fa0" & X"0" & X"fa0" & X"0" & X"fa0" & eclat_add(X"0" & X"fa0" & X"1770") & eclat_false;
                      \$v1397_init_done\ := eclat_true;
                    end if;
                    case state_var3001 is
                    when \$1410_forever\ =>
                      state_var3001 <= \$1410_forever\;
                    when \$1452_loop\ =>
                      \$v2594\ := eclat_ge(\$1452_loop_arg\(0 to 15) & eclat_add(\$1452_loop_arg\(48 to 63) & X"000" & X"1"));
                      if \$v2594\(0) = '1' then
                        \$1452_loop_result\ := eclat_unit;
                        \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$v412\(0 to 30),16)));
                        \$ram_write_request\ <= '1';
                        \$ram_write\ <= eclat_resize(copy_root_in_ram_arg(32 to 47),31) & eclat_false;
                        state_var3001 <= pause_setI2596;
                      else
                        \$ram_ptr\ <= to_integer(unsigned(eclat_add(\$1452_loop_arg\(32 to 47) & \$1452_loop_arg\(0 to 15))));
                        state_var3001 <= pause_getI2592;
                      end if;
                    when \$1489_loop\ =>
                      \$v2633\ := eclat_ge(\$1489_loop_arg\(0 to 15) & eclat_add(\$1489_loop_arg\(48 to 63) & X"000" & X"1"));
                      if \$v2633\(0) = '1' then
                        \$1489_loop_result\ := eclat_unit;
                        \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(wait_arg(33 to 63),16)));
                        \$ram_write_request\ <= '1';
                        \$ram_write\ <= eclat_resize(\$v1408\(32 to 47),31) & eclat_false;
                        state_var3001 <= pause_setI2635;
                      else
                        \$ram_ptr\ <= to_integer(unsigned(eclat_add(\$1489_loop_arg\(32 to 47) & \$1489_loop_arg\(0 to 15))));
                        state_var3001 <= pause_getI2631;
                      end if;
                    when \$1526_loop\ =>
                      \$v2646\ := eclat_ge(\$1526_loop_arg\(0 to 15) & eclat_add(\$1526_loop_arg\(48 to 63) & X"000" & X"1"));
                      if \$v2646\(0) = '1' then
                        \$1526_loop_result\ := eclat_unit;
                        \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(wait_arg(1 to 31),16)));
                        \$ram_write_request\ <= '1';
                        \$ram_write\ <= eclat_resize(\$v1397\(112 to 127),31) & eclat_false;
                        state_var3001 <= pause_setI2648;
                      else
                        \$ram_ptr\ <= to_integer(unsigned(eclat_add(\$1526_loop_arg\(32 to 47) & \$1526_loop_arg\(0 to 15))));
                        state_var3001 <= pause_getI2644;
                      end if;
                    when \$581_loop\ =>
                      \$v2611\ := eclat_ge(\$581_loop_arg\(0 to 15) & eclat_add(\$581_loop_arg\(48 to 63) & X"000" & X"1"));
                      if \$v2611\(0) = '1' then
                        \$581_loop_result\ := eclat_unit;
                        \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$v400\(0 to 30),16)));
                        \$ram_write_request\ <= '1';
                        \$ram_write\ <= eclat_resize(loop_arg(16 to 31),31) & eclat_false;
                        state_var3001 <= pause_setI2613;
                      else
                        \$ram_ptr\ <= to_integer(unsigned(eclat_add(\$581_loop_arg\(32 to 47) & \$581_loop_arg\(0 to 15))));
                        state_var3001 <= pause_getI2609;
                      end if;
                    when aux =>
                      eclat_print_string(of_string("     scan="));
                      
                      eclat_print_int(aux_arg(0 to 15));
                      
                      eclat_print_string(of_string(" | next="));
                      
                      eclat_print_int(aux_arg(16 to 31));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$v2626\ := eclat_ge(aux_arg(0 to 15) & aux_arg(16 to 31));
                      if \$v2626\(0) = '1' then
                        aux_result := aux_arg(16 to 31);
                        \$558_next\ := aux_result;
                        eclat_print_string(of_string("memory copied in to_space : "));
                        
                        eclat_print_int(eclat_sub(\$558_next\ & \$v1397\(112 to 127)));
                        
                        eclat_print_string(of_string(" words"));
                        
                        eclat_print_newline(eclat_unit);
                        
                        \$v2627\ := eclat_gt(eclat_sub(\$558_next\ & \$v1397\(112 to 127)) & X"1770");
                        if \$v2627\(0) = '1' then
                          eclat_print_string(of_string("fatal error: "));
                          
                          eclat_print_string(of_string("Out of memory"));
                          
                          eclat_print_newline(eclat_unit);
                          
                          state_var3001 <= \$1410_forever\;
                        else
                          \$v1400\ := \$v1408\(0 to 31) & \$v1409\(0 to 31) & \$558_next\;
                          eclat_print_newline(eclat_unit);
                          
                          eclat_print_newline(eclat_unit);
                          
                          eclat_print_string(of_string("[================= GC END ======================]"));
                          
                          eclat_print_newline(eclat_unit);
                          
                          eclat_print_newline(eclat_unit);
                          
                          result2587 := \$v1400\(0 to 31) & \$v1400\(32 to 63) & \$v1400\(64 to 79) & eclat_add(\$v1400\(64 to 79) & wait_arg(81 to 96)) & \$v1397\(112 to 127) & \$v1397\(96 to 111);
                          rdy2588 := eclat_true;
                          state_var3001 <= compute2589;
                        end if;
                      else
                        \$ram_ptr\ <= to_integer(unsigned(aux_arg(0 to 15)));
                        state_var3001 <= pause_getI2624;
                      end if;
                    when copy_root_in_ram =>
                      \$v2606\ := eclat_ge(copy_root_in_ram_arg(0 to 15) & copy_root_in_ram_arg(16 to 31));
                      if \$v2606\(0) = '1' then
                        copy_root_in_ram_result := copy_root_in_ram_arg(32 to 47);
                        case copy_root_in_ram_id is
                        when X"00" & X"6" =>
                          \$557_next\ := copy_root_in_ram_result;
                          eclat_print_string(of_string("======================================="));
                          
                          eclat_print_newline(eclat_unit);
                          
                          aux_arg := \$v1397\(112 to 127) & \$557_next\ & \$v1397\(96 to 111) & \$v1397\(112 to 127);
                          state_var3001 <= aux;
                        when X"00" & X"7" =>
                          \$556_next\ := copy_root_in_ram_result;
                          \$global_end_ptr\ <= 0;
                          state_var3001 <= pause_getI2628;
                        when others =>
                          
                        end case;
                      else
                        eclat_print_string(of_string("racine:"));
                        
                        eclat_print_int(copy_root_in_ram_arg(0 to 15));
                        
                        eclat_print_newline(eclat_unit);
                        
                        \$ram_ptr\ <= to_integer(unsigned(copy_root_in_ram_arg(0 to 15)));
                        state_var3001 <= pause_getI2604;
                      end if;
                    when \loop\ =>
                      \$v2623\ := eclat_ge(loop_arg(0 to 15) & eclat_add(loop_arg(64 to 79) & X"000" & X"1"));
                      if \$v2623\(0) = '1' then
                        loop_result := loop_arg(16 to 31);
                        \$562_next\ := loop_result;
                        aux_arg := eclat_add(aux_arg(0 to 15) & eclat_add(eclat_resize(eclat_lsr(eclat_resize(eclat_resize(\$v402\(0 to 30),16),31) & "000"& X"000000" & X"2"),16) & X"000" & X"1")) & \$562_next\ & aux_arg(32 to 47) & aux_arg(48 to 63);
                        state_var3001 <= aux;
                      else
                        \$ram_ptr\ <= to_integer(unsigned(eclat_add(loop_arg(80 to 95) & loop_arg(0 to 15))));
                        state_var3001 <= pause_getI2621;
                      end if;
                    when pause_getI2592 =>
                      state_var3001 <= pause_getII2593;
                    when pause_getI2598 =>
                      state_var3001 <= pause_getII2599;
                    when pause_getI2601 =>
                      state_var3001 <= pause_getII2602;
                    when pause_getI2604 =>
                      state_var3001 <= pause_getII2605;
                    when pause_getI2609 =>
                      state_var3001 <= pause_getII2610;
                    when pause_getI2615 =>
                      state_var3001 <= pause_getII2616;
                    when pause_getI2618 =>
                      state_var3001 <= pause_getII2619;
                    when pause_getI2621 =>
                      state_var3001 <= pause_getII2622;
                    when pause_getI2624 =>
                      state_var3001 <= pause_getII2625;
                    when pause_getI2628 =>
                      state_var3001 <= pause_getII2629;
                    when pause_getI2631 =>
                      state_var3001 <= pause_getII2632;
                    when pause_getI2637 =>
                      state_var3001 <= pause_getII2638;
                    when pause_getI2640 =>
                      state_var3001 <= pause_getII2641;
                    when pause_getI2644 =>
                      state_var3001 <= pause_getII2645;
                    when pause_getI2650 =>
                      state_var3001 <= pause_getII2651;
                    when pause_getI2653 =>
                      state_var3001 <= pause_getII2654;
                    when pause_getII2593 =>
                      \$1464\ := \$ram_value\;
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(\$1452_loop_arg\(16 to 31) & \$1452_loop_arg\(0 to 15))));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$1464\;
                      state_var3001 <= pause_setI2591;
                    when pause_getII2599 =>
                      \$1449_hd\ := \$ram_value\;
                      eclat_print_string(of_string("bloc "));
                      
                      eclat_print_int(eclat_resize(\$v412\(0 to 30),16));
                      
                      eclat_print_string(of_string(" of size "));
                      
                      eclat_print_int(eclat_add(eclat_resize(eclat_lsr(\$1449_hd\(0 to 30) & "000"& X"000000" & X"2"),16) & X"000" & X"1"));
                      
                      eclat_print_string(of_string(" from "));
                      
                      eclat_print_int(eclat_resize(\$v412\(0 to 30),16));
                      
                      eclat_print_string(of_string(" to "));
                      
                      eclat_print_int(copy_root_in_ram_arg(32 to 47));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$ram_ptr_write\ <= to_integer(unsigned(copy_root_in_ram_arg(32 to 47)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$1449_hd\;
                      state_var3001 <= pause_setI2597;
                    when pause_getII2602 =>
                      \$1447_w\ := \$ram_value\;
                      \$v2600\ := eclat_if(eclat_not(""&\$1447_w\(31)) & 
                                  eclat_if(eclat_le(copy_root_in_ram_arg(64 to 79) & eclat_resize(\$1447_w\(0 to 30),16)) & eclat_lt(eclat_resize(\$1447_w\(0 to 30),16) & eclat_add(copy_root_in_ram_arg(64 to 79) & X"1770")) & eclat_false) & eclat_false);
                      if \$v2600\(0) = '1' then
                        \$v1468\ := \$1447_w\ & copy_root_in_ram_arg(32 to 47);
                        \$ram_ptr_write\ <= to_integer(unsigned(copy_root_in_ram_arg(0 to 15)));
                        \$ram_write_request\ <= '1';
                        \$ram_write\ <= \$v1468\(0 to 31);
                        state_var3001 <= pause_setI2590;
                      else
                        \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$v412\(0 to 30),16)));
                        state_var3001 <= pause_getI2598;
                      end if;
                    when pause_getII2605 =>
                      \$v412\ := \$ram_value\;
                      \$v2603\ := eclat_not(eclat_if(eclat_not(""&\$v412\(31)) & 
                                            eclat_if(eclat_le(copy_root_in_ram_arg(48 to 63) & eclat_resize(\$v412\(0 to 30),16)) & eclat_lt(eclat_resize(\$v412\(0 to 30),16) & eclat_add(copy_root_in_ram_arg(48 to 63) & X"1770")) & eclat_false) & eclat_false));
                      if \$v2603\(0) = '1' then
                        \$v1468\ := \$v412\ & copy_root_in_ram_arg(32 to 47);
                        \$ram_ptr_write\ <= to_integer(unsigned(copy_root_in_ram_arg(0 to 15)));
                        \$ram_write_request\ <= '1';
                        \$ram_write\ <= \$v1468\(0 to 31);
                        state_var3001 <= pause_setI2590;
                      else
                        \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_resize(\$v412\(0 to 30),16) & X"000" & X"1")));
                        state_var3001 <= pause_getI2601;
                      end if;
                    when pause_getII2610 =>
                      \$v426\ := \$ram_value\;
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(\$581_loop_arg\(16 to 31) & \$581_loop_arg\(0 to 15))));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v426\;
                      state_var3001 <= pause_setI2608;
                    when pause_getII2616 =>
                      \$579_hd\ := \$ram_value\;
                      eclat_print_string(of_string("bloc "));
                      
                      eclat_print_int(eclat_resize(\$v400\(0 to 30),16));
                      
                      eclat_print_string(of_string(" of size "));
                      
                      eclat_print_int(eclat_add(eclat_resize(eclat_lsr(\$579_hd\(0 to 30) & "000"& X"000000" & X"2"),16) & X"000" & X"1"));
                      
                      eclat_print_string(of_string(" from "));
                      
                      eclat_print_int(eclat_resize(\$v400\(0 to 30),16));
                      
                      eclat_print_string(of_string(" to "));
                      
                      eclat_print_int(loop_arg(16 to 31));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$ram_ptr_write\ <= to_integer(unsigned(loop_arg(16 to 31)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$579_hd\;
                      state_var3001 <= pause_setI2614;
                    when pause_getII2619 =>
                      \$578_w\ := \$ram_value\;
                      \$v2617\ := eclat_if(eclat_not(""&\$578_w\(31)) & 
                                  eclat_if(eclat_le(loop_arg(48 to 63) & eclat_resize(\$578_w\(0 to 30),16)) & eclat_lt(eclat_resize(\$578_w\(0 to 30),16) & eclat_add(loop_arg(48 to 63) & X"1770")) & eclat_false) & eclat_false);
                      if \$v2617\(0) = '1' then
                        \$v1433\ := \$578_w\ & loop_arg(16 to 31);
                        \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(loop_arg(80 to 95) & loop_arg(0 to 15))));
                        \$ram_write_request\ <= '1';
                        \$ram_write\ <= \$v1433\(0 to 31);
                        state_var3001 <= pause_setI2607;
                      else
                        \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$v400\(0 to 30),16)));
                        state_var3001 <= pause_getI2615;
                      end if;
                    when pause_getII2622 =>
                      \$v400\ := \$ram_value\;
                      \$v2620\ := eclat_not(eclat_if(eclat_not(""&\$v400\(31)) & 
                                            eclat_if(eclat_le(loop_arg(32 to 47) & eclat_resize(\$v400\(0 to 30),16)) & eclat_lt(eclat_resize(\$v400\(0 to 30),16) & eclat_add(loop_arg(32 to 47) & X"1770")) & eclat_false) & eclat_false));
                      if \$v2620\(0) = '1' then
                        \$v1433\ := \$v400\ & loop_arg(16 to 31);
                        \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(loop_arg(80 to 95) & loop_arg(0 to 15))));
                        \$ram_write_request\ <= '1';
                        \$ram_write\ <= \$v1433\(0 to 31);
                        state_var3001 <= pause_setI2607;
                      else
                        \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_resize(\$v400\(0 to 30),16) & X"000" & X"1")));
                        state_var3001 <= pause_getI2618;
                      end if;
                    when pause_getII2625 =>
                      \$v402\ := \$ram_value\;
                      loop_arg := X"000" & X"1" & aux_arg(16 to 31) & aux_arg(32 to 47) & aux_arg(48 to 63) & eclat_resize(eclat_lsr(eclat_resize(eclat_resize(\$v402\(0 to 30),16),31) & "000"& X"000000" & X"2"),16) & aux_arg(0 to 15);
                      state_var3001 <= \loop\;
                    when pause_getII2629 =>
                      \$v407\ := \$global_end_value\;
                      copy_root_in_ram_id := X"00" & X"6";
                      copy_root_in_ram_arg := X"3e80" & \$v407\ & \$556_next\ & \$v1397\(96 to 111) & \$v1397\(112 to 127);
                      state_var3001 <= copy_root_in_ram;
                    when pause_getII2632 =>
                      \$1501\ := \$ram_value\;
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(\$1489_loop_arg\(16 to 31) & \$1489_loop_arg\(0 to 15))));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$1501\;
                      state_var3001 <= pause_setI2630;
                    when pause_getII2638 =>
                      \$1486_hd\ := \$ram_value\;
                      eclat_print_string(of_string("bloc "));
                      
                      eclat_print_int(eclat_resize(wait_arg(33 to 63),16));
                      
                      eclat_print_string(of_string(" of size "));
                      
                      eclat_print_int(eclat_add(eclat_resize(eclat_lsr(\$1486_hd\(0 to 30) & "000"& X"000000" & X"2"),16) & X"000" & X"1"));
                      
                      eclat_print_string(of_string(" from "));
                      
                      eclat_print_int(eclat_resize(wait_arg(33 to 63),16));
                      
                      eclat_print_string(of_string(" to "));
                      
                      eclat_print_int(\$v1408\(32 to 47));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v1408\(32 to 47)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$1486_hd\;
                      state_var3001 <= pause_setI2636;
                    when pause_getII2641 =>
                      \$1484_w\ := \$ram_value\;
                      \$v2639\ := eclat_if(eclat_not(""&\$1484_w\(31)) & 
                                  eclat_if(eclat_le(\$v1397\(112 to 127) & eclat_resize(\$1484_w\(0 to 30),16)) & eclat_lt(eclat_resize(\$1484_w\(0 to 30),16) & eclat_add(\$v1397\(112 to 127) & X"1770")) & eclat_false) & eclat_false);
                      if \$v2639\(0) = '1' then
                        \$v1409\ := \$1484_w\ & \$v1408\(32 to 47);
                        copy_root_in_ram_id := X"00" & X"7";
                        copy_root_in_ram_arg := X"0" & X"3e8" & wait_arg(65 to 80) & \$v1409\(32 to 47) & \$v1397\(96 to 111) & \$v1397\(112 to 127);
                        state_var3001 <= copy_root_in_ram;
                      else
                        \$ram_ptr\ <= to_integer(unsigned(eclat_resize(wait_arg(33 to 63),16)));
                        state_var3001 <= pause_getI2637;
                      end if;
                    when pause_getII2645 =>
                      \$1538\ := \$ram_value\;
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(\$1526_loop_arg\(16 to 31) & \$1526_loop_arg\(0 to 15))));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$1538\;
                      state_var3001 <= pause_setI2643;
                    when pause_getII2651 =>
                      \$1523_hd\ := \$ram_value\;
                      eclat_print_string(of_string("bloc "));
                      
                      eclat_print_int(eclat_resize(wait_arg(1 to 31),16));
                      
                      eclat_print_string(of_string(" of size "));
                      
                      eclat_print_int(eclat_add(eclat_resize(eclat_lsr(\$1523_hd\(0 to 30) & "000"& X"000000" & X"2"),16) & X"000" & X"1"));
                      
                      eclat_print_string(of_string(" from "));
                      
                      eclat_print_int(eclat_resize(wait_arg(1 to 31),16));
                      
                      eclat_print_string(of_string(" to "));
                      
                      eclat_print_int(\$v1397\(112 to 127));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v1397\(112 to 127)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$1523_hd\;
                      state_var3001 <= pause_setI2649;
                    when pause_getII2654 =>
                      \$1521_w\ := \$ram_value\;
                      \$v2652\ := eclat_if(eclat_not(""&\$1521_w\(31)) & 
                                  eclat_if(eclat_le(\$v1397\(112 to 127) & eclat_resize(\$1521_w\(0 to 30),16)) & eclat_lt(eclat_resize(\$1521_w\(0 to 30),16) & eclat_add(\$v1397\(112 to 127) & X"1770")) & eclat_false) & eclat_false);
                      if \$v2652\(0) = '1' then
                        \$v1408\ := \$1521_w\ & \$v1397\(112 to 127);
                        \$v2642\ := eclat_not(eclat_if(eclat_not(""&wait_arg(64)) & 
                                              eclat_if(eclat_le(\$v1397\(96 to 111) & eclat_resize(wait_arg(33 to 63),16)) & eclat_lt(eclat_resize(wait_arg(33 to 63),16) & eclat_add(\$v1397\(96 to 111) & X"1770")) & eclat_false) & eclat_false));
                        if \$v2642\(0) = '1' then
                          \$v1409\ := wait_arg(33 to 64) & \$v1408\(32 to 47);
                          copy_root_in_ram_id := X"00" & X"7";
                          copy_root_in_ram_arg := X"0" & X"3e8" & wait_arg(65 to 80) & \$v1409\(32 to 47) & \$v1397\(96 to 111) & \$v1397\(112 to 127);
                          state_var3001 <= copy_root_in_ram;
                        else
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_resize(wait_arg(33 to 63),16) & X"000" & X"1")));
                          state_var3001 <= pause_getI2640;
                        end if;
                      else
                        \$ram_ptr\ <= to_integer(unsigned(eclat_resize(wait_arg(1 to 31),16)));
                        state_var3001 <= pause_getI2650;
                      end if;
                    when pause_setI2590 =>
                      \$ram_write_request\ <= '0';
                      eclat_print_string(of_string(" next="));
                      
                      eclat_print_int(\$v1468\(32 to 47));
                      
                      eclat_print_newline(eclat_unit);
                      
                      copy_root_in_ram_arg := eclat_add(copy_root_in_ram_arg(0 to 15) & X"000" & X"1") & copy_root_in_ram_arg(16 to 31) & \$v1468\(32 to 47) & copy_root_in_ram_arg(48 to 63) & copy_root_in_ram_arg(64 to 79);
                      state_var3001 <= copy_root_in_ram;
                    when pause_setI2591 =>
                      \$ram_write_request\ <= '0';
                      \$1452_loop_arg\ := eclat_add(\$1452_loop_arg\(0 to 15) & X"000" & X"1") & \$1452_loop_arg\(16 to 31) & \$1452_loop_arg\(32 to 47) & \$1452_loop_arg\(48 to 63);
                      state_var3001 <= \$1452_loop\;
                    when pause_setI2595 =>
                      \$ram_write_request\ <= '0';
                      \$v1468\ := eclat_resize(copy_root_in_ram_arg(32 to 47),31) & eclat_false & eclat_add(copy_root_in_ram_arg(32 to 47) & eclat_add(eclat_resize(eclat_lsr(\$1449_hd\(0 to 30) & "000"& X"000000" & X"2"),16) & X"000" & X"1"));
                      \$ram_ptr_write\ <= to_integer(unsigned(copy_root_in_ram_arg(0 to 15)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v1468\(0 to 31);
                      state_var3001 <= pause_setI2590;
                    when pause_setI2596 =>
                      \$ram_write_request\ <= '0';
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_resize(\$v412\(0 to 30),16) & X"000" & X"1")));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= eclat_resize(copy_root_in_ram_arg(32 to 47),31) & eclat_false;
                      state_var3001 <= pause_setI2595;
                    when pause_setI2597 =>
                      \$ram_write_request\ <= '0';
                      \$1452_loop_arg\ := X"000" & X"1" & copy_root_in_ram_arg(32 to 47) & eclat_resize(\$v412\(0 to 30),16) & eclat_resize(eclat_lsr(\$1449_hd\(0 to 30) & "000"& X"000000" & X"2"),16);
                      state_var3001 <= \$1452_loop\;
                    when pause_setI2607 =>
                      \$ram_write_request\ <= '0';
                      loop_arg := eclat_add(loop_arg(0 to 15) & X"000" & X"1") & \$v1433\(32 to 47) & loop_arg(32 to 47) & loop_arg(48 to 63) & loop_arg(64 to 79) & loop_arg(80 to 95);
                      state_var3001 <= \loop\;
                    when pause_setI2608 =>
                      \$ram_write_request\ <= '0';
                      \$581_loop_arg\ := eclat_add(\$581_loop_arg\(0 to 15) & X"000" & X"1") & \$581_loop_arg\(16 to 31) & \$581_loop_arg\(32 to 47) & \$581_loop_arg\(48 to 63);
                      state_var3001 <= \$581_loop\;
                    when pause_setI2612 =>
                      \$ram_write_request\ <= '0';
                      \$v1433\ := eclat_resize(loop_arg(16 to 31),31) & eclat_false & eclat_add(loop_arg(16 to 31) & eclat_add(eclat_resize(eclat_lsr(\$579_hd\(0 to 30) & "000"& X"000000" & X"2"),16) & X"000" & X"1"));
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(loop_arg(80 to 95) & loop_arg(0 to 15))));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v1433\(0 to 31);
                      state_var3001 <= pause_setI2607;
                    when pause_setI2613 =>
                      \$ram_write_request\ <= '0';
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_resize(\$v400\(0 to 30),16) & X"000" & X"1")));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= eclat_resize(loop_arg(16 to 31),31) & eclat_false;
                      state_var3001 <= pause_setI2612;
                    when pause_setI2614 =>
                      \$ram_write_request\ <= '0';
                      \$581_loop_arg\ := X"000" & X"1" & loop_arg(16 to 31) & eclat_resize(\$v400\(0 to 30),16) & eclat_resize(eclat_lsr(\$579_hd\(0 to 30) & "000"& X"000000" & X"2"),16);
                      state_var3001 <= \$581_loop\;
                    when pause_setI2630 =>
                      \$ram_write_request\ <= '0';
                      \$1489_loop_arg\ := eclat_add(\$1489_loop_arg\(0 to 15) & X"000" & X"1") & \$1489_loop_arg\(16 to 31) & \$1489_loop_arg\(32 to 47) & \$1489_loop_arg\(48 to 63);
                      state_var3001 <= \$1489_loop\;
                    when pause_setI2634 =>
                      \$ram_write_request\ <= '0';
                      \$v1409\ := eclat_resize(\$v1408\(32 to 47),31) & eclat_false & eclat_add(\$v1408\(32 to 47) & eclat_add(eclat_resize(eclat_lsr(\$1486_hd\(0 to 30) & "000"& X"000000" & X"2"),16) & X"000" & X"1"));
                      copy_root_in_ram_id := X"00" & X"7";
                      copy_root_in_ram_arg := X"0" & X"3e8" & wait_arg(65 to 80) & \$v1409\(32 to 47) & \$v1397\(96 to 111) & \$v1397\(112 to 127);
                      state_var3001 <= copy_root_in_ram;
                    when pause_setI2635 =>
                      \$ram_write_request\ <= '0';
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_resize(wait_arg(33 to 63),16) & X"000" & X"1")));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= eclat_resize(\$v1408\(32 to 47),31) & eclat_false;
                      state_var3001 <= pause_setI2634;
                    when pause_setI2636 =>
                      \$ram_write_request\ <= '0';
                      \$1489_loop_arg\ := X"000" & X"1" & \$v1408\(32 to 47) & eclat_resize(wait_arg(33 to 63),16) & eclat_resize(eclat_lsr(\$1486_hd\(0 to 30) & "000"& X"000000" & X"2"),16);
                      state_var3001 <= \$1489_loop\;
                    when pause_setI2643 =>
                      \$ram_write_request\ <= '0';
                      \$1526_loop_arg\ := eclat_add(\$1526_loop_arg\(0 to 15) & X"000" & X"1") & \$1526_loop_arg\(16 to 31) & \$1526_loop_arg\(32 to 47) & \$1526_loop_arg\(48 to 63);
                      state_var3001 <= \$1526_loop\;
                    when pause_setI2647 =>
                      \$ram_write_request\ <= '0';
                      \$v1408\ := eclat_resize(\$v1397\(112 to 127),31) & eclat_false & eclat_add(\$v1397\(112 to 127) & eclat_add(eclat_resize(eclat_lsr(\$1523_hd\(0 to 30) & "000"& X"000000" & X"2"),16) & X"000" & X"1"));
                      \$v2642\ := eclat_not(eclat_if(eclat_not(""&wait_arg(64)) & 
                                            eclat_if(eclat_le(\$v1397\(96 to 111) & eclat_resize(wait_arg(33 to 63),16)) & eclat_lt(eclat_resize(wait_arg(33 to 63),16) & eclat_add(\$v1397\(96 to 111) & X"1770")) & eclat_false) & eclat_false));
                      if \$v2642\(0) = '1' then
                        \$v1409\ := wait_arg(33 to 64) & \$v1408\(32 to 47);
                        copy_root_in_ram_id := X"00" & X"7";
                        copy_root_in_ram_arg := X"0" & X"3e8" & wait_arg(65 to 80) & \$v1409\(32 to 47) & \$v1397\(96 to 111) & \$v1397\(112 to 127);
                        state_var3001 <= copy_root_in_ram;
                      else
                        \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_resize(wait_arg(33 to 63),16) & X"000" & X"1")));
                        state_var3001 <= pause_getI2640;
                      end if;
                    when pause_setI2648 =>
                      \$ram_write_request\ <= '0';
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_resize(wait_arg(1 to 31),16) & X"000" & X"1")));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= eclat_resize(\$v1397\(112 to 127),31) & eclat_false;
                      state_var3001 <= pause_setI2647;
                    when pause_setI2649 =>
                      \$ram_write_request\ <= '0';
                      \$1526_loop_arg\ := X"000" & X"1" & \$v1397\(112 to 127) & eclat_resize(wait_arg(1 to 31),16) & eclat_resize(eclat_lsr(\$1523_hd\(0 to 30) & "000"& X"000000" & X"2"),16);
                      state_var3001 <= \$1526_loop\;
                    when compute2589 =>
                      rdy2588 := eclat_false;
                      \$v2656\ := eclat_gt(eclat_add(\$v1397\(80 to 95) & wait_arg(81 to 96)) & eclat_add(\$v1397\(96 to 111) & X"1770"));
                      if \$v2656\(0) = '1' then
                        eclat_print_newline(eclat_unit);
                        
                        eclat_print_newline(eclat_unit);
                        
                        eclat_print_string(of_string("[================= GC START ======================]"));
                        
                        eclat_print_newline(eclat_unit);
                        
                        eclat_print_newline(eclat_unit);
                        
                        \$v2655\ := eclat_not(eclat_if(eclat_not(""&wait_arg(32)) & 
                                              eclat_if(eclat_le(\$v1397\(96 to 111) & eclat_resize(wait_arg(1 to 31),16)) & eclat_lt(eclat_resize(wait_arg(1 to 31),16) & eclat_add(\$v1397\(96 to 111) & X"1770")) & eclat_false) & eclat_false));
                        if \$v2655\(0) = '1' then
                          \$v1408\ := wait_arg(1 to 32) & \$v1397\(112 to 127);
                          \$v2642\ := eclat_not(eclat_if(eclat_not(""&wait_arg(64)) & 
                                                eclat_if(eclat_le(\$v1397\(96 to 111) & eclat_resize(wait_arg(33 to 63),16)) & eclat_lt(eclat_resize(wait_arg(33 to 63),16) & eclat_add(\$v1397\(96 to 111) & X"1770")) & eclat_false) & eclat_false));
                          if \$v2642\(0) = '1' then
                            \$v1409\ := wait_arg(33 to 64) & \$v1408\(32 to 47);
                            copy_root_in_ram_id := X"00" & X"7";
                            copy_root_in_ram_arg := X"0" & X"3e8" & wait_arg(65 to 80) & \$v1409\(32 to 47) & \$v1397\(96 to 111) & \$v1397\(112 to 127);
                            state_var3001 <= copy_root_in_ram;
                          else
                            \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_resize(wait_arg(33 to 63),16) & X"000" & X"1")));
                            state_var3001 <= pause_getI2640;
                          end if;
                        else
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_resize(wait_arg(1 to 31),16) & X"000" & X"1")));
                          state_var3001 <= pause_getI2653;
                        end if;
                      else
                        result2587 := wait_arg(1 to 32) & wait_arg(33 to 64) & \$v1397\(80 to 95) & eclat_add(\$v1397\(80 to 95) & wait_arg(81 to 96)) & \$v1397\(96 to 111) & \$v1397\(112 to 127);
                        rdy2588 := eclat_true;
                        state_var3001 <= compute2589;
                      end if;
                    end case;
                    \$v2658\ := eclat_not(rdy2588);
                    if \$v2658\(0) = '1' then
                      result2587 := \$v1397\(0 to 31) & \$v1397\(32 to 63) & \$v1397\(64 to 79) & \$v1397\(80 to 95) & \$v1397\(96 to 111) & \$v1397\(112 to 127);
                    end if;
                    \$v1397\ := result2587 & rdy2588;
                    \$v1395\ := \$v1397\;
                    \$v2586\ := ""&\$v1395\(128);
                    if \$v2586\(0) = '1' then
                      wait_result := \$v1395\(0 to 31) & \$v1395\(32 to 63) & \$v1395\(64 to 79);
                      \$v1380\ := wait_result;
                      eclat_print_string(of_string("size:"));
                      
                      eclat_print_int(eclat_if(eclat_eq(make_block_arg(88 to 103) & X"000" & X"0") & X"000" & X"1" & make_block_arg(88 to 103)));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v1380\(64 to 79)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= eclat_lor(eclat_lsl(eclat_resize(make_block_arg(80 to 87),31) & "000"& X"00000" & X"18") & eclat_lsl(eclat_resize(
                      eclat_if(eclat_eq(make_block_arg(88 to 103) & X"000" & X"0") & X"000" & X"1" & make_block_arg(88 to 103)),31) & "000"& X"000000" & X"2")) & eclat_true;
                      state_var3000 <= pause_setI2585;
                    else
                      wait_arg := eclat_unit & wait_arg(1 to 32) & wait_arg(33 to 64) & wait_arg(65 to 80) & wait_arg(81 to 96);
                      state_var3000 <= \wait\;
                    end if;
                  when compute2584 =>
                    rdy2583 := eclat_false;
                    eclat_print_string(of_string("pc:"));
                    
                    eclat_print_int(\$v522\(0 to 15));
                    
                    eclat_print_string(of_string("|acc:"));
                    
                    eclat_print_int(\$v522\(16 to 46));
                    
                    eclat_print_string(of_string("<"));
                    
                    \$v2991\ := ""&\$v522\(47);
                    if \$v2991\(0) = '1' then
                      eclat_print_string(of_string("int"));
                      
                      eclat_print_string(of_string(">"));
                      
                      eclat_print_string(of_string("|sp:"));
                      
                      eclat_print_int(\$v522\(48 to 63));
                      
                      eclat_print_string(of_string("|env:"));
                      
                      eclat_print_int(\$v522\(64 to 94));
                      
                      eclat_print_string(of_string("<"));
                      
                      \$v2990\ := ""&\$v522\(95);
                      if \$v2990\(0) = '1' then
                        eclat_print_string(of_string("int"));
                        
                        eclat_print_string(of_string(">"));
                        
                        eclat_print_newline(eclat_unit);
                        
                        assert eclat_lt(\$v522\(0 to 15) & std_logic_vector(to_unsigned(code'length,16))) = eclat_true report "assertion failed" severity error;
                        
                        \$code_ptr\ <= to_integer(unsigned(\$v522\(0 to 15)));
                        state_var3000 <= pause_getI2988;
                      else
                        eclat_print_string(of_string("ptr"));
                        
                        eclat_print_string(of_string(">"));
                        
                        eclat_print_newline(eclat_unit);
                        
                        assert eclat_lt(\$v522\(0 to 15) & std_logic_vector(to_unsigned(code'length,16))) = eclat_true report "assertion failed" severity error;
                        
                        \$code_ptr\ <= to_integer(unsigned(\$v522\(0 to 15)));
                        state_var3000 <= pause_getI2988;
                      end if;
                    else
                      eclat_print_string(of_string("ptr"));
                      
                      eclat_print_string(of_string(">"));
                      
                      eclat_print_string(of_string("|sp:"));
                      
                      eclat_print_int(\$v522\(48 to 63));
                      
                      eclat_print_string(of_string("|env:"));
                      
                      eclat_print_int(\$v522\(64 to 94));
                      
                      eclat_print_string(of_string("<"));
                      
                      \$v2990\ := ""&\$v522\(95);
                      if \$v2990\(0) = '1' then
                        eclat_print_string(of_string("int"));
                        
                        eclat_print_string(of_string(">"));
                        
                        eclat_print_newline(eclat_unit);
                        
                        assert eclat_lt(\$v522\(0 to 15) & std_logic_vector(to_unsigned(code'length,16))) = eclat_true report "assertion failed" severity error;
                        
                        \$code_ptr\ <= to_integer(unsigned(\$v522\(0 to 15)));
                        state_var3000 <= pause_getI2988;
                      else
                        eclat_print_string(of_string("ptr"));
                        
                        eclat_print_string(of_string(">"));
                        
                        eclat_print_newline(eclat_unit);
                        
                        assert eclat_lt(\$v522\(0 to 15) & std_logic_vector(to_unsigned(code'length,16))) = eclat_true report "assertion failed" severity error;
                        
                        \$code_ptr\ <= to_integer(unsigned(\$v522\(0 to 15)));
                        state_var3000 <= pause_getI2988;
                      end if;
                    end if;
                  end case;
                  \$v2993\ := eclat_not(rdy2583);
                  if \$v2993\(0) = '1' then
                    result2582 := \$v522\(0 to 121);
                  end if;
                  \$v524\ := result2582 & rdy2583;
                  \$v522\ := \$v524\(0 to 121) & ""&\$v524\(122);
                end if;
                \$v518\ := \$v522\;
                \$v516\ := ""&\$v518\(120) & ""&\$v518\(122) & ""&\$v516\(2) & ""&\$v518\(121);
              end if;
              \$v515\ := \$v516\;
              \$v509\ := ""&\$v515\(0) & eclat_not(""&\$v515\(1)) & ""&\$v515\(3);
              \$v2136\ := ""&\$v509\(0);
              if \$v2136\(0) = '1' then
                eclat_print_string(of_string("(cy="));
                
                eclat_print_int(cy);
                
                eclat_print_string(of_string(")"));
                
                eclat_print_newline(eclat_unit);
                
                \$v2135\ := eclat_not(\$v511_init_done\);
                if \$v2135\(0) = '1' then
                  \$v511\ := X"0000000" & X"0";
                  \$v511_init_done\ := eclat_true;
                end if;
                \$v511\ := eclat_if(eclat_eq(\$v511\ & eclat_add(X"00" & X"989680" & X"00" & X"989680")) & X"0000000" & X"0" & eclat_add(\$v511\ & X"0000000" & X"1"));
                \$v18\ := \$v511\;
                b := eclat_gt(\$v18\ & X"00" & X"989680");
                result2132 := ""&\$v509\(0) & ""&\$v509\(1) & b & ""&\$v509\(2) & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & X"0" & X"3" & X"0" & X"3" & X"0" & X"3" & X"0" & X"3" & X"0" & X"3" & X"0" & X"3";
                rdy2133 := eclat_true;
                state <= compute2134;
              else
                \$v2135\ := eclat_not(\$v511_init_done\);
                if \$v2135\(0) = '1' then
                  \$v511\ := X"0000000" & X"0";
                  \$v511_init_done\ := eclat_true;
                end if;
                \$v511\ := eclat_if(eclat_eq(\$v511\ & eclat_add(X"00" & X"989680" & X"00" & X"989680")) & X"0000000" & X"0" & eclat_add(\$v511\ & X"0000000" & X"1"));
                \$v18\ := \$v511\;
                b := eclat_gt(\$v18\ & X"00" & X"989680");
                result2132 := ""&\$v509\(0) & ""&\$v509\(1) & b & ""&\$v509\(2) & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & X"0" & X"3" & X"0" & X"3" & X"0" & X"3" & X"0" & X"3" & X"0" & X"3" & X"0" & X"3";
                rdy2133 := eclat_true;
                state <= compute2134;
              end if;
            end if;
          end case;
          
          result <= result2132;
          rdy <= rdy2133;
          
        end if;
      end if;
    end if;
  end process;
end architecture;
