-- code generated from the following source code:
--   stdlib.ecl
--   ../ocaml-vm/vm/mlvalue.ecl
--   ../ocaml-vm/vm/fail.ecl
--   ../ocaml-vm/vm/ram.ecl
--   ../ocaml-vm/vm/runtime.ecl
--   ../ocaml-vm/vm/debug.ecl
--   ../ocaml-vm/vm/alloc.ecl
--   ../ocaml-vm/vm/prims.ecl
--   ../ocaml-vm/bytecode.ecl
--   ../ocaml-vm/vm/vm.ecl
--   ../ocaml-vm/vm/target-specific/intel-max10/IOs.ecl
--   ../ocaml-vm/vm/target-specific/intel-max10/main.ecl
--
-- with the following command:
--
--    ./eclat -arg ((true,true,true,true,true,true,true,true,true,true),(true,false)) ../ocaml-vm/vm/mlvalue.ecl ../ocaml-vm/vm/fail.ecl ../ocaml-vm/vm/ram.ecl ../ocaml-vm/vm/runtime.ecl ../ocaml-vm/vm/debug.ecl ../ocaml-vm/vm/alloc.ecl ../ocaml-vm/vm/prims.ecl ../ocaml-vm/bytecode.ecl ../ocaml-vm/vm/vm.ecl ../ocaml-vm/vm/target-specific/intel-max10/IOs.ecl ../ocaml-vm/vm/target-specific/intel-max10/main.ecl

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.runtime.all;


entity main is
  
  port(signal clk    : in std_logic;
       signal reset  : in std_logic;
       signal argument : in value(0 to 11);
       signal result : out value(0 to 57));
       
end entity;
architecture rtl of main is

  type t_state is (IDLE4401, \$18437_LOOP666\, \$18438_LOOP665\, \$18439_WAIT662\, \$18440_MAKE_BLOCK579\, PAUSE_GET4405, PAUSE_GET4421, PAUSE_GET4425, PAUSE_GET4429, PAUSE_SET4402, PAUSE_SET4409, PAUSE_SET4412, PAUSE_SET4415, PAUSE_SET4418, PAUSE_SET4560, Q_WAIT4403, Q_WAIT4406, Q_WAIT4410, Q_WAIT4413, Q_WAIT4416, Q_WAIT4419, Q_WAIT4422, Q_WAIT4426, Q_WAIT4430, Q_WAIT4561);
  signal \state%now\, \state%next\: t_state;
  type t_state_var5924 is (IDLE4436, \$19779_LOOP666\, \$19780_LOOP665\, \$19781_AUX664\, \$19808_FOREVER6704342\, \$19811_COPY_ROOT_IN_RAM6634341\, \$19838_COPY_ROOT_IN_RAM6634340\, PAUSE_GET4440, PAUSE_GET4456, PAUSE_GET4460, PAUSE_GET4464, PAUSE_GET4468, PAUSE_GET4485, PAUSE_GET4489, PAUSE_GET4493, PAUSE_GET4497, PAUSE_GET4512, PAUSE_GET4516, PAUSE_GET4520, PAUSE_GET4533, PAUSE_GET4537, PAUSE_GET4550, PAUSE_GET4554, PAUSE_SET4437, PAUSE_SET4444, PAUSE_SET4447, PAUSE_SET4450, PAUSE_SET4453, PAUSE_SET4473, PAUSE_SET4476, PAUSE_SET4479, PAUSE_SET4482, PAUSE_SET4500, PAUSE_SET4503, PAUSE_SET4506, PAUSE_SET4509, PAUSE_SET4524, PAUSE_SET4527, PAUSE_SET4530, PAUSE_SET4541, PAUSE_SET4544, PAUSE_SET4547, Q_WAIT4438, Q_WAIT4441, Q_WAIT4445, Q_WAIT4448, Q_WAIT4451, Q_WAIT4454, Q_WAIT4457, Q_WAIT4461, Q_WAIT4465, Q_WAIT4469, Q_WAIT4474, Q_WAIT4477, Q_WAIT4480, Q_WAIT4483, Q_WAIT4486, Q_WAIT4490, Q_WAIT4494, Q_WAIT4498, Q_WAIT4501, Q_WAIT4504, Q_WAIT4507, Q_WAIT4510, Q_WAIT4513, Q_WAIT4517, Q_WAIT4521, Q_WAIT4525, Q_WAIT4528, Q_WAIT4531, Q_WAIT4534, Q_WAIT4538, Q_WAIT4542, Q_WAIT4545, Q_WAIT4548, Q_WAIT4551, Q_WAIT4555);
  signal \state_var5924%now\, \state_var5924%next\: t_state_var5924;
  type t_state_var5923 is (IDLE4609, \$18521_LOOP666\, \$18522_LOOP665\, \$18523_AUX664\, \$18524_LOOP666\, \$18525_LOOP665\, \$18526_AUX664\, \$18553_FOREVER6704348\, \$18556_FOREVER6704344\, \$18559_COPY_ROOT_IN_RAM6634347\, \$18571_COPY_ROOT_IN_RAM6634345\, \$18613_COPY_ROOT_IN_RAM6634346\, \$18625_COPY_ROOT_IN_RAM6634345\, PAUSE_GET4613, PAUSE_GET4629, PAUSE_GET4633, PAUSE_GET4637, PAUSE_GET4641, PAUSE_GET4648, PAUSE_GET4664, PAUSE_GET4668, PAUSE_GET4672, PAUSE_GET4676, PAUSE_GET4693, PAUSE_GET4697, PAUSE_GET4701, PAUSE_GET4717, PAUSE_GET4721, PAUSE_GET4725, PAUSE_GET4729, PAUSE_GET4744, PAUSE_GET4748, PAUSE_GET4752, PAUSE_GET4768, PAUSE_GET4772, PAUSE_GET4776, PAUSE_GET4789, PAUSE_GET4793, PAUSE_GET4806, PAUSE_GET4810, PAUSE_SET4610, PAUSE_SET4617, PAUSE_SET4620, PAUSE_SET4623, PAUSE_SET4626, PAUSE_SET4645, PAUSE_SET4652, PAUSE_SET4655, PAUSE_SET4658, PAUSE_SET4661, PAUSE_SET4681, PAUSE_SET4684, PAUSE_SET4687, PAUSE_SET4690, PAUSE_SET4705, PAUSE_SET4708, PAUSE_SET4711, PAUSE_SET4714, PAUSE_SET4732, PAUSE_SET4735, PAUSE_SET4738, PAUSE_SET4741, PAUSE_SET4756, PAUSE_SET4759, PAUSE_SET4762, PAUSE_SET4765, PAUSE_SET4780, PAUSE_SET4783, PAUSE_SET4786, PAUSE_SET4797, PAUSE_SET4800, PAUSE_SET4803, Q_WAIT4611, Q_WAIT4614, Q_WAIT4618, Q_WAIT4621, Q_WAIT4624, Q_WAIT4627, Q_WAIT4630, Q_WAIT4634, Q_WAIT4638, Q_WAIT4642, Q_WAIT4646, Q_WAIT4649, Q_WAIT4653, Q_WAIT4656, Q_WAIT4659, Q_WAIT4662, Q_WAIT4665, Q_WAIT4669, Q_WAIT4673, Q_WAIT4677, Q_WAIT4682, Q_WAIT4685, Q_WAIT4688, Q_WAIT4691, Q_WAIT4694, Q_WAIT4698, Q_WAIT4702, Q_WAIT4706, Q_WAIT4709, Q_WAIT4712, Q_WAIT4715, Q_WAIT4718, Q_WAIT4722, Q_WAIT4726, Q_WAIT4730, Q_WAIT4733, Q_WAIT4736, Q_WAIT4739, Q_WAIT4742, Q_WAIT4745, Q_WAIT4749, Q_WAIT4753, Q_WAIT4757, Q_WAIT4760, Q_WAIT4763, Q_WAIT4766, Q_WAIT4769, Q_WAIT4773, Q_WAIT4777, Q_WAIT4781, Q_WAIT4784, Q_WAIT4787, Q_WAIT4790, Q_WAIT4794, Q_WAIT4798, Q_WAIT4801, Q_WAIT4804, Q_WAIT4807, Q_WAIT4811);
  signal \state_var5923%now\, \state_var5923%next\: t_state_var5923;
  type t_state_var5922 is (IDLE4574, \$18466_LOOP666\, \$18467_LOOP665\, \$18468_WAIT662\, \$18469_MAKE_BLOCK579\, PAUSE_GET4578, PAUSE_GET4594, PAUSE_GET4598, PAUSE_GET4602, PAUSE_SET4575, PAUSE_SET4582, PAUSE_SET4585, PAUSE_SET4588, PAUSE_SET4591, PAUSE_SET4816, PAUSE_SET4819, PAUSE_SET4822, PAUSE_SET4825, PAUSE_SET4828, PAUSE_SET4831, PAUSE_SET4834, PAUSE_SET4837, PAUSE_SET4840, PAUSE_SET4843, PAUSE_SET4846, PAUSE_SET4849, PAUSE_SET4852, PAUSE_SET4855, PAUSE_SET4858, PAUSE_SET4861, PAUSE_SET4864, PAUSE_SET4867, PAUSE_SET4870, PAUSE_SET4873, PAUSE_SET4876, PAUSE_SET4879, PAUSE_SET4882, PAUSE_SET4885, PAUSE_SET4888, PAUSE_SET4891, PAUSE_SET4894, PAUSE_SET4897, PAUSE_SET4900, PAUSE_SET4903, PAUSE_SET4906, PAUSE_SET4909, PAUSE_SET4912, PAUSE_SET4915, PAUSE_SET4918, PAUSE_SET4921, PAUSE_SET4924, Q_WAIT4576, Q_WAIT4579, Q_WAIT4583, Q_WAIT4586, Q_WAIT4589, Q_WAIT4592, Q_WAIT4595, Q_WAIT4599, Q_WAIT4603, Q_WAIT4817, Q_WAIT4820, Q_WAIT4823, Q_WAIT4826, Q_WAIT4829, Q_WAIT4832, Q_WAIT4835, Q_WAIT4838, Q_WAIT4841, Q_WAIT4844, Q_WAIT4847, Q_WAIT4850, Q_WAIT4853, Q_WAIT4856, Q_WAIT4859, Q_WAIT4862, Q_WAIT4865, Q_WAIT4868, Q_WAIT4871, Q_WAIT4874, Q_WAIT4877, Q_WAIT4880, Q_WAIT4883, Q_WAIT4886, Q_WAIT4889, Q_WAIT4892, Q_WAIT4895, Q_WAIT4898, Q_WAIT4901, Q_WAIT4904, Q_WAIT4907, Q_WAIT4910, Q_WAIT4913, Q_WAIT4916, Q_WAIT4919, Q_WAIT4922, Q_WAIT4925);
  signal \state_var5922%now\, \state_var5922%next\: t_state_var5922;
  type t_state_var5921 is (IDLE4965, \$19494_LOOP666\, \$19495_LOOP665\, \$19496_AUX664\, \$19497_LOOP666\, \$19498_LOOP665\, \$19499_AUX664\, \$19526_FOREVER6704355\, \$19529_FOREVER6704351\, \$19532_FOREVER6704350\, \$19535_COPY_ROOT_IN_RAM6634354\, \$19547_COPY_ROOT_IN_RAM6634352\, \$19589_COPY_ROOT_IN_RAM6634353\, \$19601_COPY_ROOT_IN_RAM6634352\, PAUSE_GET4969, PAUSE_GET4985, PAUSE_GET4989, PAUSE_GET4993, PAUSE_GET4997, PAUSE_GET5004, PAUSE_GET5020, PAUSE_GET5024, PAUSE_GET5028, PAUSE_GET5032, PAUSE_GET5049, PAUSE_GET5053, PAUSE_GET5057, PAUSE_GET5073, PAUSE_GET5077, PAUSE_GET5081, PAUSE_GET5085, PAUSE_GET5100, PAUSE_GET5104, PAUSE_GET5108, PAUSE_GET5124, PAUSE_GET5128, PAUSE_GET5132, PAUSE_GET5145, PAUSE_GET5149, PAUSE_GET5162, PAUSE_GET5166, PAUSE_SET4966, PAUSE_SET4973, PAUSE_SET4976, PAUSE_SET4979, PAUSE_SET4982, PAUSE_SET5001, PAUSE_SET5008, PAUSE_SET5011, PAUSE_SET5014, PAUSE_SET5017, PAUSE_SET5037, PAUSE_SET5040, PAUSE_SET5043, PAUSE_SET5046, PAUSE_SET5061, PAUSE_SET5064, PAUSE_SET5067, PAUSE_SET5070, PAUSE_SET5088, PAUSE_SET5091, PAUSE_SET5094, PAUSE_SET5097, PAUSE_SET5112, PAUSE_SET5115, PAUSE_SET5118, PAUSE_SET5121, PAUSE_SET5136, PAUSE_SET5139, PAUSE_SET5142, PAUSE_SET5153, PAUSE_SET5156, PAUSE_SET5159, Q_WAIT4967, Q_WAIT4970, Q_WAIT4974, Q_WAIT4977, Q_WAIT4980, Q_WAIT4983, Q_WAIT4986, Q_WAIT4990, Q_WAIT4994, Q_WAIT4998, Q_WAIT5002, Q_WAIT5005, Q_WAIT5009, Q_WAIT5012, Q_WAIT5015, Q_WAIT5018, Q_WAIT5021, Q_WAIT5025, Q_WAIT5029, Q_WAIT5033, Q_WAIT5038, Q_WAIT5041, Q_WAIT5044, Q_WAIT5047, Q_WAIT5050, Q_WAIT5054, Q_WAIT5058, Q_WAIT5062, Q_WAIT5065, Q_WAIT5068, Q_WAIT5071, Q_WAIT5074, Q_WAIT5078, Q_WAIT5082, Q_WAIT5086, Q_WAIT5089, Q_WAIT5092, Q_WAIT5095, Q_WAIT5098, Q_WAIT5101, Q_WAIT5105, Q_WAIT5109, Q_WAIT5113, Q_WAIT5116, Q_WAIT5119, Q_WAIT5122, Q_WAIT5125, Q_WAIT5129, Q_WAIT5133, Q_WAIT5137, Q_WAIT5140, Q_WAIT5143, Q_WAIT5146, Q_WAIT5150, Q_WAIT5154, Q_WAIT5157, Q_WAIT5160, Q_WAIT5163, Q_WAIT5167);
  signal \state_var5921%now\, \state_var5921%next\: t_state_var5921;
  type t_state_var5920 is (IDLE4930, \$18790_LOOP666\, \$18791_LOOP665\, \$18792_WAIT662\, \$18793_MAKE_BLOCK579\, \$18794_APPLY638\, \$18795_OFFSETCLOSURE_N639\, \$18796_MAKE_BLOCK_N646\, \$18797_BRANCH_IF648\, \$18798_W652\, \$18799_W1656\, \$18856_LOOP_PUSH6494360\, \$18901_BINOP_INT6434361\, \$18907_MODULO6684356\, \$18910_MODULO6684349\, \$18914_MODULO6684357\, \$18917_MODULO6684349\, \$18920_BINOP_INT6434362\, \$18926_MODULO6684356\, \$18929_MODULO6684349\, \$18933_MODULO6684357\, \$18936_MODULO6684349\, \$18939_BINOP_INT6434363\, \$18945_MODULO6684356\, \$18948_MODULO6684349\, \$18952_MODULO6684357\, \$18955_MODULO6684349\, \$18958_BINOP_INT6434364\, \$18964_MODULO6684356\, \$18967_MODULO6684349\, \$18971_MODULO6684357\, \$18974_MODULO6684349\, \$18977_BINOP_INT6434365\, \$18983_MODULO6684356\, \$18986_MODULO6684349\, \$18990_MODULO6684357\, \$18993_MODULO6684349\, \$18996_BINOP_INT6434366\, \$19002_MODULO6684356\, \$19005_MODULO6684349\, \$19009_MODULO6684357\, \$19012_MODULO6684349\, \$19015_BINOP_INT6434367\, \$19021_MODULO6684356\, \$19024_MODULO6684349\, \$19028_MODULO6684357\, \$19031_MODULO6684349\, \$19034_BINOP_INT6434368\, \$19040_MODULO6684356\, \$19043_MODULO6684349\, \$19047_MODULO6684357\, \$19050_MODULO6684349\, \$19053_BINOP_INT6434369\, \$19059_MODULO6684356\, \$19062_MODULO6684349\, \$19066_MODULO6684357\, \$19069_MODULO6684349\, \$19072_BINOP_INT6434370\, \$19078_MODULO6684356\, \$19081_MODULO6684349\, \$19085_MODULO6684357\, \$19088_MODULO6684349\, \$19091_BINOP_INT6434371\, \$19097_MODULO6684356\, \$19100_MODULO6684349\, \$19104_MODULO6684357\, \$19107_MODULO6684349\, \$19113_FOREVER6704372\, \$19116_BINOP_INT6434373\, \$19122_MODULO6684356\, \$19125_MODULO6684349\, \$19129_MODULO6684357\, \$19132_MODULO6684349\, \$19135_BINOP_INT6434374\, \$19141_MODULO6684356\, \$19144_MODULO6684349\, \$19148_MODULO6684357\, \$19151_MODULO6684349\, \$19157_FOREVER6704375\, \$19163_FOREVER6704376\, \$19166_BINOP_COMPARE6454377\, \$19171_COMPARE6444358\, \$19174_BINOP_COMPARE6454378\, \$19179_COMPARE6444358\, \$19182_BINOP_COMPARE6454379\, \$19187_COMPARE6444358\, \$19190_BINOP_COMPARE6454380\, \$19195_COMPARE6444358\, \$19198_BINOP_COMPARE6454381\, \$19203_COMPARE6444358\, \$19206_BINOP_COMPARE6454382\, \$19211_COMPARE6444358\, \$19238_W6514383\, \$19252_FOREVER6704384\, \$19262_FOREVER6704385\, \$19320_FOREVER6704386\, \$19326_COMPBRANCH6504387\, \$19330_COMPARE6444359\, \$19333_COMPBRANCH6504388\, \$19337_COMPARE6444359\, \$19347_FILL6534389\, \$19361_FILL6544390\, \$19366_COMPBRANCH6504391\, \$19370_COMPARE6444359\, \$19373_COMPBRANCH6504392\, \$19377_COMPARE6444359\, \$19380_COMPBRANCH6504393\, \$19384_COMPARE6444359\, \$19387_COMPBRANCH6504394\, \$19391_COMPARE6444359\, \$19394_COMPBRANCH6504395\, \$19398_COMPARE6444359\, \$19401_COMPBRANCH6504396\, \$19405_COMPARE6444359\, \$19416_W36574398\, \$19420_W06554397\, PAUSE_GET4934, PAUSE_GET4950, PAUSE_GET4954, PAUSE_GET4958, PAUSE_GET5175, PAUSE_GET5200, PAUSE_GET5204, PAUSE_GET5208, PAUSE_GET5216, PAUSE_GET5223, PAUSE_GET5231, PAUSE_GET5238, PAUSE_GET5245, PAUSE_GET5252, PAUSE_GET5255, PAUSE_GET5258, PAUSE_GET5261, PAUSE_GET5264, PAUSE_GET5267, PAUSE_GET5270, PAUSE_GET5273, PAUSE_GET5282, PAUSE_GET5288, PAUSE_GET5294, PAUSE_GET5300, PAUSE_GET5306, PAUSE_GET5312, PAUSE_GET5318, PAUSE_GET5324, PAUSE_GET5327, PAUSE_GET5330, PAUSE_GET5333, PAUSE_GET5336, PAUSE_GET5342, PAUSE_GET5348, PAUSE_GET5354, PAUSE_GET5360, PAUSE_GET5366, PAUSE_GET5370, PAUSE_GET5385, PAUSE_GET5388, PAUSE_GET5391, PAUSE_GET5394, PAUSE_GET5400, PAUSE_GET5406, PAUSE_GET5412, PAUSE_GET5418, PAUSE_GET5421, PAUSE_GET5424, PAUSE_GET5427, PAUSE_GET5433, PAUSE_GET5436, PAUSE_GET5439, PAUSE_GET5442, PAUSE_GET5448, PAUSE_GET5451, PAUSE_GET5454, PAUSE_GET5457, PAUSE_GET5460, PAUSE_GET5463, PAUSE_GET5466, PAUSE_GET5488, PAUSE_GET5498, PAUSE_GET5508, PAUSE_GET5518, PAUSE_GET5528, PAUSE_GET5538, PAUSE_GET5548, PAUSE_GET5558, PAUSE_GET5568, PAUSE_GET5578, PAUSE_GET5588, PAUSE_GET5598, PAUSE_GET5608, PAUSE_GET5612, PAUSE_GET5616, PAUSE_GET5620, PAUSE_GET5624, PAUSE_GET5628, PAUSE_GET5632, PAUSE_GET5635, PAUSE_GET5638, PAUSE_GET5647, PAUSE_GET5650, PAUSE_GET5665, PAUSE_GET5668, PAUSE_GET5671, PAUSE_GET5674, PAUSE_GET5677, PAUSE_GET5681, PAUSE_GET5684, PAUSE_GET5687, PAUSE_GET5693, PAUSE_GET5707, PAUSE_GET5710, PAUSE_GET5722, PAUSE_GET5728, PAUSE_GET5731, PAUSE_GET5734, PAUSE_GET5750, PAUSE_GET5757, PAUSE_GET5764, PAUSE_GET5767, PAUSE_GET5774, PAUSE_GET5777, PAUSE_GET5780, PAUSE_GET5787, PAUSE_GET5790, PAUSE_GET5793, PAUSE_GET5796, PAUSE_GET5803, PAUSE_GET5806, PAUSE_GET5809, PAUSE_GET5812, PAUSE_GET5821, PAUSE_GET5826, PAUSE_GET5832, PAUSE_GET5843, PAUSE_GET5846, PAUSE_GET5849, PAUSE_GET5852, PAUSE_GET5861, PAUSE_GET5884, PAUSE_GET5895, PAUSE_GET5899, PAUSE_GET5903, PAUSE_GET5907, PAUSE_GET5911, PAUSE_SET4931, PAUSE_SET4938, PAUSE_SET4941, PAUSE_SET4944, PAUSE_SET4947, PAUSE_SET5172, PAUSE_SET5178, PAUSE_SET5182, PAUSE_SET5186, PAUSE_SET5190, PAUSE_SET5193, PAUSE_SET5196, PAUSE_SET5213, PAUSE_SET5220, PAUSE_SET5227, PAUSE_SET5235, PAUSE_SET5242, PAUSE_SET5248, PAUSE_SET5276, PAUSE_SET5279, PAUSE_SET5285, PAUSE_SET5291, PAUSE_SET5297, PAUSE_SET5303, PAUSE_SET5309, PAUSE_SET5315, PAUSE_SET5321, PAUSE_SET5339, PAUSE_SET5345, PAUSE_SET5351, PAUSE_SET5357, PAUSE_SET5363, PAUSE_SET5373, PAUSE_SET5376, PAUSE_SET5379, PAUSE_SET5382, PAUSE_SET5397, PAUSE_SET5403, PAUSE_SET5409, PAUSE_SET5415, PAUSE_SET5430, PAUSE_SET5445, PAUSE_SET5469, PAUSE_SET5472, PAUSE_SET5475, PAUSE_SET5478, PAUSE_SET5641, PAUSE_SET5644, PAUSE_SET5653, PAUSE_SET5656, PAUSE_SET5659, PAUSE_SET5662, PAUSE_SET5690, PAUSE_SET5697, PAUSE_SET5700, PAUSE_SET5704, PAUSE_SET5713, PAUSE_SET5716, PAUSE_SET5719, PAUSE_SET5725, PAUSE_SET5738, PAUSE_SET5741, PAUSE_SET5744, PAUSE_SET5747, PAUSE_SET5754, PAUSE_SET5761, PAUSE_SET5771, PAUSE_SET5784, PAUSE_SET5800, PAUSE_SET5815, PAUSE_SET5818, PAUSE_SET5829, PAUSE_SET5836, PAUSE_SET5839, PAUSE_SET5855, PAUSE_SET5858, PAUSE_SET5865, PAUSE_SET5874, PAUSE_SET5878, PAUSE_SET5881, PAUSE_SET5888, PAUSE_SET5891, Q_WAIT4932, Q_WAIT4935, Q_WAIT4939, Q_WAIT4942, Q_WAIT4945, Q_WAIT4948, Q_WAIT4951, Q_WAIT4955, Q_WAIT4959, Q_WAIT5173, Q_WAIT5176, Q_WAIT5179, Q_WAIT5183, Q_WAIT5187, Q_WAIT5191, Q_WAIT5194, Q_WAIT5197, Q_WAIT5201, Q_WAIT5205, Q_WAIT5209, Q_WAIT5214, Q_WAIT5217, Q_WAIT5221, Q_WAIT5224, Q_WAIT5228, Q_WAIT5232, Q_WAIT5236, Q_WAIT5239, Q_WAIT5243, Q_WAIT5246, Q_WAIT5249, Q_WAIT5253, Q_WAIT5256, Q_WAIT5259, Q_WAIT5262, Q_WAIT5265, Q_WAIT5268, Q_WAIT5271, Q_WAIT5274, Q_WAIT5277, Q_WAIT5280, Q_WAIT5283, Q_WAIT5286, Q_WAIT5289, Q_WAIT5292, Q_WAIT5295, Q_WAIT5298, Q_WAIT5301, Q_WAIT5304, Q_WAIT5307, Q_WAIT5310, Q_WAIT5313, Q_WAIT5316, Q_WAIT5319, Q_WAIT5322, Q_WAIT5325, Q_WAIT5328, Q_WAIT5331, Q_WAIT5334, Q_WAIT5337, Q_WAIT5340, Q_WAIT5343, Q_WAIT5346, Q_WAIT5349, Q_WAIT5352, Q_WAIT5355, Q_WAIT5358, Q_WAIT5361, Q_WAIT5364, Q_WAIT5367, Q_WAIT5371, Q_WAIT5374, Q_WAIT5377, Q_WAIT5380, Q_WAIT5383, Q_WAIT5386, Q_WAIT5389, Q_WAIT5392, Q_WAIT5395, Q_WAIT5398, Q_WAIT5401, Q_WAIT5404, Q_WAIT5407, Q_WAIT5410, Q_WAIT5413, Q_WAIT5416, Q_WAIT5419, Q_WAIT5422, Q_WAIT5425, Q_WAIT5428, Q_WAIT5431, Q_WAIT5434, Q_WAIT5437, Q_WAIT5440, Q_WAIT5443, Q_WAIT5446, Q_WAIT5449, Q_WAIT5452, Q_WAIT5455, Q_WAIT5458, Q_WAIT5461, Q_WAIT5464, Q_WAIT5467, Q_WAIT5470, Q_WAIT5473, Q_WAIT5476, Q_WAIT5479, Q_WAIT5489, Q_WAIT5499, Q_WAIT5509, Q_WAIT5519, Q_WAIT5529, Q_WAIT5539, Q_WAIT5549, Q_WAIT5559, Q_WAIT5569, Q_WAIT5579, Q_WAIT5589, Q_WAIT5599, Q_WAIT5609, Q_WAIT5613, Q_WAIT5617, Q_WAIT5621, Q_WAIT5625, Q_WAIT5629, Q_WAIT5633, Q_WAIT5636, Q_WAIT5639, Q_WAIT5642, Q_WAIT5645, Q_WAIT5648, Q_WAIT5651, Q_WAIT5654, Q_WAIT5657, Q_WAIT5660, Q_WAIT5663, Q_WAIT5666, Q_WAIT5669, Q_WAIT5672, Q_WAIT5675, Q_WAIT5678, Q_WAIT5682, Q_WAIT5685, Q_WAIT5688, Q_WAIT5691, Q_WAIT5694, Q_WAIT5698, Q_WAIT5701, Q_WAIT5705, Q_WAIT5708, Q_WAIT5711, Q_WAIT5714, Q_WAIT5717, Q_WAIT5720, Q_WAIT5723, Q_WAIT5726, Q_WAIT5729, Q_WAIT5732, Q_WAIT5735, Q_WAIT5739, Q_WAIT5742, Q_WAIT5745, Q_WAIT5748, Q_WAIT5751, Q_WAIT5755, Q_WAIT5758, Q_WAIT5762, Q_WAIT5765, Q_WAIT5768, Q_WAIT5772, Q_WAIT5775, Q_WAIT5778, Q_WAIT5781, Q_WAIT5785, Q_WAIT5788, Q_WAIT5791, Q_WAIT5794, Q_WAIT5797, Q_WAIT5801, Q_WAIT5804, Q_WAIT5807, Q_WAIT5810, Q_WAIT5813, Q_WAIT5816, Q_WAIT5819, Q_WAIT5822, Q_WAIT5827, Q_WAIT5830, Q_WAIT5833, Q_WAIT5837, Q_WAIT5840, Q_WAIT5844, Q_WAIT5847, Q_WAIT5850, Q_WAIT5853, Q_WAIT5856, Q_WAIT5859, Q_WAIT5862, Q_WAIT5866, Q_WAIT5875, Q_WAIT5879, Q_WAIT5882, Q_WAIT5885, Q_WAIT5889, Q_WAIT5892, Q_WAIT5896, Q_WAIT5900, Q_WAIT5904, Q_WAIT5908, Q_WAIT5912);
  signal \state_var5920%now\, \state_var5920%next\: t_state_var5920;
  type array_value_16 is array (natural range <>) of value(0 to 15);
  type array_value_31 is array (natural range <>) of value(0 to 30);
  type array_value_32 is array (natural range <>) of value(0 to 31);
  signal ram : array_value_32(0 to 16383);
  signal \$ram_value\ : value(0 to 31) := (others => '0');
  signal \$ram_ptr\ : natural range 0 to 16383 := 0;
  signal \$ram_ptr_write\ : natural range 0 to 16383 := 0;
  signal \$ram_write\ : value(0 to 31) := (others => '0');
  signal \$ram_write_request\ : std_logic := '0';
  signal global_end : array_value_16(0 to 0);
  signal \$global_end_value\ : value(0 to 15) := (others => '0');
  signal \$global_end_ptr\ : natural range 0 to 0 := 0;
  signal \$global_end_ptr_write\ : natural range 0 to 0 := 0;
  signal \$global_end_write\ : value(0 to 15) := (others => '0');
  signal \$global_end_write_request\ : std_logic := '0';
  signal code : array_value_31(0 to 34);
  signal \$code_value\ : value(0 to 30) := (others => '0');
  signal \$code_ptr\ : natural range 0 to 34 := 0;
  signal \$code_ptr_write\ : natural range 0 to 34 := 0;
  signal \$code_write\ : value(0 to 30) := (others => '0');
  signal \$code_write_request\ : std_logic := '0';
  signal \$18463%next\, \$18463%now\ : value(0 to 1) := (others => '0');
  signal \$19410%next\, \$19410%now\, \$18469_make_block579_result%next\, 
         \$18469_make_block579_result%now\, \$19420_w06554397_arg%next\, 
         \$19420_w06554397_arg%now\, \$18440_make_block579_result%next\, 
         \$18440_make_block579_result%now\, \$19344%next\, \$19344%now\, 
         \$18525_loop665_arg%next\, \$18525_loop665_arg%now\, \$19231%next\, 
         \$19231%now\, \$18438_loop665_arg%next\, \$18438_loop665_arg%now\, 
         \$18522_loop665_arg%next\, \$18522_loop665_arg%now\, \$19444%next\, 
         \$19444%now\, \$19498_loop665_arg%next\, \$19498_loop665_arg%now\, 
         \$18467_loop665_arg%next\, \$18467_loop665_arg%now\, 
         \$18791_loop665_arg%next\, \$18791_loop665_arg%now\, 
         \$19780_loop665_arg%next\, \$19780_loop665_arg%now\, 
         \$19495_loop665_arg%next\, \$19495_loop665_arg%now\, \$19358%next\, 
         \$19358%now\, \$18793_make_block579_result%next\, 
         \$18793_make_block579_result%now\ : value(0 to 95) := (others => '0');
  signal \$19195_compare6444358_arg%next\, \$19195_compare6444358_arg%now\, 
         \$19330_compare6444359_arg%next\, \$19330_compare6444359_arg%now\, 
         \$19398_compare6444359_arg%next\, \$19398_compare6444359_arg%now\, 
         \$19384_compare6444359_arg%next\, \$19384_compare6444359_arg%now\, 
         \$19377_compare6444359_arg%next\, \$19377_compare6444359_arg%now\, 
         \$19370_compare6444359_arg%next\, \$19370_compare6444359_arg%now\, 
         \$19171_compare6444358_arg%next\, \$19171_compare6444358_arg%now\, 
         \$19391_compare6444359_arg%next\, \$19391_compare6444359_arg%now\, 
         \$19203_compare6444358_arg%next\, \$19203_compare6444358_arg%now\, 
         \$19405_compare6444359_arg%next\, \$19405_compare6444359_arg%now\, 
         \$19211_compare6444358_arg%next\, \$19211_compare6444358_arg%now\, 
         \$19337_compare6444359_arg%next\, \$19337_compare6444359_arg%now\, 
         \$19187_compare6444358_arg%next\, \$19187_compare6444358_arg%now\, 
         \$19179_compare6444358_arg%next\, \$19179_compare6444358_arg%now\ : value(0 to 93) := (others => '0');
  signal \$19742%next\, \$19742%now\, \$19608%next\, \$19608%now\, 
         \$18632%next\, \$18632%now\, \$18532%next\, \$18532%now\, 
         \$19506%next\, \$19506%now\, \$19931%next\, \$19931%now\, 
         \$18448_dis%next\, \$18448_dis%now\, \$18766%next\, \$18766%now\, 
         \$18533%next\, \$18533%now\, \$19462%next\, \$19462%now\, 
         \$19907%next\, \$19907%now\, \$19818%next\, \$19818%now\, 
         \$19788%next\, \$19788%now\, \$19542%next\, \$19542%now\, 
         \$19787%next\, \$19787%now\, \$19554%next\, \$19554%now\, 
         \$19718%next\, \$19718%now\, \$19463%next\, \$19463%now\, 
         \$18742%next\, \$18742%now\, \$19505%next\, \$19505%now\, 
         \$19596%next\, \$19596%now\, \$18566%next\, \$18566%now\, 
         \$19845%next\, \$19845%now\, \$18709%next\, \$18709%now\, 
         \$18620%next\, \$18620%now\, \$18578%next\, \$18578%now\, 
         \$19685%next\, \$19685%now\, \$19464%next\, \$19464%now\ : value(0 to 47) := (others => '0');
  signal \$18790_loop666_arg%next\, \$18790_loop666_arg%now\, 
         \$18523_aux664_arg%next\, \$18523_aux664_arg%now\, 
         \$18798_w652_arg%next\, \$18798_w652_arg%now\, 
         \$18466_loop666_arg%next\, \$18466_loop666_arg%now\, 
         \$19494_loop666_arg%next\, \$19494_loop666_arg%now\, 
         \$19781_aux664_arg%next\, \$19781_aux664_arg%now\, 
         \$19497_loop666_arg%next\, \$19497_loop666_arg%now\, 
         \$18524_loop666_arg%next\, \$18524_loop666_arg%now\, 
         \$18437_loop666_arg%next\, \$18437_loop666_arg%now\, 
         \$18526_aux664_arg%next\, \$18526_aux664_arg%now\, 
         \$19499_aux664_arg%next\, \$19499_aux664_arg%now\, 
         \$18856_loop_push6494360_arg%next\, 
         \$18856_loop_push6494360_arg%now\, \$19779_loop666_arg%next\, 
         \$19779_loop666_arg%now\, \$19238_w6514383_arg%next\, 
         \$19238_w6514383_arg%now\, \$19496_aux664_arg%next\, 
         \$19496_aux664_arg%now\, \$18521_loop666_arg%next\, 
         \$18521_loop666_arg%now\ : value(0 to 63) := (others => '0');
  signal \$18452%next\, \$18452%now\, \$18451%next\, \$18451%now\, 
         \$18454%next\, \$18454%now\, \$v5902%next\, \$v5902%now\, 
         \$v5910%next\, \$v5910%now\, \$v5898%next\, \$v5898%now\, 
         \$v5906%next\, \$v5906%now\, \$18453%next\, \$18453%now\, 
         \$18456%next\, \$18456%now\, \$18455%next\, \$18455%now\ : value(0 to 7) := (others => '0');
  signal \$18797_branch_if648_arg%next\, \$18797_branch_if648_arg%now\, 
         \$18787%next\, \$18787%now\, \$18789%next\, \$18789%now\, 
         \$18788%next\, \$18788%now\ : value(0 to 122) := (others => '0');
  signal \$18541%next\, \$18541%now\, \$19360_sp%next\, \$19360_sp%now\, 
         \$19415_sp%next\, \$19415_sp%now\, \$19499_aux664_result%next\, 
         \$19499_aux664_result%now\, \$18705_next%next\, \$18705_next%now\, 
         \$19780_loop665_result%next\, \$19780_loop665_result%now\, 
         \$19343_sp%next\, \$19343_sp%now\, \$19446_sp%next\, 
         \$19446_sp%now\, \$18526_aux664_result%next\, 
         \$18526_aux664_result%now\, \$19465_sp%next\, \$19465_sp%now\, 
         \$18625_copy_root_in_ram6634345_result%next\, 
         \$18625_copy_root_in_ram6634345_result%now\, \$19468_sp%next\, 
         \$19468_sp%now\, \$19265_ofs%next\, \$19265_ofs%now\, 
         \$18534_next%next\, \$18534_next%now\, 
         \$18856_loop_push6494360_result%next\, 
         \$18856_loop_push6494360_result%now\, \$19903_next%next\, 
         \$19903_next%now\, \$19346_sp%next\, \$19346_sp%now\, 
         \$18523_aux664_result%next\, \$18523_aux664_result%now\, 
         \$19781_aux664_result%next\, \$19781_aux664_result%now\, 
         \$19535_copy_root_in_ram6634354_result%next\, 
         \$19535_copy_root_in_ram6634354_result%now\, \$19514%next\, 
         \$19514%now\, \$19347_fill6534389_result%next\, 
         \$19347_fill6534389_result%now\, \$18467_loop665_result%next\, 
         \$18467_loop665_result%now\, \$19518_next%next\, \$19518_next%now\, 
         \$18571_copy_root_in_ram6634345_result%next\, 
         \$18571_copy_root_in_ram6634345_result%now\, 
         \$18438_loop665_result%next\, \$18438_loop665_result%now\, 
         \$18522_loop665_result%next\, \$18522_loop665_result%now\, 
         \$18542_next%next\, \$18542_next%now\, \$19447_sp%next\, 
         \$19447_sp%now\, \$18545_next%next\, \$18545_next%now\, 
         \$19811_copy_root_in_ram6634341_result%next\, 
         \$19811_copy_root_in_ram6634341_result%now\, \$19234_sp%next\, 
         \$19234_sp%now\, \$19409_sp%next\, \$19409_sp%now\, 
         \$19498_loop665_result%next\, \$19498_loop665_result%now\, 
         \$19466_sp%next\, \$19466_sp%now\, \$19796%next\, \$19796%now\, 
         \$19789_next%next\, \$19789_next%now\, \$19507_next%next\, 
         \$19507_next%now\, \$19496_aux664_result%next\, 
         \$19496_aux664_result%now\, \$19412_sp%next\, \$19412_sp%now\, 
         \$19420_w06554397_result%next\, \$19420_w06554397_result%now\, 
         \$19589_copy_root_in_ram6634353_result%next\, 
         \$19589_copy_root_in_ram6634353_result%now\, \$18854_sp%next\, 
         \$18854_sp%now\, \$19467_sp%next\, \$19467_sp%now\, 
         \$18613_copy_root_in_ram6634346_result%next\, 
         \$18613_copy_root_in_ram6634346_result%now\, 
         \$19361_fill6544390_result%next\, \$19361_fill6544390_result%now\, 
         \$19601_copy_root_in_ram6634352_result%next\, 
         \$19601_copy_root_in_ram6634352_result%now\, 
         \$18791_loop665_result%next\, \$18791_loop665_result%now\, 
         \$19238_w6514383_result%next\, \$19238_w6514383_result%now\, 
         \$18525_loop665_result%next\, \$18525_loop665_result%now\, 
         \$19681_next%next\, \$19681_next%now\, 
         \$19547_copy_root_in_ram6634352_result%next\, 
         \$19547_copy_root_in_ram6634352_result%now\, 
         \$18559_copy_root_in_ram6634347_result%next\, 
         \$18559_copy_root_in_ram6634347_result%now\, \$19800_next%next\, 
         \$19800_next%now\, \$19495_loop665_result%next\, 
         \$19495_loop665_result%now\, \$19515_next%next\, \$19515_next%now\, 
         \$19838_copy_root_in_ram6634340_result%next\, 
         \$19838_copy_root_in_ram6634340_result%now\, \$19714_next%next\, 
         \$19714_next%now\, \$19797_next%next\, \$19797_next%now\, 
         \$18738_next%next\, \$18738_next%now\, 
         \$19416_w36574398_result%next\, \$19416_w36574398_result%now\ : value(0 to 15) := (others => '0');
  signal \$18926_modulo6684356_arg%next\, \$18926_modulo6684356_arg%now\, 
         \$19125_modulo6684349_arg%next\, \$19125_modulo6684349_arg%now\, 
         \$18955_modulo6684349_arg%next\, \$18955_modulo6684349_arg%now\, 
         \$18910_modulo6684349_arg%next\, \$18910_modulo6684349_arg%now\, 
         \$19050_modulo6684349_arg%next\, \$19050_modulo6684349_arg%now\, 
         \$19028_modulo6684357_arg%next\, \$19028_modulo6684357_arg%now\, 
         \$18990_modulo6684357_arg%next\, \$18990_modulo6684357_arg%now\, 
         \$19122_modulo6684356_arg%next\, \$19122_modulo6684356_arg%now\, 
         \$19144_modulo6684349_arg%next\, \$19144_modulo6684349_arg%now\, 
         \$19047_modulo6684357_arg%next\, \$19047_modulo6684357_arg%now\, 
         \$18983_modulo6684356_arg%next\, \$18983_modulo6684356_arg%now\, 
         \$19151_modulo6684349_arg%next\, \$19151_modulo6684349_arg%now\, 
         \$19024_modulo6684349_arg%next\, \$19024_modulo6684349_arg%now\, 
         \$19012_modulo6684349_arg%next\, \$19012_modulo6684349_arg%now\, 
         \$18964_modulo6684356_arg%next\, \$18964_modulo6684356_arg%now\, 
         \$19040_modulo6684356_arg%next\, \$19040_modulo6684356_arg%now\, 
         \$19062_modulo6684349_arg%next\, \$19062_modulo6684349_arg%now\, 
         \$19132_modulo6684349_arg%next\, \$19132_modulo6684349_arg%now\, 
         \$19021_modulo6684356_arg%next\, \$19021_modulo6684356_arg%now\, 
         \$19031_modulo6684349_arg%next\, \$19031_modulo6684349_arg%now\, 
         \$18917_modulo6684349_arg%next\, \$18917_modulo6684349_arg%now\, 
         \$19104_modulo6684357_arg%next\, \$19104_modulo6684357_arg%now\, 
         \$19009_modulo6684357_arg%next\, \$19009_modulo6684357_arg%now\, 
         \$18929_modulo6684349_arg%next\, \$18929_modulo6684349_arg%now\, 
         \$18971_modulo6684357_arg%next\, \$18971_modulo6684357_arg%now\, 
         \$19141_modulo6684356_arg%next\, \$19141_modulo6684356_arg%now\, 
         \$19097_modulo6684356_arg%next\, \$19097_modulo6684356_arg%now\, 
         \$19100_modulo6684349_arg%next\, \$19100_modulo6684349_arg%now\, 
         \$19005_modulo6684349_arg%next\, \$19005_modulo6684349_arg%now\, 
         \$19085_modulo6684357_arg%next\, \$19085_modulo6684357_arg%now\, 
         \$19148_modulo6684357_arg%next\, \$19148_modulo6684357_arg%now\, 
         \$19078_modulo6684356_arg%next\, \$19078_modulo6684356_arg%now\, 
         \$19107_modulo6684349_arg%next\, \$19107_modulo6684349_arg%now\, 
         \$19129_modulo6684357_arg%next\, \$19129_modulo6684357_arg%now\, 
         \$18907_modulo6684356_arg%next\, \$18907_modulo6684356_arg%now\, 
         \$19069_modulo6684349_arg%next\, \$19069_modulo6684349_arg%now\, 
         \$19059_modulo6684356_arg%next\, \$19059_modulo6684356_arg%now\, 
         \$19088_modulo6684349_arg%next\, \$19088_modulo6684349_arg%now\, 
         \$18952_modulo6684357_arg%next\, \$18952_modulo6684357_arg%now\, 
         \$18933_modulo6684357_arg%next\, \$18933_modulo6684357_arg%now\, 
         \$19066_modulo6684357_arg%next\, \$19066_modulo6684357_arg%now\, 
         \$18936_modulo6684349_arg%next\, \$18936_modulo6684349_arg%now\, 
         \$18967_modulo6684349_arg%next\, \$18967_modulo6684349_arg%now\, 
         \$19043_modulo6684349_arg%next\, \$19043_modulo6684349_arg%now\, 
         \$18948_modulo6684349_arg%next\, \$18948_modulo6684349_arg%now\, 
         \$18914_modulo6684357_arg%next\, \$18914_modulo6684357_arg%now\, 
         \$18993_modulo6684349_arg%next\, \$18993_modulo6684349_arg%now\, 
         \$18986_modulo6684349_arg%next\, \$18986_modulo6684349_arg%now\, 
         \$19002_modulo6684356_arg%next\, \$19002_modulo6684356_arg%now\, 
         \$18974_modulo6684349_arg%next\, \$18974_modulo6684349_arg%now\, 
         \$19081_modulo6684349_arg%next\, \$19081_modulo6684349_arg%now\, 
         \$18945_modulo6684356_arg%next\, \$18945_modulo6684356_arg%now\ : value(0 to 61) := (others => '0');
  signal \$18468_wait662_arg%next\, \$18468_wait662_arg%now\, 
         \$18792_wait662_arg%next\, \$18792_wait662_arg%now\, 
         \$18439_wait662_arg%next\, \$18439_wait662_arg%now\ : value(0 to 96) := (others => '0');
  signal \result4399%next\, \result4399%now\ : value(0 to 57) := (others => '0');
  signal \$v4564%next\, \$v4564%now\, \$v4566%next\, \$v4566%now\, 
         \$v4567%next\, \$v4567%now\, \$18443%next\, \$18443%now\, 
         \$18462%next\, \$18462%now\, \$v4565%next\, \$v4565%now\, 
         \$v4568%next\, \$v4568%now\, \$v4563%next\, \$v4563%now\ : value(0 to 3) := (others => '0');
  signal \$19380_compbranch6504393_arg%next\, 
         \$19380_compbranch6504393_arg%now\, 
         \$19373_compbranch6504392_arg%next\, 
         \$19373_compbranch6504392_arg%now\, 
         \$19401_compbranch6504396_arg%next\, 
         \$19401_compbranch6504396_arg%now\, 
         \$19387_compbranch6504394_arg%next\, 
         \$19387_compbranch6504394_arg%now\, 
         \$19366_compbranch6504391_arg%next\, 
         \$19366_compbranch6504391_arg%now\, 
         \$19326_compbranch6504387_arg%next\, 
         \$19326_compbranch6504387_arg%now\, 
         \$19333_compbranch6504388_arg%next\, 
         \$19333_compbranch6504388_arg%now\, 
         \$19394_compbranch6504395_arg%next\, 
         \$19394_compbranch6504395_arg%now\ : value(0 to 215) := (others => '0');
  signal \$18952_modulo6684357_id%next\, \$18952_modulo6684357_id%now\, 
         \$19107_modulo6684349_id%next\, \$19107_modulo6684349_id%now\, 
         \$19141_modulo6684356_id%next\, \$19141_modulo6684356_id%now\, 
         \$18917_modulo6684349_id%next\, \$18917_modulo6684349_id%now\, 
         \$19347_fill6534389_id%next\, \$19347_fill6534389_id%now\, 
         \$18901_binop_int6434361_id%next\, \$18901_binop_int6434361_id%now\, 
         \$19085_modulo6684357_id%next\, \$19085_modulo6684357_id%now\, 
         \$18798_w652_id%next\, \$18798_w652_id%now\, 
         \$19416_w36574398_id%next\, \$19416_w36574398_id%now\, 
         \$19198_binop_compare6454381_id%next\, 
         \$19198_binop_compare6454381_id%now\, 
         \$18929_modulo6684349_id%next\, \$18929_modulo6684349_id%now\, 
         \$19498_loop665_id%next\, \$19498_loop665_id%now\, 
         \$19405_compare6444359_id%next\, \$19405_compare6444359_id%now\, 
         \$19009_modulo6684357_id%next\, \$19009_modulo6684357_id%now\, 
         \$18524_loop666_id%next\, \$18524_loop666_id%now\, 
         \$18967_modulo6684349_id%next\, \$18967_modulo6684349_id%now\, 
         \$19116_binop_int6434373_id%next\, \$19116_binop_int6434373_id%now\, 
         \$18792_wait662_id%next\, \$18792_wait662_id%now\, 
         \$19034_binop_int6434368_id%next\, \$19034_binop_int6434368_id%now\, 
         \$18468_wait662_id%next\, \$18468_wait662_id%now\, 
         \$18986_modulo6684349_id%next\, \$18986_modulo6684349_id%now\, 
         \$19195_compare6444358_id%next\, \$19195_compare6444358_id%now\, 
         \$19377_compare6444359_id%next\, \$19377_compare6444359_id%now\, 
         \$18920_binop_int6434362_id%next\, \$18920_binop_int6434362_id%now\, 
         \$18983_modulo6684356_id%next\, \$18983_modulo6684356_id%now\, 
         \$19401_compbranch6504396_id%next\, 
         \$19401_compbranch6504396_id%now\, 
         \$19206_binop_compare6454382_id%next\, 
         \$19206_binop_compare6454382_id%now\, 
         \$19050_modulo6684349_id%next\, \$19050_modulo6684349_id%now\, 
         \$19151_modulo6684349_id%next\, \$19151_modulo6684349_id%now\, 
         \$19002_modulo6684356_id%next\, \$19002_modulo6684356_id%now\, 
         \$19053_binop_int6434369_id%next\, \$19053_binop_int6434369_id%now\, 
         \$19529_forever6704351_id%next\, \$19529_forever6704351_id%now\, 
         \$19494_loop666_id%next\, \$19494_loop666_id%now\, 
         \$19808_forever6704342_id%next\, \$19808_forever6704342_id%now\, 
         \$19373_compbranch6504392_id%next\, 
         \$19373_compbranch6504392_id%now\, \$19122_modulo6684356_id%next\, 
         \$19122_modulo6684356_id%now\, 
         \$19838_copy_root_in_ram6634340_id%next\, 
         \$19838_copy_root_in_ram6634340_id%now\, \$19780_loop665_id%next\, 
         \$19780_loop665_id%now\, \$19174_binop_compare6454378_id%next\, 
         \$19174_binop_compare6454378_id%now\, 
         \$19366_compbranch6504391_id%next\, 
         \$19366_compbranch6504391_id%now\, 
         \$18856_loop_push6494360_id%next\, \$18856_loop_push6494360_id%now\, 
         \$19394_compbranch6504395_id%next\, 
         \$19394_compbranch6504395_id%now\, \$19081_modulo6684349_id%next\, 
         \$19081_modulo6684349_id%now\, \$18955_modulo6684349_id%next\, 
         \$18955_modulo6684349_id%now\, \$19398_compare6444359_id%next\, 
         \$19398_compare6444359_id%now\, \$19059_modulo6684356_id%next\, 
         \$19059_modulo6684356_id%now\, \$19420_w06554397_id%next\, 
         \$19420_w06554397_id%now\, \$19135_binop_int6434374_id%next\, 
         \$19135_binop_int6434374_id%now\, 
         \$19547_copy_root_in_ram6634352_id%next\, 
         \$19547_copy_root_in_ram6634352_id%now\, 
         \$19182_binop_compare6454379_id%next\, 
         \$19182_binop_compare6454379_id%now\, 
         \$19148_modulo6684357_id%next\, \$19148_modulo6684357_id%now\, 
         \$19113_forever6704372_id%next\, \$19113_forever6704372_id%now\, 
         \$19072_binop_int6434370_id%next\, \$19072_binop_int6434370_id%now\, 
         \$18439_wait662_id%next\, \$18439_wait662_id%now\, 
         \$18556_forever6704344_id%next\, \$18556_forever6704344_id%now\, 
         \$18625_copy_root_in_ram6634345_id%next\, 
         \$18625_copy_root_in_ram6634345_id%now\, 
         \$19252_forever6704384_id%next\, \$19252_forever6704384_id%now\, 
         \$19024_modulo6684349_id%next\, \$19024_modulo6684349_id%now\, 
         \$19781_aux664_id%next\, \$19781_aux664_id%now\, 
         \$18914_modulo6684357_id%next\, \$18914_modulo6684357_id%now\, 
         \$19005_modulo6684349_id%next\, \$19005_modulo6684349_id%now\, 
         \$19166_binop_compare6454377_id%next\, 
         \$19166_binop_compare6454377_id%now\, 
         \$18553_forever6704348_id%next\, \$18553_forever6704348_id%now\, 
         \$19526_forever6704355_id%next\, \$19526_forever6704355_id%now\, 
         \$19031_modulo6684349_id%next\, \$19031_modulo6684349_id%now\, 
         \$19047_modulo6684357_id%next\, \$19047_modulo6684357_id%now\, 
         \$18525_loop665_id%next\, \$18525_loop665_id%now\, 
         \$19091_binop_int6434371_id%next\, \$19091_binop_int6434371_id%now\, 
         \$19028_modulo6684357_id%next\, \$19028_modulo6684357_id%now\, 
         \$18795_offsetclosure_n639_id%next\, 
         \$18795_offsetclosure_n639_id%now\, \$19125_modulo6684349_id%next\, 
         \$19125_modulo6684349_id%now\, 
         \$18559_copy_root_in_ram6634347_id%next\, 
         \$18559_copy_root_in_ram6634347_id%now\, 
         \$19100_modulo6684349_id%next\, \$19100_modulo6684349_id%now\, 
         \$18948_modulo6684349_id%next\, \$18948_modulo6684349_id%now\, 
         \$19361_fill6544390_id%next\, \$19361_fill6544390_id%now\, 
         \$19326_compbranch6504387_id%next\, 
         \$19326_compbranch6504387_id%now\, \$19203_compare6444358_id%next\, 
         \$19203_compare6444358_id%now\, \$18437_loop666_id%next\, 
         \$18437_loop666_id%now\, \$19097_modulo6684356_id%next\, 
         \$19097_modulo6684356_id%now\, \$18945_modulo6684356_id%next\, 
         \$18945_modulo6684356_id%now\, \$19066_modulo6684357_id%next\, 
         \$19066_modulo6684357_id%now\, 
         \$19601_copy_root_in_ram6634352_id%next\, 
         \$19601_copy_root_in_ram6634352_id%now\, 
         \$19370_compare6444359_id%next\, \$19370_compare6444359_id%now\, 
         \$18522_loop665_id%next\, \$18522_loop665_id%now\, 
         \$19171_compare6444358_id%next\, \$19171_compare6444358_id%now\, 
         \$18936_modulo6684349_id%next\, \$18936_modulo6684349_id%now\, 
         \$19144_modulo6684349_id%next\, \$19144_modulo6684349_id%now\, 
         \$19190_binop_compare6454380_id%next\, 
         \$19190_binop_compare6454380_id%now\, 
         \$18939_binop_int6434363_id%next\, \$18939_binop_int6434363_id%now\, 
         \$18797_branch_if648_id%next\, \$18797_branch_if648_id%now\, 
         \$18971_modulo6684357_id%next\, \$18971_modulo6684357_id%now\, 
         \$19262_forever6704385_id%next\, \$19262_forever6704385_id%now\, 
         \$19330_compare6444359_id%next\, \$19330_compare6444359_id%now\, 
         \$19497_loop666_id%next\, \$19497_loop666_id%now\, 
         \$18794_apply638_id%next\, \$18794_apply638_id%now\, 
         \$19238_w6514383_id%next\, \$19238_w6514383_id%now\, 
         \$18526_aux664_id%next\, \$18526_aux664_id%now\, 
         \$19532_forever6704350_id%next\, \$19532_forever6704350_id%now\, 
         \$19043_modulo6684349_id%next\, \$19043_modulo6684349_id%now\, 
         \$18990_modulo6684357_id%next\, \$18990_modulo6684357_id%now\, 
         \$18799_w1656_id%next\, \$18799_w1656_id%now\, 
         \$19333_compbranch6504388_id%next\, 
         \$19333_compbranch6504388_id%now\, \$19320_forever6704386_id%next\, 
         \$19320_forever6704386_id%now\, \$18958_binop_int6434364_id%next\, 
         \$18958_binop_int6434364_id%now\, \$18907_modulo6684356_id%next\, 
         \$18907_modulo6684356_id%now\, \$18790_loop666_id%next\, 
         \$18790_loop666_id%now\, \$18964_modulo6684356_id%next\, 
         \$18964_modulo6684356_id%now\, \$18977_binop_int6434365_id%next\, 
         \$18977_binop_int6434365_id%now\, \$18996_binop_int6434366_id%next\, 
         \$18996_binop_int6434366_id%now\, \$19012_modulo6684349_id%next\, 
         \$19012_modulo6684349_id%now\, \$19088_modulo6684349_id%next\, 
         \$19088_modulo6684349_id%now\, \$19021_modulo6684356_id%next\, 
         \$19021_modulo6684356_id%now\, \$18993_modulo6684349_id%next\, 
         \$18993_modulo6684349_id%now\, \$19384_compare6444359_id%next\, 
         \$19384_compare6444359_id%now\, \$19179_compare6444358_id%next\, 
         \$19179_compare6444358_id%now\, \$19078_modulo6684356_id%next\, 
         \$19078_modulo6684356_id%now\, \$19211_compare6444358_id%next\, 
         \$19211_compare6444358_id%now\, 
         \$18571_copy_root_in_ram6634345_id%next\, 
         \$18571_copy_root_in_ram6634345_id%now\, 
         \$18796_make_block_n646_id%next\, \$18796_make_block_n646_id%now\, 
         \$18521_loop666_id%next\, \$18521_loop666_id%now\, 
         \$19387_compbranch6504394_id%next\, 
         \$19387_compbranch6504394_id%now\, 
         \$19535_copy_root_in_ram6634354_id%next\, 
         \$19535_copy_root_in_ram6634354_id%now\, 
         \$19391_compare6444359_id%next\, \$19391_compare6444359_id%now\, 
         \$19337_compare6444359_id%next\, \$19337_compare6444359_id%now\, 
         \$18613_copy_root_in_ram6634346_id%next\, 
         \$18613_copy_root_in_ram6634346_id%now\, \$19495_loop665_id%next\, 
         \$19495_loop665_id%now\, \$19157_forever6704375_id%next\, 
         \$19157_forever6704375_id%now\, \$19062_modulo6684349_id%next\, 
         \$19062_modulo6684349_id%now\, \$18466_loop666_id%next\, 
         \$18466_loop666_id%now\, \$18926_modulo6684356_id%next\, 
         \$18926_modulo6684356_id%now\, \$19187_compare6444358_id%next\, 
         \$19187_compare6444358_id%now\, \$19163_forever6704376_id%next\, 
         \$19163_forever6704376_id%now\, \$19015_binop_int6434367_id%next\, 
         \$19015_binop_int6434367_id%now\, 
         \$19811_copy_root_in_ram6634341_id%next\, 
         \$19811_copy_root_in_ram6634341_id%now\, 
         \$18793_make_block579_id%next\, \$18793_make_block579_id%now\, 
         \$19129_modulo6684357_id%next\, \$19129_modulo6684357_id%now\, 
         \$19589_copy_root_in_ram6634353_id%next\, 
         \$19589_copy_root_in_ram6634353_id%now\, 
         \$19040_modulo6684356_id%next\, \$19040_modulo6684356_id%now\, 
         \$19104_modulo6684357_id%next\, \$19104_modulo6684357_id%now\, 
         \$19499_aux664_id%next\, \$19499_aux664_id%now\, 
         \$19132_modulo6684349_id%next\, \$19132_modulo6684349_id%now\, 
         \$19380_compbranch6504393_id%next\, 
         \$19380_compbranch6504393_id%now\, \$18933_modulo6684357_id%next\, 
         \$18933_modulo6684357_id%now\, \$18974_modulo6684349_id%next\, 
         \$18974_modulo6684349_id%now\, \$19779_loop666_id%next\, 
         \$19779_loop666_id%now\, \$19069_modulo6684349_id%next\, 
         \$19069_modulo6684349_id%now\, \$18910_modulo6684349_id%next\, 
         \$18910_modulo6684349_id%now\ : value(0 to 11) := (others => '0');
  signal \$19008_r%next\, \$19008_r%now\, \$18943_res%next\, 
         \$18943_res%now\, \$18917_modulo6684349_result%next\, 
         \$18917_modulo6684349_result%now\, \$18981_res%next\, 
         \$18981_res%now\, \$18929_modulo6684349_result%next\, 
         \$18929_modulo6684349_result%now\, 
         \$18910_modulo6684349_result%next\, 
         \$18910_modulo6684349_result%now\, 
         \$19059_modulo6684356_result%next\, 
         \$19059_modulo6684356_result%now\, \$19058_r%next\, \$19058_r%now\, 
         \$19050_modulo6684349_result%next\, 
         \$19050_modulo6684349_result%now\, \$v5783%next\, \$v5783%now\, 
         \$18989_r%next\, \$18989_r%now\, \$18964_modulo6684356_result%next\, 
         \$18964_modulo6684356_result%now\, \$18932_r%next\, \$18932_r%now\, 
         \$19132_modulo6684349_result%next\, 
         \$19132_modulo6684349_result%now\, \$19215_argument1%next\, 
         \$19215_argument1%now\, \$19129_modulo6684357_result%next\, 
         \$19129_modulo6684357_result%now\, \$19065_r%next\, \$19065_r%now\, 
         \$18970_r%next\, \$18970_r%now\, \$19151_modulo6684349_result%next\, 
         \$19151_modulo6684349_result%now\, \$19039_r%next\, \$19039_r%now\, 
         \$19002_modulo6684356_result%next\, 
         \$19002_modulo6684356_result%now\, \$19340_argument2%next\, 
         \$19340_argument2%now\, \$19069_modulo6684349_result%next\, 
         \$19069_modulo6684349_result%now\, \$19121_r%next\, \$19121_r%now\, 
         \$19107_modulo6684349_result%next\, 
         \$19107_modulo6684349_result%now\, \$19095_res%next\, 
         \$19095_res%now\, \$18983_modulo6684356_result%next\, 
         \$18983_modulo6684356_result%now\, \$19103_r%next\, \$19103_r%now\, 
         \$19000_res%next\, \$19000_res%now\, 
         \$18936_modulo6684349_result%next\, 
         \$18936_modulo6684349_result%now\, \$v5770%next\, \$v5770%now\, 
         \$19148_modulo6684357_result%next\, 
         \$19148_modulo6684357_result%now\, \$19433%next\, \$19433%now\, 
         \$19100_modulo6684349_result%next\, 
         \$19100_modulo6684349_result%now\, 
         \$19005_modulo6684349_result%next\, 
         \$19005_modulo6684349_result%now\, \$18951_r%next\, \$18951_r%now\, 
         \$18963_r%next\, \$18963_r%now\, \$18914_modulo6684357_result%next\, 
         \$18914_modulo6684357_result%now\, 
         \$18971_modulo6684357_result%next\, 
         \$18971_modulo6684357_result%now\, \$v5753%next\, \$v5753%now\, 
         \$18967_modulo6684349_result%next\, 
         \$18967_modulo6684349_result%now\, 
         \$19021_modulo6684356_result%next\, 
         \$19021_modulo6684356_result%now\, \$19147_r%next\, \$19147_r%now\, 
         \$19084_r%next\, \$19084_r%now\, \$19266%next\, \$19266%now\, 
         \$18986_modulo6684349_result%next\, 
         \$18986_modulo6684349_result%now\, 
         \$19078_modulo6684356_result%next\, 
         \$19078_modulo6684356_result%now\, 
         \$18907_modulo6684356_result%next\, 
         \$18907_modulo6684356_result%now\, 
         \$19012_modulo6684349_result%next\, 
         \$19012_modulo6684349_result%now\, 
         \$19009_modulo6684357_result%next\, 
         \$19009_modulo6684357_result%now\, 
         \$19047_modulo6684357_result%next\, 
         \$19047_modulo6684357_result%now\, 
         \$18955_modulo6684349_result%next\, 
         \$18955_modulo6684349_result%now\, \$19027_r%next\, \$19027_r%now\, 
         \$19031_modulo6684349_result%next\, 
         \$19031_modulo6684349_result%now\, 
         \$19144_modulo6684349_result%next\, 
         \$19144_modulo6684349_result%now\, 
         \$19125_modulo6684349_result%next\, 
         \$19125_modulo6684349_result%now\, \$v5799%next\, \$v5799%now\, 
         \$19046_r%next\, \$19046_r%now\, \$18944_r%next\, \$18944_r%now\, 
         \$19104_modulo6684357_result%next\, 
         \$19104_modulo6684357_result%now\, 
         \$19141_modulo6684356_result%next\, 
         \$19141_modulo6684356_result%now\, \$19120_res%next\, 
         \$19120_res%now\, \$19040_modulo6684356_result%next\, 
         \$19040_modulo6684356_result%now\, \$18925_r%next\, \$18925_r%now\, 
         \$19038_res%next\, \$19038_res%now\, \$19057_res%next\, 
         \$19057_res%now\, \$18926_modulo6684356_result%next\, 
         \$18926_modulo6684356_result%now\, \$19441_arg%next\, 
         \$19441_arg%now\, \$19077_r%next\, \$19077_r%now\, \$19020_r%next\, 
         \$19020_r%now\, \$19097_modulo6684356_result%next\, 
         \$19097_modulo6684356_result%now\, \$19128_r%next\, \$19128_r%now\, 
         \$19019_res%next\, \$19019_res%now\, \$18905_res%next\, 
         \$18905_res%now\, \$18948_modulo6684349_result%next\, 
         \$18948_modulo6684349_result%now\, \$18982_r%next\, \$18982_r%now\, 
         \$19096_r%next\, \$19096_r%now\, \$18816%next\, \$18816%now\, 
         \$18933_modulo6684357_result%next\, 
         \$18933_modulo6684357_result%now\, \$18962_res%next\, 
         \$18962_res%now\, \$19408_argument3%next\, \$19408_argument3%now\, 
         \$18913_r%next\, \$18913_r%now\, \$18906_r%next\, \$18906_r%now\, 
         \$19139_res%next\, \$19139_res%now\, 
         \$18952_modulo6684357_result%next\, 
         \$18952_modulo6684357_result%now\, 
         \$19081_modulo6684349_result%next\, 
         \$19081_modulo6684349_result%now\, 
         \$19088_modulo6684349_result%next\, 
         \$19088_modulo6684349_result%now\, 
         \$19062_modulo6684349_result%next\, 
         \$19062_modulo6684349_result%now\, \$19076_res%next\, 
         \$19076_res%now\, \$18974_modulo6684349_result%next\, 
         \$18974_modulo6684349_result%now\, \$v5760%next\, \$v5760%now\, 
         \$19066_modulo6684357_result%next\, 
         \$19066_modulo6684357_result%now\, \$19427%next\, \$19427%now\, 
         \$19043_modulo6684349_result%next\, 
         \$19043_modulo6684349_result%now\, 
         \$18990_modulo6684357_result%next\, 
         \$18990_modulo6684357_result%now\, 
         \$19028_modulo6684357_result%next\, 
         \$19028_modulo6684357_result%now\, \$18924_res%next\, 
         \$18924_res%now\, \$19122_modulo6684356_result%next\, 
         \$19122_modulo6684356_result%now\, \$19001_r%next\, \$19001_r%now\, 
         \$19140_r%next\, \$19140_r%now\, \$19024_modulo6684349_result%next\, 
         \$19024_modulo6684349_result%now\, 
         \$18993_modulo6684349_result%next\, 
         \$18993_modulo6684349_result%now\, 
         \$19085_modulo6684357_result%next\, 
         \$19085_modulo6684357_result%now\, 
         \$18945_modulo6684356_result%next\, 
         \$18945_modulo6684356_result%now\ : value(0 to 30) := (others => '0');
  signal \$18795_offsetclosure_n639_arg%next\, 
         \$18795_offsetclosure_n639_arg%now\ : value(0 to 137) := (others => '0');
  signal \$18793_make_block579_arg%next\, \$18793_make_block579_arg%now\ : value(0 to 103) := (others => '0');
  signal \$18469_make_block579_arg%next\, \$18469_make_block579_arg%now\, 
         \result4963%next\, \result4963%now\, \result4607%next\, 
         \result4607%now\, \result4434%next\, \result4434%now\, 
         \$18440_make_block579_arg%next\, \$18440_make_block579_arg%now\ : value(0 to 127) := (others => '0');
  signal \$code_lock%next\, \$code_lock%now\, \$global_end_lock%next\, 
         \$global_end_lock%now\, \$ram_lock%next\, \$ram_lock%now\, 
         \$19630%next\, \$19630%now\, \$19699%next\, \$19699%now\, 
         \$18862%next\, \$18862%now\, \$19669%next\, \$19669%now\, 
         \$v5535%next\, \$v5535%now\, \$v5667%next\, \$v5667%now\, 
         \$v4731%next\, \$v4731%now\, \$v5230%next\, \$v5230%now\, 
         \$v5350%next\, \$v5350%now\, \$19567%next\, \$19567%now\, 
         \$v5438%next\, \$v5438%now\, \$19805%next\, \$19805%now\, 
         \$19252_forever6704384_arg%next\, \$19252_forever6704384_arg%now\, 
         \$19729%next\, \$19729%now\, \$19573%next\, \$19573%now\, 
         \$19862%next\, \$19862%now\, \$v4404%next\, \$v4404%now\, 
         \$v5520%next\, \$v5520%now\, \$v5661%next\, \$v5661%now\, 
         \$v4896%next\, \$v4896%now\, \$19370_compare6444359_result%next\, 
         \$19370_compare6444359_result%now\, \$19692%next\, \$19692%now\, 
         \$19555%next\, \$19555%now\, \$19513%next\, \$19513%now\, 
         \$18543%next\, \$18543%now\, \$v4622%next\, \$v4622%now\, 
         \$v5590%next\, \$v5590%now\, \$v4869%next\, \$v4869%now\, 
         \$v4625%next\, \$v4625%now\, \$18568%next\, \$18568%now\, 
         \$19593%next\, \$19593%now\, \$v4848%next\, \$v4848%now\, 
         \$v4971%next\, \$v4971%now\, \$19782%next\, \$19782%now\, 
         \$18491%next\, \$18491%now\, \$19171_compare6444358_result%next\, 
         \$19171_compare6444358_result%now\, \$18588%next\, \$18588%now\, 
         \$18496%next\, \$18496%now\, \$19693%next\, \$19693%now\, 
         \$18656%next\, \$18656%now\, \$19516%next\, \$19516%now\, 
         \$v5240%next\, \$v5240%now\, \$19224%next\, \$19224%now\, 
         \$19221%next\, \$19221%now\, \$19802%next\, \$19802%now\, 
         \$19633%next\, \$19633%now\, \$v4933%next\, \$v4933%now\, 
         \$19635%next\, \$19635%now\, \$18477%next\, \$18477%now\, 
         \$19262_forever6704385_arg%next\, \$19262_forever6704385_arg%now\, 
         \$v5480%next\, \$v5480%now\, \$19792%next\, \$19792%now\, 
         \$v5917%next\, \$v5917%now\, \$19627%next\, \$19627%now\, 
         \$v5093%next\, \$v5093%now\, \$v5207%next\, \$v5207%now\, 
         \$v4508%next\, \$v4508%now\, \$19808_forever6704342_arg%next\, 
         \$19808_forever6704342_arg%now\, \$18811%next\, \$18811%now\, 
         \$v4808%next\, \$v4808%now\, \$v5399%next\, \$v5399%now\, 
         \$18499%next\, \$18499%now\, \$19223%next\, \$19223%now\, 
         \$19277%next\, \$19277%now\, \$v5779%next\, \$v5779%now\, 
         \$v5503%next\, \$v5503%now\, \$v4439%next\, \$v4439%now\, 
         \$v5056%next\, \$v5056%now\, \$19484%next\, \$19484%now\, 
         \$18634%next\, \$18634%now\, \$v5417%next\, \$v5417%now\, 
         \$19940%next\, \$19940%now\, \$18719%next\, \$18719%now\, 
         \$18692%next\, \$18692%now\, \$v5075%next\, \$v5075%now\, 
         \$v5553%next\, \$v5553%now\, \$18847%next\, \$18847%now\, 
         \$v5165%next\, \$v5165%now\, \$18833%next\, \$18833%now\, 
         \$19429%next\, \$19429%now\, \$19733%next\, \$19733%now\, 
         \$v5215%next\, \$v5215%now\, \$v5423%next\, \$v5423%now\, 
         \$18530%next\, \$18530%now\, \$v5087%next\, \$v5087%now\, 
         \$18700%next\, \$18700%now\, \$18675%next\, \$18675%now\, 
         \$v5554%next\, \$v5554%now\, \$v5016%next\, \$v5016%now\, 
         \$v5798%next\, \$v5798%now\, \$v5914%next\, \$v5914%now\, 
         \$v5886%next\, \$v5886%now\, \$v5864%next\, \$v5864%now\, 
         \$v5786%next\, \$v5786%now\, \$19690%next\, \$19690%now\, 
         \$v5854%next\, \$v5854%now\, \$18503%next\, \$18503%now\, 
         \$v4580%next\, \$v4580%now\, \$v4723%next\, \$v4723%now\, 
         \$19568%next\, \$19568%now\, \$v5834%next\, \$v5834%now\, 
         \$19708%next\, \$19708%now\, \$18774%next\, \$18774%now\, 
         \$19481%next\, \$19481%now\, \$19831%next\, \$19831%now\, 
         \$v5048%next\, \$v5048%now\, \$v5746%next\, \$v5746%now\, 
         \$v5583%next\, \$v5583%now\, \$19502%next\, \$19502%now\, 
         \$18804%next\, \$18804%now\, \$v5006%next\, \$v5006%now\, 
         \$19195_compare6444358_result%next\, 
         \$19195_compare6444358_result%now\, \$19606%next\, \$19606%now\, 
         \$19652%next\, \$19652%now\, \$19696%next\, \$19696%now\, 
         \$v4522%next\, \$v4522%now\, \$v5504%next\, \$v5504%now\, 
         \$19511%next\, \$19511%now\, \$v5842%next\, \$v5842%now\, 
         \$19654%next\, \$19654%now\, \$v4962%next\, \$v4962%now\, 
         \$v5338%next\, \$v5338%now\, \$19283%next\, \$19283%now\, 
         \$18528%next\, \$18528%now\, \$v4764%next\, \$v4764%now\, 
         \$18501%next\, \$18501%now\, \$18486%next\, \$18486%now\, 
         \$v5706%next\, \$v5706%now\, \$v5435%next\, \$v5435%now\, 
         \$v5901%next\, \$v5901%now\, \$18471%next\, \$18471%now\, 
         \$19691%next\, \$19691%now\, \$18481%next\, \$18481%now\, 
         \$19369_b%next\, \$19369_b%now\, \$19424%next\, \$19424%now\, 
         \$v5877%next\, \$v5877%now\, \$v5680%next\, \$v5680%now\, 
         \$18594%next\, \$18594%now\, \$v5241%next\, \$v5241%now\, 
         \$v4778%next\, \$v4778%now\, \$19289%next\, \$19289%now\, 
         \$18592%next\, \$18592%now\, \$v5600%next\, \$v5600%now\, 
         \$19330_compare6444359_result%next\, 
         \$19330_compare6444359_result%now\, 
         \$18556_forever6704344_arg%next\, \$18556_forever6704344_arg%now\, 
         \$19841%next\, \$19841%now\, \$19712%next\, \$19712%now\, 
         \$v5676%next\, \$v5676%now\, \$18710%next\, \$18710%now\, 
         \$v4452%next\, \$v4452%now\, \$18665%next\, \$18665%now\, 
         \$19730%next\, \$19730%now\, \$v4956%next\, \$v4956%now\, 
         \$18513%next\, \$18513%now\, \$19935%next\, \$19935%now\, 
         \$18722%next\, \$18722%now\, \$v4644%next\, \$v4644%now\, 
         \$v5521%next\, \$v5521%now\, \$v4875%next\, \$v4875%now\, 
         \$19520%next\, \$19520%now\, \$v4788%next\, \$v4788%now\, 
         \$19655%next\, \$19655%now\, \$v4427%next\, \$v4427%now\, 
         \$v5740%next\, \$v5740%now\, \$18773%next\, \$18773%now\, 
         \$18641%next\, \$18641%now\, \$19577%next\, \$19577%now\, 
         \$v5372%next\, \$v5372%now\, \$19943%next\, \$19943%now\, 
         \$19946%next\, \$19946%now\, \$v4463%next\, \$v4463%now\, 
         \$v4914%next\, \$v4914%now\, \$19911%next\, \$19911%now\, 
         \$18538%next\, \$18538%now\, \$19562%next\, \$19562%now\, 
         \$18628%next\, \$18628%now\, \$18772%next\, \$18772%now\, 
         \$18548%next\, \$18548%now\, \$19318%next\, \$19318%now\, 
         \$19473%next\, \$19473%now\, \$19270%next\, \$19270%now\, 
         \$19323%next\, \$19323%now\, \$v5501%next\, \$v5501%now\, 
         \$v4657%next\, \$v4657%now\, \$19640%next\, \$19640%now\, 
         \$18466_loop666_result%next\, \$18466_loop666_result%now\, 
         \$v4999%next\, \$v4999%now\, \$v5581%next\, \$v5581%now\, 
         \$v4643%next\, \$v4643%now\, \$18860%next\, \$18860%now\, 
         \$v5375%next\, \$v5375%now\, \$18490%next\, \$18490%now\, 
         \$19756%next\, \$19756%now\, \$v5219%next\, \$v5219%now\, 
         \$v5155%next\, \$v5155%now\, \$19645%next\, \$19645%now\, 
         \$18547%next\, \$18547%now\, \$19411%next\, \$19411%now\, 
         \$19618%next\, \$19618%now\, \$19219%next\, \$19219%now\, 
         \$19545%next\, \$19545%now\, \$18587%next\, \$18587%now\, 
         \$19624%next\, \$19624%now\, \$v4446%next\, \$v4446%now\, 
         \$19404_b%next\, \$19404_b%now\, \$v5718%next\, \$v5718%now\, 
         \$19472%next\, \$19472%now\, \$v4686%next\, \$v4686%now\, 
         \$v4968%next\, \$v4968%now\, \$v5022%next\, \$v5022%now\, 
         \$v5820%next\, \$v5820%now\, \$18878%next\, \$18878%now\, 
         \$18445_x%next\, \$18445_x%now\, \$v5474%next\, \$v5474%now\, 
         \$v5381%next\, \$v5381%now\, \$v4747%next\, \$v4747%now\, 
         \$v5575%next\, \$v5575%now\, \$19426%next\, \$19426%now\, 
         \$18437_loop666_result%next\, \$18437_loop666_result%now\, 
         \$18597%next\, \$18597%now\, \$18693%next\, \$18693%now\, 
         \$v5106%next\, \$v5106%now\, \$v5792%next\, \$v5792%now\, 
         \$v4635%next\, \$v4635%now\, \$18771%next\, \$18771%now\, 
         \$18616%next\, \$18616%now\, \$18713%next\, \$18713%now\, 
         \$19225%next\, \$19225%now\, \$18611%next\, \$18611%now\, 
         \$18636%next\, \$18636%now\, \$19938%next\, \$19938%now\, 
         \$18617%next\, \$18617%now\, \$18672%next\, \$18672%now\, 
         \$v5887%next\, \$v5887%now\, \$19830%next\, \$19830%now\, 
         \$v4987%next\, \$v4987%now\, \$19847%next\, \$19847%now\, 
         \$v4785%next\, \$v4785%now\, \$19612%next\, \$19612%now\, 
         \$18586%next\, \$18586%now\, \$19111%next\, \$19111%now\, 
         \$19898%next\, \$19898%now\, \$19900%next\, \$19900%now\, 
         \$19869%next\, \$19869%now\, \$19510%next\, \$19510%now\, 
         \$v5805%next\, \$v5805%now\, \$19604%next\, \$19604%now\, 
         \$19791%next\, \$19791%now\, \$18743%next\, \$18743%now\, 
         \$19912%next\, \$19912%now\, \$v4755%next\, \$v4755%now\, 
         \$18690%next\, \$18690%now\, \rdy4964%next\, \rdy4964%now\, 
         \$v4411%next\, \$v4411%now\, \$19337_compare6444359_result%next\, 
         \$19337_compare6444359_result%now\, \$v5302%next\, \$v5302%now\, 
         \$v5229%next\, \$v5229%now\, \$18593%next\, \$18593%now\, 
         \$19632%next\, \$19632%now\, \$v5493%next\, \$v5493%now\, 
         \$v4526%next\, \$v4526%now\, \$18686%next\, \$18686%now\, 
         \$18671%next\, \$18671%now\, \$v5110%next\, \$v5110%now\, 
         \$18736%next\, \$18736%now\, \$19705%next\, \$19705%now\, 
         \$19459%next\, \$19459%now\, \$18633%next\, \$18633%now\, 
         \$v5593%next\, \$v5593%now\, \$19405_compare6444359_result%next\, 
         \$19405_compare6444359_result%now\, \$v5808%next\, \$v5808%now\, 
         \$19711%next\, \$19711%now\, \$19556%next\, \$19556%now\, 
         \$19457%next\, \$19457%now\, \$19670%next\, \$19670%now\, 
         \$19738%next\, \$19738%now\, \$18814%next\, \$18814%now\, 
         \$v5408%next\, \$v5408%now\, \$v5918%next\, \$v5918%now\, 
         \$19899%next\, \$19899%now\, \$v5500%next\, \$v5500%now\, 
         \$19622%next\, \$19622%now\, \$v5712%next\, \$v5712%now\, 
         \$v4737%next\, \$v4737%now\, \$v4707%next\, \$v4707%now\, 
         \$v5177%next\, \$v5177%now\, \$19695%next\, \$19695%now\, 
         \$v5841%next\, \$v5841%now\, \$19846%next\, \$19846%now\, 
         \$18691%next\, \$18691%now\, \$18803%next\, \$18803%now\, 
         \$19857%next\, \$19857%now\, \$v4332%next\, \$v4332%now\, 
         \$v5736%next\, \$v5736%now\, \$19365%next\, \$19365%now\, 
         \$v4432%next\, \$v4432%now\, \$18585%next\, \$18585%now\, 
         \$19634%next\, \$19634%now\, \$v5483%next\, \$v5483%now\, 
         \$19919%next\, \$19919%now\, \$19587%next\, \$19587%now\, 
         \$v4600%next\, \$v4600%now\, \$18589%next\, \$18589%now\, 
         \$v4890%next\, \$v4890%now\, \$v5531%next\, \$v5531%now\, 
         \$v5211%next\, \$v5211%now\, \$v5591%next\, \$v5591%now\, 
         \$v4991%next\, \$v4991%now\, \$18861%next\, \$18861%now\, 
         \$v5218%next\, \$v5218%now\, \$v4553%next\, \$v4553%now\, 
         \$18596%next\, \$18596%now\, \$v4905%next\, \$v4905%now\, 
         \$v5362%next\, \$v5362%now\, \$19113_forever6704372_arg%next\, 
         \$19113_forever6704372_arg%now\, \$v5848%next\, \$v5848%now\, 
         \$18753%next\, \$18753%now\, \$v5510%next\, \$v5510%now\, 
         \$19822%next\, \$19822%now\, \$18678%next\, \$18678%now\, 
         \$v5111%next\, \$v5111%now\, \$v5851%next\, \$v5851%now\, 
         \$18658%next\, \$18658%now\, \$18716%next\, \$18716%now\, 
         \$v5626%next\, \$v5626%now\, \$v5341%next\, \$v5341%now\, 
         \$18839%next\, \$18839%now\, \$19461%next\, \$19461%now\, 
         \$v5192%next\, \$v5192%now\, \$v5114%next\, \$v5114%now\, 
         \$v5756%next\, \$v5756%now\, \$v5572%next\, \$v5572%now\, 
         \$v4333%next\, \$v4333%now\, \$v5030%next\, \$v5030%now\, 
         \$v5880%next\, \$v5880%now\, \$v4670%next\, \$v4670%now\, 
         \$v5045%next\, \$v5045%now\, \$v5332%next\, \$v5332%now\, 
         \$18871%next\, \$18871%now\, \$19663%next\, \$19663%now\, 
         \$19160%next\, \$19160%now\, \$19178_res%next\, \$19178_res%now\, 
         \$v5562%next\, \$v5562%now\, \result4572%next\, \result4572%now\, 
         \$v4720%next\, \$v4720%now\, \$19258%next\, \$19258%now\, 
         \$v4487%next\, \$v4487%now\, \$v4536%next\, \$v4536%now\, 
         \$19757%next\, \$19757%now\, \$v4557%next\, \$v4557%now\, 
         \$18800%next\, \$18800%now\, \$18874%next\, \$18874%now\, 
         \$19305%next\, \$19305%now\, \$v4459%next\, \$v4459%now\, 
         \$18757%next\, \$18757%now\, \$19552%next\, \$19552%now\, 
         \$18720%next\, \$18720%now\, \$18609%next\, \$18609%now\, 
         \rdy4435%next\, \rdy4435%now\, \$19278%next\, \$19278%now\, 
         \$v5561%next\, \$v5561%now\, \$19428%next\, \$19428%now\, 
         \$v5695%next\, \$v5695%now\, \$19762%next\, \$19762%now\, 
         \$v5919%next\, \$v5919%now\, \$v4774%next\, \$v4774%now\, 
         \$19598%next\, \$19598%now\, \$18621%next\, \$18621%now\, 
         \$v4505%next\, \$v4505%now\, \$v5495%next\, \$v5495%now\, 
         \$v4478%next\, \$v4478%now\, \$v5782%next\, \$v5782%now\, 
         \$v5181%next\, \$v5181%now\, \$19767%next\, \$19767%now\, 
         \$v5459%next\, \$v5459%now\, \$19284%next\, \$19284%now\, 
         \$19494_loop666_result%next\, \$19494_loop666_result%now\, 
         \$v5585%next\, \$v5585%now\, \$19247%next\, \$19247%now\, 
         \$19524%next\, \$19524%now\, \$v5444%next\, \$v5444%now\, 
         \$18579%next\, \$18579%now\, \$18493%next\, \$18493%now\, 
         \$v5773%next\, \$v5773%now\, \$18544%next\, \$18544%now\, 
         \$v5602%next\, \$v5602%now\, \$v5387%next\, \$v5387%now\, 
         \$19576%next\, \$19576%now\, \$v5890%next\, \$v5890%now\, 
         \$18827%next\, \$18827%now\, \$v5126%next\, \$v5126%now\, 
         \$19271%next\, \$19271%now\, \$v4771%next\, \$v4771%now\, 
         \$v4981%next\, \$v4981%now\, \$v5894%next\, \$v5894%now\, 
         \$19753%next\, \$19753%now\, \$18607%next\, \$18607%now\, 
         \$v4488%next\, \$v4488%now\, \$v4758%next\, \$v4758%now\, 
         \$v5863%next\, \$v5863%now\, \$v4884%next\, \$v4884%now\, 
         \$19285%next\, \$19285%now\, \$19747%next\, \$19747%now\, 
         \$v4824%next\, \$v4824%now\, \$v4466%next\, \$v4466%now\, 
         \$19945%next\, \$19945%now\, \$v4795%next\, \$v4795%now\, 
         \$v4881%next\, \$v4881%now\, \$v5566%next\, \$v5566%now\, 
         \$19261%next\, \$19261%now\, \$18758%next\, \$18758%now\, 
         \$19621%next\, \$19621%now\, \$19286%next\, \$19286%now\, 
         \$v4857%next\, \$v4857%now\, \$18536%next\, \$18536%now\, 
         \$19497_loop666_result%next\, \$19497_loop666_result%now\, 
         \$v5556%next\, \$v5556%now\, \$19529_forever6704351_arg%next\, 
         \$19529_forever6704351_arg%now\, \$v5543%next\, \$v5543%now\, 
         \$18812%next\, \$18812%now\, \$19889%next\, \$19889%now\, 
         \$v5630%next\, \$v5630%now\, \$v5679%next\, \$v5679%now\, 
         \$v5051%next\, \$v5051%now\, \$v4597%next\, \$v4597%now\, 
         \$19893%next\, \$19893%now\, \$19580%next\, \$19580%now\, 
         \$19470%next\, \$19470%now\, \$19460%next\, \$19460%now\, 
         \$v4953%next\, \$v4953%now\, \$v5353%next\, \$v5353%now\, 
         \$19475%next\, \$19475%now\, \$19722%next\, \$19722%now\, 
         \$19341%next\, \$19341%now\, \$v5396%next\, \$v5396%now\, 
         \$v4716%next\, \$v4716%now\, \$18640%next\, \$18640%now\, 
         \$v4836%next\, \$v4836%now\, \$19605%next\, \$19605%now\, 
         \$18899%next\, \$18899%now\, \$v4902%next\, \$v4902%now\, 
         \$19941%next\, \$19941%now\, \$v4809%next\, \$v4809%now\, 
         \$19768%next\, \$19768%now\, \$19795%next\, \$19795%now\, 
         \$19749%next\, \$19749%now\, \$v5079%next\, \$v5079%now\, 
         \$18574%next\, \$18574%now\, \$19668%next\, \$19668%now\, 
         \$v5494%next\, \$v5494%now\, \$v5368%next\, \$v5368%now\, 
         \$19302%next\, \$19302%now\, \$v4917%next\, \$v4917%now\, 
         \$v5802%next\, \$v5802%now\, \$v4827%next\, \$v4827%now\, 
         \$19860%next\, \$19860%now\, \$v5099%next\, \$v5099%now\, 
         \$19864%next\, \$19864%now\, \$v4719%next\, \$v4719%now\, 
         \$19921%next\, \$19921%now\, \$v5670%next\, \$v5670%now\, 
         \$v5606%next\, \$v5606%now\, \$19876%next\, \$19876%now\, 
         \$v5251%next\, \$v5251%now\, \$v5689%next\, \$v5689%now\, 
         \$18714%next\, \$18714%now\, \$v5296%next\, \$v5296%now\, 
         \$19677%next\, \$19677%now\, \$v5039%next\, \$v5039%now\, 
         \$18735%next\, \$18735%now\, \$v4423%next\, \$v4423%now\, 
         \$19697%next\, \$19697%now\, \$19917%next\, \$19917%now\, 
         \$v5709%next\, \$v5709%now\, \$19586%next\, \$19586%now\, 
         \$18701%next\, \$18701%now\, \$19820%next\, \$19820%now\, 
         \$v4654%next\, \$v4654%now\, \$v5084%next\, \$v5084%now\, 
         \$18489%next\, \$18489%now\, \$18550%next\, \$18550%now\, 
         \$18777%next\, \$18777%now\, \$19719%next\, \$19719%now\, 
         \$19915%next\, \$19915%now\, \$v4782%next\, \$v4782%now\, 
         \$v5222%next\, \$v5222%now\, \$v5034%next\, \$v5034%now\, 
         \$v5185%next\, \$v5185%now\, \$v5000%next\, \$v5000%now\, 
         \$19833%next\, \$19833%now\, \$19646%next\, \$19646%now\, 
         \$v5867%next\, \$v5867%now\, \$v5505%next\, \$v5505%now\, 
         \$19799%next\, \$19799%now\, \$18715%next\, \$18715%now\, 
         \$18808%next\, \$18808%now\, \$18651%next\, \$18651%now\, 
         \$18780%next\, \$18780%now\, \$v5724%next\, \$v5724%now\, 
         \$19202_res%next\, \$19202_res%now\, 
         \$19398_compare6444359_result%next\, 
         \$19398_compare6444359_result%now\, \$18748%next\, \$18748%now\, 
         \$19592%next\, \$19592%now\, \$18786%next\, \$18786%now\, 
         \$v5525%next\, \$v5525%now\, \$v5293%next\, \$v5293%now\, 
         \$19927%next\, \$19927%now\, \$18595%next\, \$18595%now\, 
         \$18674%next\, \$18674%now\, \$v4960%next\, \$v4960%now\, 
         \$v5023%next\, \$v5023%now\, \$v5584%next\, \$v5584%now\, 
         \$v5356%next\, \$v5356%now\, \$v5909%next\, \$v5909%now\, 
         \$19456%next\, \$19456%now\, \$18497%next\, \$18497%now\, 
         \$18756%next\, \$18756%now\, \$v5411%next\, \$v5411%now\, 
         \$v5347%next\, \$v5347%now\, \$v4492%next\, \$v4492%now\, 
         \$19316%next\, \$19316%now\, \$v4514%next\, \$v4514%now\, 
         \$18676%next\, \$18676%now\, \$19615%next\, \$19615%now\, 
         \$19942%next\, \$19942%now\, \$19584%next\, \$19584%now\, 
         \$19383_b%next\, \$19383_b%now\, \$v5876%next\, \$v5876%now\, 
         \$v5652%next\, \$v5652%now\, \$v5491%next\, \$v5491%now\, 
         \$19345%next\, \$19345%now\, \$v5544%next\, \$v5544%now\, 
         \$18752%next\, \$18752%now\, \$19539%next\, \$19539%now\, 
         \$19242%next\, \$19242%now\, \$19807%next\, \$19807%now\, 
         \$19951%next\, \$19951%now\, \$v4689%next\, \$v4689%now\, 
         \$18515%next\, \$18515%now\, \$v5131%next\, \$v5131%now\, 
         \$19853%next\, \$19853%now\, \$v5605%next\, \$v5605%now\, 
         \$19260%next\, \$19260%now\, \$v5845%next\, \$v5845%now\, 
         \$v5814%next\, \$v5814%now\, \$v5502%next\, \$v5502%now\, 
         \$18516%next\, \$18516%now\, \$19879%next\, \$19879%now\, 
         \$v5441%next\, \$v5441%now\, \$18886%next\, \$18886%now\, 
         \$19585%next\, \$19585%now\, \$19451%next\, \$19451%now\, 
         \$19617%next\, \$19617%now\, \$v5540%next\, \$v5540%now\, 
         \$v5314%next\, \$v5314%now\, \$19642%next\, \$19642%now\, 
         \$v5432%next\, \$v5432%now\, \$v4813%next\, \$v4813%now\, 
         \$v5102%next\, \$v5102%now\, \$v4984%next\, \$v4984%now\, 
         \$18781%next\, \$18781%now\, \$v5107%next\, \$v5107%now\, 
         \$v4675%next\, \$v4675%now\, \$v5477%next\, \$v5477%now\, 
         \$v4496%next\, \$v4496%now\, \$18897%next\, \$18897%now\, 
         \$18702%next\, \$18702%now\, \$19649%next\, \$19649%now\, 
         \$19414%next\, \$19414%now\, \$v5743%next\, \$v5743%now\, 
         \$v4911%next\, \$v4911%now\, \$18654%next\, \$18654%now\, 
         \$19233%next\, \$19233%now\, \$19755%next\, \$19755%now\, 
         \$18487%next\, \$18487%now\, \$v4751%next\, \$v4751%now\, 
         \$v5560%next\, \$v5560%now\, \$19856%next\, \$19856%now\, 
         \$v5524%next\, \$v5524%now\, \$v4746%next\, \$v4746%now\, 
         \$v4791%next\, \$v4791%now\, \$v4833%next\, \$v4833%now\, 
         \$19500%next\, \$19500%now\, \$19351%next\, \$19351%now\, 
         \$19665%next\, \$19665%now\, \$19355%next\, \$19355%now\, 
         \$19293%next\, \$19293%now\, \$19425%next\, \$19425%now\, 
         \$18724%next\, \$18724%now\, \$19769%next\, \$19769%now\, 
         \$19700%next\, \$19700%now\, \$19834%next\, \$19834%now\, 
         \$v5335%next\, \$v5335%now\, \$18564%next\, \$18564%now\, 
         \$v4562%next\, \$v4562%now\, \$18498%next\, \$18498%now\, 
         \$18666%next\, \$18666%now\, \$v4539%next\, \$v4539%now\, 
         \$v4605%next\, \$v4605%now\, \$v4449%next\, \$v4449%now\, 
         \$18562%next\, \$18562%now\, \$19154%next\, \$19154%now\, 
         \$18639%next\, \$18639%now\, \$v5141%next\, \$v5141%now\, 
         \$v4606%next\, \$v4606%now\, \$19563%next\, \$19563%now\, 
         \$v5359%next\, \$v5359%now\, \$v5096%next\, \$v5096%now\, 
         \$v4337%next\, \$v4337%now\, \$19566%next\, \$19566%now\, 
         \$19214%next\, \$19214%now\, \$v4558%next\, \$v4558%now\, 
         \$19766%next\, \$19766%now\, \$18673%next\, \$18673%now\, 
         \$v5260%next\, \$v5260%now\, \$v4532%next\, \$v4532%now\, 
         \$v4339%next\, \$v4339%now\, \$19892%next\, \$19892%now\, 
         \$18642%next\, \$18642%now\, \$v5275%next\, \$v5275%now\, 
         \$v5254%next\, \$v5254%now\, \$v4754%next\, \$v4754%now\, 
         \$19872%next\, \$19872%now\, \$v4972%next\, \$v4972%now\, 
         \$v5138%next\, \$v5138%now\, \$v5188%next\, \$v5188%now\, 
         \$v5622%next\, \$v5622%now\, \$v5405%next\, \$v5405%now\, 
         \$19678%next\, \$19678%now\, \$19110%next\, \$19110%now\, 
         \$19315%next\, \$19315%now\, \$18508%next\, \$18508%now\, 
         \$v4640%next\, \$v4640%now\, \$v4455%next\, \$v4455%now\, 
         \$19832%next\, \$19832%now\, \$19521%next\, \$19521%now\, 
         \$19594%next\, \$19594%now\, \$v5596%next\, \$v5596%now\, 
         \$19329_b%next\, \$19329_b%now\, \$19636%next\, \$19636%now\, 
         \$18464_rdy%next\, \$18464_rdy%now\, \$19779_loop666_result%next\, 
         \$19779_loop666_result%now\, \$v5305%next\, \$v5305%now\, 
         \$v4937%next\, \$v4937%now\, \$18679%next\, \$18679%now\, 
         \$18663%next\, \$18663%now\, \$19868%next\, \$19868%now\, 
         \$18500%next\, \$18500%now\, \$v5664%next\, \$v5664%now\, 
         \$v4821%next\, \$v4821%now\, \$19638%next\, \$19638%now\, 
         \$v4540%next\, \$v4540%now\, \$19870%next\, \$19870%now\, 
         \$19519%next\, \$19519%now\, \$v4713%next\, \$v4713%now\, 
         \$v4775%next\, \$v4775%now\, \$19743%next\, \$19743%now\, 
         \$v4750%next\, \$v4750%now\, \$v4818%next\, \$v4818%now\, 
         \$19660%next\, \$19660%now\, \$19806%next\, \$19806%now\, 
         \$19561%next\, \$19561%now\, \$v4796%next\, \$v4796%now\, 
         \$19877%next\, \$19877%now\, \$19882%next\, \$19882%now\, 
         \$v5727%next\, \$v5727%now\, \$19772%next\, \$19772%now\, 
         \$19268%next\, \$19268%now\, \$v4940%next\, \$v4940%now\, 
         \$v4700%next\, \$v4700%now\, \$19532_forever6704350_arg%next\, 
         \$19532_forever6704350_arg%now\, \$19843%next\, \$19843%now\, 
         \$v5492%next\, \$v5492%now\, \$19728%next\, \$19728%now\, 
         \rdy4608%next\, \rdy4608%now\, \$18687%next\, \$18687%now\, 
         \$v4327%next\, \$v4327%now\, \$v5066%next\, \$v5066%now\, 
         \$19878%next\, \$19878%now\, \rdy4573%next\, \rdy4573%now\, 
         \$18660%next\, \$18660%now\, \$18669%next\, \$18669%now\, 
         \$19449%next\, \$19449%now\, \$19731%next\, \$19731%now\, 
         \$v5453%next\, \$v5453%now\, \$v4556%next\, \$v4556%now\, 
         \$v4887%next\, \$v4887%now\, \$18629%next\, \$18629%now\, 
         \$19922%next\, \$19922%now\, \$v5072%next\, \$v5072%now\, 
         \$18478%next\, \$18478%now\, \$v5897%next\, \$v5897%now\, 
         \$v5563%next\, \$v5563%now\, \$19391_compare6444359_result%next\, 
         \$19391_compare6444359_result%now\, \$18898%next\, \$18898%now\, 
         \$19572%next\, \$19572%now\, \$v5384%next\, \$v5384%now\, 
         \$19937%next\, \$19937%now\, \$v4615%next\, \$v4615%now\, 
         \$v5571%next\, \$v5571%now\, \$18492%next\, \$18492%now\, 
         \$19156%next\, \$19156%now\, \$19161%next\, \$19161%now\, 
         \$v4581%next\, \$v4581%now\, \$v5198%next\, \$v5198%now\, 
         \$18476%next\, \$18476%now\, \$19503%next\, \$19503%now\, 
         \$v5696%next\, \$v5696%now\, \$19815%next\, \$19815%now\, 
         \$19310%next\, \$19310%now\, \$18470%next\, \$18470%now\, 
         \$19639%next\, \$19639%now\, \$19875%next\, \$19875%now\, 
         \$v5471%next\, \$v5471%now\, \$18618%next\, \$18618%now\, 
         \$18732%next\, \$18732%now\, \$19725%next\, \$19725%now\, 
         \$v4471%next\, \$v4471%now\, \$19512%next\, \$19512%now\, 
         \$v5811%next\, \$v5811%now\, \$v5552%next\, \$v5552%now\, 
         \$v5915%next\, \$v5915%now\, \$v4335%next\, \$v4335%now\, 
         \$v5184%next\, \$v5184%now\, \$18649%next\, \$18649%now\, 
         \$v4683%next\, \$v4683%now\, \$18567%next\, \$18567%now\, 
         \$v4639%next\, \$v4639%now\, \$v4802%next\, \$v4802%now\, 
         \$18531%next\, \$18531%now\, \$v4502%next\, \$v4502%now\, 
         \$18546%next\, \$18546%now\, \$19619%next\, \$19619%now\, 
         \$19709%next\, \$19709%now\, \$19336_b%next\, \$19336_b%now\, 
         \$v4957%next\, \$v4957%now\, \$v4632%next\, \$v4632%now\, 
         \$v5233%next\, \$v5233%now\, \$18845%next\, \$18845%now\, 
         \$v4679%next\, \$v4679%now\, \$v4839%next\, \$v4839%now\, 
         \$v4529%next\, \$v4529%now\, \$v5168%next\, \$v5168%now\, 
         \$19543%next\, \$19543%now\, \$19701%next\, \$19701%now\, 
         \$v5365%next\, \$v5365%now\, \$18603%next\, \$18603%now\, 
         \$19932%next\, \$19932%now\, \$v5134%next\, \$v5134%now\, 
         \$18473%next\, \$18473%now\, \$19259%next\, \$19259%now\, 
         \$18695%next\, \$18695%now\, \$v4593%next\, \$v4593%now\, 
         \$19667%next\, \$19667%now\, \$v4519%next\, \$v4519%now\, 
         \$18622%next\, \$18622%now\, \$19804%next\, \$19804%now\, 
         \$18790_loop666_result%next\, \$18790_loop666_result%now\, 
         \$19211_compare6444358_result%next\, 
         \$19211_compare6444358_result%now\, \$v4678%next\, \$v4678%now\, 
         \$v4667%next\, \$v4667%now\, \$18813%next\, \$18813%now\, 
         \$v5042%next\, \$v5042%now\, \rdy4400%next\, \rdy4400%now\, 
         \$19783%next\, \$19783%now\, \$v5522%next\, \$v5522%now\, 
         \$19774%next\, \$19774%now\, \$v5055%next\, \$v5055%now\, 
         \$v4428%next\, \$v4428%now\, \$v5257%next\, \$v5257%now\, 
         \$18659%next\, \$18659%now\, \$v5490%next\, \$v5490%now\, 
         \$18869%next\, \$18869%now\, \$18880%next\, \$18880%now\, 
         \$19944%next\, \$19944%now\, \$18810%next\, \$18810%now\, 
         \$v4920%next\, \$v4920%now\, \$v4978%next\, \$v4978%now\, 
         \$19571%next\, \$19571%now\, \$v5429%next\, \$v5429%now\, 
         \$19837%next\, \$19837%now\, \$18444%next\, \$18444%now\, 
         \$v5574%next\, \$v5574%now\, \$v4812%next\, \$v4812%now\, 
         \$v4636%next\, \$v4636%now\, \$v4779%next\, \$v4779%now\, 
         \$v4546%next\, \$v4546%now\, \$v5281%next\, \$v5281%now\, 
         \$v4330%next\, \$v4330%now\, \$18891%next\, \$18891%now\, 
         \$v4647%next\, \$v4647%now\, \$v4866%next\, \$v4866%now\, 
         \$18806%next\, \$18806%now\, \$18825%next\, \$18825%now\, 
         \$v5036%next\, \$v5036%now\, \$v4996%next\, \$v4996%now\, 
         \$v5026%next\, \$v5026%now\, \$18657%next\, \$18657%now\, 
         \$v5059%next\, \$v5059%now\, \$v5206%next\, \$v5206%now\, 
         \$18461%next\, \$18461%now\, \$19748%next\, \$19748%now\, 
         \$19384_compare6444359_result%next\, 
         \$19384_compare6444359_result%now\, \$v4338%next\, \$v4338%now\, 
         \$19581%next\, \$19581%now\, \$19597%next\, \$19597%now\, 
         \$18539%next\, \$18539%now\, \$v5299%next\, \$v5299%now\, 
         \$v5536%next\, \$v5536%now\, \$19842%next\, \$19842%now\, 
         \$v5673%next\, \$v5673%now\, \$19793%next\, \$19793%now\, 
         \$18648%next\, \$18648%now\, \$18527%next\, \$18527%now\, 
         \$19325%next\, \$19325%now\, \$19859%next\, \$19859%now\, 
         \$19276%next\, \$19276%now\, \$v5658%next\, \$v5658%now\, 
         \$18551%next\, \$18551%now\, \$18495%next\, \$18495%now\, 
         \$19650%next\, \$19650%now\, \$19939%next\, \$19939%now\, 
         \$v4587%next\, \$v4587%now\, \$18661%next\, \$18661%now\, 
         \$19155%next\, \$19155%now\, \$18647%next\, \$18647%now\, 
         \$v5769%next\, \$v5769%now\, \$v4424%next\, \$v4424%now\, 
         \$19773%next\, \$19773%now\, \$v5482%next\, \$v5482%now\, 
         \$19886%next\, \$19886%now\, \$v5576%next\, \$v5576%now\, 
         \$19625%next\, \$19625%now\, \$v4420%next\, \$v4420%now\, 
         \$19487%next\, \$19487%now\, \$v4671%next\, \$v4671%now\, 
         \$18511%next\, \$18511%now\, \$19317%next\, \$19317%now\, 
         \$18608%next\, \$18608%now\, \$v5311%next\, \$v5311%now\, 
         \$19914%next\, \$19914%now\, \$v5462%next\, \$v5462%now\, 
         \$v5390%next\, \$v5390%now\, \$v4704%next\, \$v4704%now\, 
         \$18721%next\, \$18721%now\, \$19471%next\, \$19471%now\, 
         \$19626%next\, \$19626%now\, \$v5550%next\, \$v5550%now\, 
         \$v5003%next\, \$v5003%now\, \$19798%next\, \$19798%now\, 
         \$v5447%next\, \$v5447%now\, \$v4407%next\, \$v4407%now\, 
         \$18688%next\, \$18688%now\, \$19376_b%next\, \$19376_b%now\, 
         \$18505%next\, \$18505%now\, \$v5523%next\, \$v5523%now\, 
         \$19304%next\, \$19304%now\, \$v4408%next\, \$v4408%now\, 
         \$v5090%next\, \$v5090%now\, \$v5402%next\, \$v5402%now\, 
         \$18747%next\, \$18747%now\, \$18514%next\, \$18514%now\, 
         \$v5169%next\, \$v5169%now\, \$19210_res%next\, \$19210_res%now\, 
         \$19913%next\, \$19913%now\, \$19801%next\, \$19801%now\, 
         \$v5637%next\, \$v5637%now\, \$v4518%next\, \$v4518%now\, 
         \$v4612%next\, \$v4612%now\, \$18580%next\, \$18580%now\, 
         \$18475%next\, \$18475%now\, \$19295%next\, \$19295%now\, 
         \$v5817%next\, \$v5817%now\, \$19540%next\, \$19540%now\, 
         \$v5083%next\, \$v5083%now\, \$18575%next\, \$18575%now\, 
         \$18540%next\, \$18540%now\, \$18604%next\, \$18604%now\, 
         \$v5468%next\, \$v5468%now\, \$18549%next\, \$18549%now\, 
         \$19901%next\, \$19901%now\, \$18521_loop666_result%next\, 
         \$18521_loop666_result%now\, \$v4651%next\, \$v4651%now\, 
         \$19888%next\, \$19888%now\, \$v4619%next\, \$v4619%now\, 
         \$19570%next\, \$19570%now\, \$v5344%next\, \$v5344%now\, 
         \$19582%next\, \$19582%now\, \$v4696%next\, \$v4696%now\, 
         \$18782%next\, \$18782%now\, \$19517%next\, \$19517%now\, 
         \$19557%next\, \$19557%now\, \$18851%next\, \$18851%now\, 
         \$19871%next\, \$19871%now\, \$19884%next\, \$19884%now\, 
         \$v4872%next\, \$v4872%now\, \$19836%next\, \$19836%now\, 
         \$19275%next\, \$19275%now\, \$v4571%next\, \$v4571%now\, 
         \$19255%next\, \$19255%now\, \$19538%next\, \$19538%now\, 
         \$19243%next\, \$19243%now\, \$19544%next\, \$19544%now\, 
         \$19522%next\, \$19522%now\, \$v5103%next\, \$v5103%now\, 
         \$19179_compare6444358_result%next\, 
         \$19179_compare6444358_result%now\, \$v4549%next\, \$v4549%now\, 
         \$19920%next\, \$19920%now\, \$v5199%next\, \$v5199%now\, 
         \$v5649%next\, \$v5649%now\, \$19891%next\, \$19891%now\, 
         \$v4442%next\, \$v4442%now\, \$v5189%next\, \$v5189%now\, 
         \$v4767%next\, \$v4767%now\, \$19546%next\, \$19546%now\, 
         \$v5266%next\, \$v5266%now\, \$19249%next\, \$19249%now\, 
         \$18677%next\, \$18677%now\, \$19883%next\, \$19883%now\, 
         \$v4458%next\, \$v4458%now\, \$v4666%next\, \$v4666%now\, 
         \$18472%next\, \$18472%now\, \rdy4929%next\, \rdy4929%now\, 
         \$19734%next\, \$19734%now\, \$18826%next\, \$18826%now\, 
         \$19785%next\, \$19785%now\, \$18537%next\, \$18537%now\, 
         \$19771%next\, \$19771%now\, \$19710%next\, \$19710%now\, 
         \$v4431%next\, \$v4431%now\, \$19637%next\, \$19637%now\, 
         \$19664%next\, \$19664%now\, \$v5570%next\, \$v5570%now\, 
         \$19203_compare6444358_result%next\, 
         \$19203_compare6444358_result%now\, 
         \$19377_compare6444359_result%next\, 
         \$19377_compare6444359_result%now\, \$v5007%next\, \$v5007%now\, 
         \$v5730%next\, \$v5730%now\, \$v4899%next\, \$v4899%now\, 
         \$v5147%next\, \$v5147%now\, \$v4495%next\, \$v4495%now\, 
         \$v5135%next\, \$v5135%now\, \$18863%next\, \$18863%now\, 
         \$19794%next\, \$19794%now\, \$18749%next\, \$18749%now\, 
         \$18849%next\, \$18849%now\, \$v4860%next\, \$v4860%now\, 
         \$v4799%next\, \$v4799%now\, \$v5618%next\, \$v5618%now\, 
         \$v5763%next\, \$v5763%now\, \$v5080%next\, \$v5080%now\, 
         \$18494%next\, \$18494%now\, \$v5174%next\, \$v5174%now\, 
         \$19821%next\, \$19821%now\, \$v5393%next\, \$v5393%now\, 
         \$v5063%next\, \$v5063%now\, \$v5225%next\, \$v5225%now\, 
         \$19320_forever6704386_arg%next\, \$19320_forever6704386_arg%now\, 
         \$v5573%next\, \$v5573%now\, \$v5496%next\, \$v5496%now\, 
         \$19873%next\, \$19873%now\, \$19509%next\, \$19509%now\, 
         \$18770%next\, \$18770%now\, \$19564%next\, \$19564%now\, 
         \$19923%next\, \$19923%now\, \$19523%next\, \$19523%now\, 
         \$v5010%next\, \$v5010%now\, \$18681%next\, \$18681%now\, 
         \$v5450%next\, \$v5450%now\, \$v5789%next\, \$v5789%now\, 
         \$19352%next\, \$19352%now\, \$v4724%next\, \$v4724%now\, 
         \$19849%next\, \$19849%now\, \$18718%next\, \$18718%now\, 
         \$18750%next\, \$18750%now\, \$v5161%next\, \$v5161%now\, 
         \$v5456%next\, \$v5456%now\, \$v5031%next\, \$v5031%now\, 
         \$v5545%next\, \$v5545%now\, \$18552%next\, \$18552%now\, 
         \$18601%next\, \$18601%now\, \$19675%next\, \$19675%now\, 
         \$v4570%next\, \$v4570%now\, \$v5511%next\, \$v5511%now\, 
         \$v5601%next\, \$v5601%now\, \$19936%next\, \$19936%now\, 
         \$v5329%next\, \$v5329%now\, \$v4893%next\, \$v4893%now\, 
         \$v5580%next\, \$v5580%now\, \$v4851%next\, \$v4851%now\, 
         \$19162%next\, \$19162%now\, \$18798_w652_result%next\, 
         \$18798_w652_result%now\, \$18799_w1656_result%next\, 
         \$18799_w1656_result%now\, \$19826%next\, \$19826%now\, 
         \$19750%next\, \$19750%now\, \$18734%next\, \$18734%now\, 
         \$v4475%next\, \$v4475%now\, \$19671%next\, \$19671%now\, 
         \$v5893%next\, \$v5893%now\, \$18479%next\, \$18479%now\, 
         \$v5534%next\, \$v5534%now\, \$v4975%next\, \$v4975%now\, 
         \$19686%next\, \$19686%now\, \$19610%next\, \$19610%now\, 
         \$19666%next\, \$19666%now\, \$v4792%next\, \$v4792%now\, 
         \$19616%next\, \$19616%now\, \$v4484%next\, \$v4484%now\, 
         \$18465%next\, \$18465%now\, \$v5512%next\, \$v5512%now\, 
         \$v5317%next\, \$v5317%now\, \$v4943%next\, \$v4943%now\, 
         \$19588%next\, \$19588%now\, \$19835%next\, \$19835%now\, 
         \$v4923%next\, \$v4923%now\, \$v5565%next\, \$v5565%now\, 
         \$v5202%next\, \$v5202%now\, \$v5795%next\, \$v5795%now\, 
         \$18755%next\, \$18755%now\, \$19694%next\, \$19694%now\, 
         \$19631%next\, \$19631%now\, \$18689%next\, \$18689%now\, 
         \$19186_res%next\, \$19186_res%now\, \$v5269%next\, \$v5269%now\, 
         \$19551%next\, \$19551%now\, \$19303%next\, \$19303%now\, 
         \$18612%next\, \$18612%now\, \$v5272%next\, \$v5272%now\, 
         \$18779%next\, \$18779%now\, \$19858%next\, \$19858%now\, 
         \$19908%next\, \$19908%now\, \$v5144%next\, \$v5144%now\, 
         \$19724%next\, \$19724%now\, \$v5546%next\, \$v5546%now\, 
         \$18459%next\, \$18459%now\, \$18725%next\, \$18725%now\, 
         \$19786%next\, \$19786%now\, \$19861%next\, \$19861%now\, 
         \$19483%next\, \$19483%now\, \$19647%next\, \$19647%now\, 
         \$19438%next\, \$19438%now\, \$v5170%next\, \$v5170%now\, 
         \$v5148%next\, \$v5148%now\, \$18717%next\, \$18717%now\, 
         \$v4462%next\, \$v4462%now\, \$19676%next\, \$19676%now\, 
         \$v5737%next\, \$v5737%now\, \$18829%next\, \$18829%now\, 
         \$v5123%next\, \$v5123%now\, \$18831%next\, \$18831%now\, 
         \$v4699%next\, \$v4699%now\, \$v5595%next\, \$v5595%now\, 
         \$v5130%next\, \$v5130%now\, \$19651%next\, \$19651%now\, 
         \$v5290%next\, \$v5290%now\, \$v5203%next\, \$v5203%now\, 
         \$18746%next\, \$18746%now\, \$18488%next\, \$18488%now\, 
         \$19746%next\, \$19746%now\, \$v4863%next\, \$v4863%now\, 
         \$19565%next\, \$19565%now\, \$v5542%next\, \$v5542%now\, 
         \$19313%next\, \$19313%now\, \$v5426%next\, \$v5426%now\, 
         \$19855%next\, \$19855%now\, \$v5180%next\, \$v5180%now\, 
         \$v5516%next\, \$v5516%now\, \$19550%next\, \$19550%now\, 
         \$v5485%next\, \$v5485%now\, \$19397_b%next\, \$19397_b%now\, 
         \$18754%next\, \$18754%now\, \$18643%next\, \$18643%now\, 
         \$18553_forever6704348_arg%next\, \$18553_forever6704348_arg%now\, 
         \$v5533%next\, \$v5533%now\, \$19852%next\, \$19852%now\, 
         \$v5237%next\, \$v5237%now\, \$v4414%next\, \$v4414%now\, 
         \$v5860%next\, \$v5860%now\, \$18684%next\, \$18684%now\, 
         \$v5069%next\, \$v5069%now\, \$18610%next\, \$18610%now\, 
         \$v5027%next\, \$v5027%now\, \$v5614%next\, \$v5614%now\, 
         \$v5835%next\, \$v5835%now\, \$v5263%next\, \$v5263%now\, 
         \$18570%next\, \$18570%now\, \$v5420%next\, \$v5420%now\, 
         \$v4543%next\, \$v4543%now\, \$v5247%next\, \$v5247%now\, 
         \$v4328%next\, \$v4328%now\, \$19918%next\, \$19918%now\, 
         \$18460%next\, \$18460%now\, \$19825%next\, \$19825%now\, 
         \$19754%next\, \$19754%now\, \$18623%next\, \$18623%now\, 
         \$v5465%next\, \$v5465%now\, \$19867%next\, \$19867%now\, 
         \$19157_forever6704375_arg%next\, \$19157_forever6704375_arg%now\, 
         \$19751%next\, \$19751%now\, \$18680%next\, \$18680%now\, 
         \$18699%next\, \$18699%now\, \$v4842%next\, \$v4842%now\, 
         \$19726%next\, \$19726%now\, \$v5555%next\, \$v5555%now\, 
         \$v5883%next\, \$v5883%now\, \$18591%next\, \$18591%now\, 
         \$v5564%next\, \$v5564%now\, \$19474%next\, \$19474%now\, 
         \$19488%next\, \$19488%now\, \$v5905%next\, \$v5905%now\, 
         \$v5284%next\, \$v5284%now\, \$v5278%next\, \$v5278%now\, 
         \$19280%next\, \$19280%now\, \$19558%next\, \$19558%now\, 
         \$18605%next\, \$18605%now\, \$19578%next\, \$19578%now\, 
         \$19526_forever6704355_arg%next\, \$19526_forever6704355_arg%now\, 
         \$19599%next\, \$19599%now\, \$18864%next\, \$18864%now\, 
         \$v4433%next\, \$v4433%now\, \$v5195%next\, \$v5195%now\, 
         \$19679%next\, \$19679%now\, \$v4878%next\, \$v4878%now\, 
         \$19359%next\, \$19359%now\, \$18767%next\, \$18767%now\, 
         \$19698%next\, \$19698%now\, \$v4584%next\, \$v4584%now\, 
         \$19413%next\, \$19413%now\, \$19662%next\, \$19662%now\, 
         \$18510%next\, \$18510%now\, \$19727%next\, \$19727%now\, 
         \$19390_b%next\, \$19390_b%now\, \$v4660%next\, \$v4660%now\, 
         \$18733%next\, \$18733%now\, \$18484%next\, \$18484%now\, 
         \$v4601%next\, \$v4601%now\, \$v4995%next\, \$v4995%now\, 
         \$v5308%next\, \$v5308%now\, \$v4740%next\, \$v4740%now\, 
         \$v5831%next\, \$v5831%now\, \$v5164%next\, \$v5164%now\, 
         \$v5823%next\, \$v5823%now\, \$19569%next\, \$19569%now\, 
         \$19269%next\, \$19269%now\, \$v5514%next\, \$v5514%now\, 
         \$v4805%next\, \$v4805%now\, \$19887%next\, \$19887%now\, 
         \$v5127%next\, \$v5127%now\, \$v4680%next\, \$v4680%now\, 
         \$19814%next\, \$19814%now\, \$19232%next\, \$19232%now\, 
         \$19848%next\, \$19848%now\, \$v4988%next\, \$v4988%now\, 
         \$19854%next\, \$19854%now\, \$v5120%next\, \$v5120%now\, 
         \$19648%next\, \$19648%now\, \$19251%next\, \$19251%now\, 
         \$18635%next\, \$18635%now\, \$v4908%next\, \$v4908%now\, 
         \$18576%next\, \$18576%now\, \$v4695%next\, \$v4695%now\, 
         \$19897%next\, \$19897%now\, \$18645%next\, \$18645%now\, 
         \$18563%next\, \$18563%now\, \$v5250%next\, \$v5250%now\, 
         \$v4674%next\, \$v4674%now\, \$18644%next\, \$18644%now\, 
         \$v5530%next\, \$v5530%now\, \$19885%next\, \$19885%now\, 
         \$19600%next\, \$19600%now\, \$v5244%next\, \$v5244%now\, 
         \$18600%next\, \$18600%now\, \$18662%next\, \$18662%now\, 
         \$v5481%next\, \$v5481%now\, \$v5702%next\, \$v5702%now\, 
         \$v4992%next\, \$v4992%now\, \$18447%next\, \$18447%now\, 
         \$v4417%next\, \$v4417%now\, \$v4936%next\, \$v4936%now\, 
         \$18485%next\, \$18485%now\, \$18646%next\, \$18646%now\, 
         \$18664%next\, \$18664%now\, \$v4946%next\, \$v4946%now\, 
         \$v5052%next\, \$v5052%now\, \$19623%next\, \$19623%now\, 
         \$v5378%next\, \$v5378%now\, \$19187_compare6444358_result%next\, 
         \$19187_compare6444358_result%now\, \$v4552%next\, \$v4552%now\, 
         \$v5060%next\, \$v5060%now\, \$v5582%next\, \$v5582%now\, 
         \$v5603%next\, \$v5603%now\, \$18685%next\, \$18685%now\, 
         \$v5035%next\, \$v5035%now\, \$v4631%next\, \$v4631%now\, 
         \$v4845%next\, \$v4845%now\, \$19816%next\, \$19816%now\, 
         \$v4761%next\, \$v4761%now\, \$19248%next\, \$19248%now\, 
         \$v5604%next\, \$v5604%now\, \$18670%next\, \$18670%now\, 
         \$18590%next\, \$18590%now\, \$v4596%next\, \$v4596%now\, 
         \$v4728%next\, \$v4728%now\, \$18762%next\, \$18762%now\, 
         \$19314%next\, \$19314%now\, \$v5640%next\, \$v5640%now\, 
         \$v4481%next\, \$v4481%now\, \$18723%next\, \$18723%now\, 
         \$v5838%next\, \$v5838%now\, \$19583%next\, \$19583%now\, 
         \$v5828%next\, \$v5828%now\, \$19294%next\, \$19294%now\, 
         \$v5655%next\, \$v5655%now\, \$18458%next\, \$18458%now\, 
         \$18480%next\, \$18480%now\, \$19656%next\, \$19656%now\, 
         \$v4734%next\, \$v4734%now\, \$v4727%next\, \$v4727%now\, 
         \$v4491%next\, \$v4491%now\, \$v5210%next\, \$v5210%now\, 
         \$18815%next\, \$18815%now\, \$19609%next\, \$19609%now\, 
         \$19732%next\, \$19732%now\, \$19434%next\, \$19434%now\, 
         \$v4770%next\, \$v4770%now\, \$18502%next\, \$18502%now\, 
         \$19784%next\, \$19784%now\, \$19611%next\, \$19611%now\, 
         \$19482%next\, \$19482%now\, \$v5749%next\, \$v5749%now\, 
         \$v4569%next\, \$v4569%now\, \$v4523%next\, \$v4523%now\, 
         \$19829%next\, \$19829%now\, \$v4926%next\, \$v4926%now\, 
         \$v5506%next\, \$v5506%now\, \$18703%next\, \$18703%now\, 
         \$v4628%next\, \$v4628%now\, \$v4854%next\, \$v4854%now\, 
         \$v5686%next\, \$v5686%now\, \$19916%next\, \$19916%now\, 
         \$18529%next\, \$18529%now\, \$v4692%next\, \$v4692%now\, 
         \$18482%next\, \$18482%now\, \$v5857%next\, \$v5857%now\, 
         \$19486%next\, \$19486%now\, \$v4949%next\, \$v4949%now\, 
         \$19217%next\, \$19217%now\, \$19803%next\, \$19803%now\, 
         \$19620%next\, \$19620%now\, \$19657%next\, \$19657%now\, 
         \$v5683%next\, \$v5683%now\, \$v5610%next\, \$v5610%now\, 
         \$v4952%next\, \$v4952%now\, \$v5646%next\, \$v5646%now\, 
         \$19319%next\, \$19319%now\, \$v5515%next\, \$v5515%now\, 
         \$19112%next\, \$19112%now\, \$18805%next\, \$18805%now\, 
         \$18569%next\, \$18569%now\, \$18837%next\, \$18837%now\, 
         \$18650%next\, \$18650%now\, \$19504%next\, \$19504%now\, 
         \$18807%next\, \$18807%now\, \$v5019%next\, \$v5019%now\, 
         \$v5776%next\, \$v5776%now\, \$19489%next\, \$19489%now\, 
         \$19819%next\, \$19819%now\, \$19894%next\, \$19894%now\, 
         \$v4616%next\, \$v4616%now\, \$19752%next\, \$19752%now\, 
         \$v5766%next\, \$v5766%now\, \$v5234%next\, \$v5234%now\, 
         \$v5586%next\, \$v5586%now\, \$19458%next\, \$19458%now\, 
         \$v5721%next\, \$v5721%now\, \$v5212%next\, \$v5212%now\, 
         \$v5320%next\, \$v5320%now\, \$v5703%next\, \$v5703%now\, 
         \$19419%next\, \$19419%now\, \$v5759%next\, \$v5759%now\, 
         \$18694%next\, \$18694%now\, \$18778%next\, \$18778%now\, 
         \$19723%next\, \$19723%now\, \$v4472%next\, \$v4472%now\, 
         \$18524_loop666_result%next\, \$18524_loop666_result%now\, 
         \$v4590%next\, \$v4590%now\, \$v4511%next\, \$v4511%now\, 
         \$19890%next\, \$19890%now\, \$18865%next\, \$18865%now\, 
         \$v5752%next\, \$v5752%now\, \$18867%next\, \$18867%now\, 
         \$19445%next\, \$19445%now\, \$v5117%next\, \$v5117%now\, 
         \$v4830%next\, \$v4830%now\, \$v5594%next\, \$v5594%now\, 
         \$v5151%next\, \$v5151%now\, \$19653%next\, \$19653%now\, 
         \$18876%next\, \$18876%now\, \$v4443%next\, \$v4443%now\, 
         \$v5414%next\, \$v5414%now\, \$19661%next\, \$19661%now\, 
         \$v5733%next\, \$v5733%now\, \$v5369%next\, \$v5369%now\, 
         \$v5158%next\, \$v5158%now\, \$19641%next\, \$19641%now\, 
         \$18474%next\, \$18474%now\, \$v5692%next\, \$v5692%now\, 
         \$19672%next\, \$19672%now\, \$19947%next\, \$19947%now\, 
         \$19194_res%next\, \$19194_res%now\, \$v5592%next\, \$v5592%now\, 
         \$18655%next\, \$18655%now\, \$v5323%next\, \$v5323%now\, 
         \$v4515%next\, \$v4515%now\, \$18509%next\, \$18509%now\, 
         \$19525%next\, \$19525%now\, \$v5013%next\, \$v5013%now\, 
         \$18582%next\, \$18582%now\, \$v5226%next\, \$v5226%now\, 
         \$v5551%next\, \$v5551%now\, \$v4535%next\, \$v4535%now\, 
         \$18630%next\, \$18630%now\, \$19432%next\, \$19432%now\, 
         \$19827%next\, \$19827%now\, \$19863%next\, \$19863%now\, 
         \$19170_res%next\, \$19170_res%now\, \$v4814%next\, \$v4814%now\, 
         \$v4710%next\, \$v4710%now\, \$18483%next\, \$18483%now\, 
         \$v4703%next\, \$v4703%now\, \$v5152%next\, \$v5152%now\, 
         \$19501%next\, \$19501%now\, \$v5532%next\, \$v5532%now\, 
         \$v5076%next\, \$v5076%now\, \$18802%next\, \$18802%now\, 
         \$v4577%next\, \$v4577%now\, \$19689%next\, \$19689%now\, 
         \$19245%next\, \$19245%now\, \$18696%next\, \$18696%now\, 
         \$v4325%next\, \$v4325%now\, \$v4470%next\, \$v4470%now\, 
         \$18900%next\, \$18900%now\, \$v4467%next\, \$v4467%now\, 
         \$v5287%next\, \$v5287%now\, \$18581%next\, \$18581%now\, 
         \$v5634%next\, \$v5634%now\, \$19292%next\, \$19292%now\, 
         \$v5699%next\, \$v5699%now\, \$v4604%next\, \$v4604%now\, 
         \$19163_forever6704376_arg%next\, \$19163_forever6704376_arg%now\, 
         \$18776%next\, \$18776%now\, \$19758%next\, \$19758%now\, 
         \$19579%next\, \$19579%now\, \$18835%next\, \$18835%now\, 
         \$v4650%next\, \$v4650%now\, \$18624%next\, \$18624%now\, 
         \$19250%next\, \$19250%now\, \$v5643%next\, \$v5643%now\, 
         \$18504%next\, \$18504%now\, \$v5484%next\, \$v5484%now\, 
         \$v5326%next\, \$v5326%now\, \$v4499%next\, \$v4499%now\, 
         \$v4961%next\, \$v4961%now\, \$19828%next\, \$19828%now\, 
         \$v5715%next\, \$v5715%now\, \$19874%next\, \$19874%now\, 
         \$18775%next\, \$18775%now\, \$18801%next\, \$18801%now\, 
         \$18729%next\, \$18729%now\, \$v5513%next\, \$v5513%now\, 
         \$v5486%next\, \$v5486%now\, \$19272%next\, \$19272%now\, 
         \$18751%next\, \$18751%now\, \$18809%next\, \$18809%now\, 
         \$v5541%next\, \$v5541%now\, \$18602%next\, \$18602%now\, 
         \$v5913%next\, \$v5913%now\, \$v4663%next\, \$v4663%now\, 
         \$v5526%next\, \$v5526%now\, \$19299%next\, \$19299%now\, 
         \$v4743%next\, \$v4743%now\, \$18606%next\, \$18606%now\ : value(0 to 0) := (others => '0');
  signal \$18794_apply638_arg%next\, \$18794_apply638_arg%now\ : value(0 to 165) := (others => '0');
  signal \$18796_make_block_n646_arg%next\, \$18796_make_block_n646_arg%now\ : value(0 to 171) := (others => '0');
  signal \$19838_copy_root_in_ram6634340_arg%next\, 
         \$19838_copy_root_in_ram6634340_arg%now\, 
         \$18468_wait662_result%next\, \$18468_wait662_result%now\, 
         \$19547_copy_root_in_ram6634352_arg%next\, 
         \$19547_copy_root_in_ram6634352_arg%now\, 
         \$18625_copy_root_in_ram6634345_arg%next\, 
         \$18625_copy_root_in_ram6634345_arg%now\, 
         \$19589_copy_root_in_ram6634353_arg%next\, 
         \$19589_copy_root_in_ram6634353_arg%now\, \$18535%next\, 
         \$18535%now\, \$19416_w36574398_arg%next\, 
         \$19416_w36574398_arg%now\, \$18799_w1656_arg%next\, 
         \$18799_w1656_arg%now\, \$18613_copy_root_in_ram6634346_arg%next\, 
         \$18613_copy_root_in_ram6634346_arg%now\, \$19770%next\, 
         \$19770%now\, \$18439_wait662_result%next\, 
         \$18439_wait662_result%now\, \$19485%next\, \$19485%now\, 
         \$18559_copy_root_in_ram6634347_arg%next\, 
         \$18559_copy_root_in_ram6634347_arg%now\, 
         \$19811_copy_root_in_ram6634341_arg%next\, 
         \$19811_copy_root_in_ram6634341_arg%now\, 
         \$19601_copy_root_in_ram6634352_arg%next\, 
         \$19601_copy_root_in_ram6634352_arg%now\, 
         \$18792_wait662_result%next\, \$18792_wait662_result%now\, 
         \$19790%next\, \$19790%now\, 
         \$19535_copy_root_in_ram6634354_arg%next\, 
         \$19535_copy_root_in_ram6634354_arg%now\, 
         \$19361_fill6544390_arg%next\, \$19361_fill6544390_arg%now\, 
         \$18571_copy_root_in_ram6634345_arg%next\, 
         \$18571_copy_root_in_ram6634345_arg%now\, 
         \$19347_fill6534389_arg%next\, \$19347_fill6534389_arg%now\, 
         \$18512%next\, \$18512%now\, \$19508%next\, \$19508%now\ : value(0 to 79) := (others => '0');
  signal \$18519%next\, \$18519%now\, \$19493%next\, \$19493%now\, 
         \$19492%next\, \$19492%now\, \$18520%next\, \$18520%now\, 
         \$19778%next\, \$19778%now\, \$19777%next\, \$19777%now\ : value(0 to 128) := (others => '0');
  signal \$v5547%next\, \$v5547%now\, \$18761%next\, \$18761%now\, 
         \$18449%next\, \$18449%now\, \$18942_v%next\, \$18942_v%now\, 
         \$19229_v%next\, \$19229_v%now\, \$19575_hd%next\, \$19575_hd%now\, 
         \$v5517%next\, \$v5517%now\, \$19688_hd%next\, \$19688_hd%now\, 
         \$18887_v%next\, \$18887_v%now\, \$19541%next\, \$19541%now\, 
         \$19644_hd%next\, \$19644_hd%now\, \$19291_v%next\, \$19291_v%now\, 
         \$19881_hd%next\, \$19881_hd%now\, \$18712_hd%next\, 
         \$18712_hd%now\, \$18653_hd%next\, \$18653_hd%now\, \$18744_w%next\, 
         \$18744_w%now\, \$19469%next\, \$19469%now\, \$18923_v%next\, 
         \$18923_v%now\, \$18704%next\, \$18704%now\, \$19477_v%next\, 
         \$19477_v%now\, \$18853_hd%next\, \$18853_hd%now\, \$v5527%next\, 
         \$v5527%now\, \$19613_w%next\, \$19613_w%now\, \$19216_v%next\, 
         \$19216_v%now\, \$19353%next\, \$19353%now\, \$19560_hd%next\, 
         \$19560_hd%now\, \$v5587%next\, \$v5587%now\, \$18866_v%next\, 
         \$18866_v%now\, \$19356%next\, \$19356%now\, \$19236_v%next\, 
         \$19236_v%now\, \$18879_v%next\, \$18879_v%now\, \$19056_v%next\, 
         \$19056_v%now\, \$v5567%next\, \$v5567%now\, \$19306_v%next\, 
         \$19306_v%now\, \$18819_v%next\, \$18819_v%now\, \$v5631%next\, 
         \$v5631%now\, \$18850%next\, \$18850%now\, \$19763%next\, 
         \$19763%now\, \$18868_v%next\, \$18868_v%now\, \$19437%next\, 
         \$19437%now\, \$18892_v%next\, \$18892_v%now\, \$18894_v%next\, 
         \$18894_v%now\, \$19745_hd%next\, \$19745_hd%now\, \$19687_w%next\, 
         \$19687_w%now\, \$19244_v%next\, \$19244_v%now\, \$18728%next\, 
         \$18728%now\, \$v5615%next\, \$v5615%now\, \$19680%next\, 
         \$19680%now\, \$18652_w%next\, \$18652_w%now\, \$18823_v%next\, 
         \$18823_v%now\, \$v5871%next\, \$v5871%now\, \$18836_v%next\, 
         \$18836_v%now\, \$19629_hd%next\, \$19629_hd%now\, \$18818_v%next\, 
         \$18818_v%now\, \$v5868%next\, \$v5868%now\, \$19037_v%next\, 
         \$19037_v%now\, \$19237_v%next\, \$19237_v%now\, \$19574_w%next\, 
         \$19574_w%now\, \$19476_v%next\, \$19476_v%now\, \$18840_v%next\, 
         \$18840_v%now\, \$18885_v%next\, \$18885_v%now\, \$18883_v%next\, 
         \$18883_v%now\, \$19193_v%next\, \$19193_v%now\, \$19744_w%next\, 
         \$19744_w%now\, \$19933_w%next\, \$19933_w%now\, \$19607%next\, 
         \$19607%now\, \$18890_v%next\, \$18890_v%now\, \$18817_v%next\, 
         \$18817_v%now\, \$18872_v%next\, \$18872_v%now\, \$19298_v%next\, 
         \$19298_v%now\, \$19287_v%next\, \$19287_v%now\, \$v5623%next\, 
         \$v5623%now\, \$18882_v%next\, \$18882_v%now\, \$18708%next\, 
         \$18708%now\, \$v5627%next\, \$v5627%now\, \$18785%next\, 
         \$18785%now\, \$18870_v%next\, \$18870_v%now\, \$19228_v%next\, 
         \$19228_v%now\, \$19823_w%next\, \$19823_w%now\, \$18741%next\, 
         \$18741%now\, \$19138_v%next\, \$19138_v%now\, \$18768_w%next\, 
         \$18768_w%now\, \$18842%next\, \$18842%now\, \$19297_v%next\, 
         \$19297_v%now\, \$19865_w%next\, \$19865_w%now\, \$18844%next\, 
         \$18844%now\, \$19241_v%next\, \$19241_v%now\, \$v5497%next\, 
         \$v5497%now\, \$18820_v%next\, \$18820_v%now\, \$19658_w%next\, 
         \$19658_w%now\, \$18838_v%next\, \$18838_v%now\, \$19737%next\, 
         \$19737%now\, \$18446_dur%next\, \$18446_dur%now\, \$18737%next\, 
         \$18737%now\, \$18896_v%next\, \$18896_v%now\, \$v5597%next\, 
         \$v5597%now\, \$19950%next\, \$19950%now\, \$18904_v%next\, 
         \$18904_v%now\, \$18682_w%next\, \$18682_w%now\, \$19684%next\, 
         \$19684%now\, \$19614_hd%next\, \$19614_hd%now\, \$19926%next\, 
         \$19926%now\, \$v5825%next\, \$v5825%now\, \$18583_w%next\, 
         \$18583_w%now\, \$19257_v%next\, \$19257_v%now\, \$19282_v%next\, 
         \$19282_v%now\, \$18889_v%next\, \$18889_v%now\, \$19226%next\, 
         \$19226%now\, \$19301_v%next\, \$19301_v%now\, \$18631%next\, 
         \$18631%now\, \$18895_v%next\, \$18895_v%now\, \$19741%next\, 
         \$19741%now\, \$19218_v%next\, \$19218_v%now\, \$19713%next\, 
         \$19713%now\, \$19018_v%next\, \$19018_v%now\, \$19230_v%next\, 
         \$19230_v%now\, \$19350_v%next\, \$19350_v%now\, \$19659_hd%next\, 
         \$19659_hd%now\, \$19844%next\, \$19844%now\, \$v5487%next\, 
         \$v5487%now\, \$19169_v%next\, \$19169_v%now\, \$19643_w%next\, 
         \$19643_w%now\, \$18841%next\, \$18841%now\, \$v5872%next\, 
         \$v5872%now\, \$19824_hd%next\, \$19824_hd%now\, \$19220%next\, 
         \$19220%now\, \$18683_hd%next\, \$18683_hd%now\, \$19308_v%next\, 
         \$19308_v%now\, \$18843%next\, \$18843%now\, \$18824_v%next\, 
         \$18824_v%now\, \$19256_v%next\, \$19256_v%now\, \$18877_v%next\, 
         \$18877_v%now\, \$19119_v%next\, \$19119_v%now\, \$19227%next\, 
         \$19227%now\, \$18832_v%next\, \$18832_v%now\, \$19717%next\, 
         \$19717%now\, \$19288_v%next\, \$19288_v%now\, \$v5873%next\, 
         \$v5873%now\, \$18888_next_acc%next\, \$18888_next_acc%now\, 
         \$18893_v%next\, \$18893_v%now\, \$18848%next\, \$18848%now\, 
         \$19324_f0%next\, \$19324_f0%now\, \$18442_cy%next\, 
         \$18442_cy%now\, \$18599_hd%next\, \$18599_hd%now\, \$18884_v%next\, 
         \$18884_v%now\, \$19559_w%next\, \$19559_w%now\, \$19595%next\, 
         \$19595%now\, \$18873_v%next\, \$18873_v%now\, \$19354_v%next\, 
         \$19354_v%now\, \$19307_v%next\, \$19307_v%now\, \$19880_w%next\, 
         \$19880_w%now\, \$19910_hd%next\, \$19910_hd%now\, \$v5611%next\, 
         \$v5611%now\, \$19177_v%next\, \$19177_v%now\, \$18598_w%next\, 
         \$18598_w%now\, \$19423_v%next\, \$19423_v%now\, \$19075_v%next\, 
         \$19075_v%now\, \$18765%next\, \$18765%now\, \$19357_v%next\, 
         \$19357_v%now\, \$19909_w%next\, \$19909_w%now\, \$18830_v%next\, 
         \$18830_v%now\, \$18711_w%next\, \$18711_w%now\, \$18450%next\, 
         \$18450%now\, \$19761%next\, \$19761%now\, \$19450_v%next\, 
         \$19450_v%now\, \$19222%next\, \$19222%now\, \$19851_hd%next\, 
         \$19851_hd%now\, \$v5870%next\, \$v5870%now\, \$18980_v%next\, 
         \$18980_v%now\, \$19279_v%next\, \$19279_v%now\, \$18577%next\, 
         \$18577%now\, \$18822_v%next\, \$18822_v%now\, \$19312_v%next\, 
         \$19312_v%now\, \$18999_v%next\, \$18999_v%now\, \$18584_hd%next\, 
         \$18584_hd%now\, \$18834_v%next\, \$18834_v%now\, \$19817%next\, 
         \$19817%now\, \$v5557%next\, \$v5557%now\, \$19267_hd%next\, 
         \$19267_hd%now\, \$v5577%next\, \$v5577%now\, \$18828_v%next\, 
         \$18828_v%now\, \$19721_hd%next\, \$19721_hd%now\, \$18457%next\, 
         \$18457%now\, \$19296_v%next\, \$19296_v%now\, \$v5607%next\, 
         \$v5607%now\, \$19246_v%next\, \$19246_v%now\, \$18638_hd%next\, 
         \$18638_hd%now\, \$19720_w%next\, \$19720_w%now\, \$18852%next\, 
         \$18852%now\, \$18668_hd%next\, \$18668_hd%now\, \$19628_w%next\, 
         \$19628_w%now\, \$19902%next\, \$19902%now\, \$v5537%next\, 
         \$v5537%now\, \$18565%next\, \$18565%now\, \$18667_w%next\, 
         \$18667_w%now\, \$19209_v%next\, \$19209_v%now\, \$19309_v%next\, 
         \$19309_v%now\, \$19342%next\, \$19342%now\, \$v5869%next\, 
         \$v5869%now\, \$19478_v%next\, \$19478_v%now\, \$18745_hd%next\, 
         \$18745_hd%now\, \$19364_v%next\, \$19364_v%now\, \$19185_v%next\, 
         \$19185_v%now\, \$19930%next\, \$19930%now\, \$19704%next\, 
         \$19704%now\, \$19274_v%next\, \$19274_v%now\, \$19201_v%next\, 
         \$19201_v%now\, \$18961_v%next\, \$18961_v%now\, \$19850_w%next\, 
         \$19850_w%now\, \$18846%next\, \$18846%now\, \$19934_hd%next\, 
         \$19934_hd%now\, \$18859%next\, \$18859%now\, 
         \$18855_next_env%next\, \$18855_next_env%now\, \$19906%next\, 
         \$19906%now\, \$19235_v%next\, \$19235_v%now\, \$18881_hd%next\, 
         \$18881_hd%now\, \$v5824%next\, \$v5824%now\, \$19094_v%next\, 
         \$19094_v%now\, \$19448_v%next\, \$19448_v%now\, \$18821_v%next\, 
         \$18821_v%now\, \$18769_hd%next\, \$18769_hd%now\, \$19866_hd%next\, 
         \$19866_hd%now\, \$18619%next\, \$18619%now\, \$18875_v%next\, 
         \$18875_v%now\, \$v5619%next\, \$v5619%now\, \$18637_w%next\, 
         \$18637_w%now\, \$19553%next\, \$19553%now\, \$v5507%next\, 
         \$v5507%now\ : value(0 to 31) := (others => '0');
  signal \$19198_binop_compare6454381_arg%next\, 
         \$19198_binop_compare6454381_arg%now\, 
         \$19174_binop_compare6454378_arg%next\, 
         \$19174_binop_compare6454378_arg%now\, 
         \$18901_binop_int6434361_arg%next\, 
         \$18901_binop_int6434361_arg%now\, 
         \$19091_binop_int6434371_arg%next\, 
         \$19091_binop_int6434371_arg%now\, 
         \$19182_binop_compare6454379_arg%next\, 
         \$19182_binop_compare6454379_arg%now\, 
         \$19053_binop_int6434369_arg%next\, 
         \$19053_binop_int6434369_arg%now\, \$19311%next\, \$19311%now\, 
         \$18958_binop_int6434364_arg%next\, 
         \$18958_binop_int6434364_arg%now\, 
         \$18939_binop_int6434363_arg%next\, 
         \$18939_binop_int6434363_arg%now\, \$19281%next\, \$19281%now\, 
         \$19116_binop_int6434373_arg%next\, 
         \$19116_binop_int6434373_arg%now\, \$19300%next\, \$19300%now\, 
         \$18920_binop_int6434362_arg%next\, 
         \$18920_binop_int6434362_arg%now\, 
         \$19206_binop_compare6454382_arg%next\, 
         \$19206_binop_compare6454382_arg%now\, 
         \$18996_binop_int6434366_arg%next\, 
         \$18996_binop_int6434366_arg%now\, 
         \$18977_binop_int6434365_arg%next\, 
         \$18977_binop_int6434365_arg%now\, 
         \$19015_binop_int6434367_arg%next\, 
         \$19015_binop_int6434367_arg%now\, 
         \$19034_binop_int6434368_arg%next\, 
         \$19034_binop_int6434368_arg%now\, 
         \$19135_binop_int6434374_arg%next\, 
         \$19135_binop_int6434374_arg%now\, 
         \$19166_binop_compare6454377_arg%next\, 
         \$19166_binop_compare6454377_arg%now\, \$19273%next\, \$19273%now\, 
         \$19290%next\, \$19290%now\, \$19072_binop_int6434370_arg%next\, 
         \$19072_binop_int6434370_arg%now\, 
         \$19190_binop_compare6454380_arg%next\, 
         \$19190_binop_compare6454380_arg%now\ : value(0 to 153) := (others => '0');
  signal \$19116_binop_int6434373_result%next\, 
         \$19116_binop_int6434373_result%now\, 
         \$19166_binop_compare6454377_result%next\, 
         \$19166_binop_compare6454377_result%now\, 
         \$19387_compbranch6504394_result%next\, 
         \$19387_compbranch6504394_result%now\, 
         \$19034_binop_int6434368_result%next\, 
         \$19034_binop_int6434368_result%now\, 
         \$18796_make_block_n646_result%next\, 
         \$18796_make_block_n646_result%now\, 
         \$18920_binop_int6434362_result%next\, 
         \$18920_binop_int6434362_result%now\, 
         \$19091_binop_int6434371_result%next\, 
         \$19091_binop_int6434371_result%now\, 
         \$19380_compbranch6504393_result%next\, 
         \$19380_compbranch6504393_result%now\, 
         \$19394_compbranch6504395_result%next\, 
         \$19394_compbranch6504395_result%now\, 
         \$18794_apply638_result%next\, \$18794_apply638_result%now\, 
         \$18901_binop_int6434361_result%next\, 
         \$18901_binop_int6434361_result%now\, 
         \$19174_binop_compare6454378_result%next\, 
         \$19174_binop_compare6454378_result%now\, 
         \$18996_binop_int6434366_result%next\, 
         \$18996_binop_int6434366_result%now\, 
         \$19198_binop_compare6454381_result%next\, 
         \$19198_binop_compare6454381_result%now\, 
         \$19053_binop_int6434369_result%next\, 
         \$19053_binop_int6434369_result%now\, 
         \$19182_binop_compare6454379_result%next\, 
         \$19182_binop_compare6454379_result%now\, 
         \$19206_binop_compare6454382_result%next\, 
         \$19206_binop_compare6454382_result%now\, 
         \$19015_binop_int6434367_result%next\, 
         \$19015_binop_int6434367_result%now\, 
         \$18977_binop_int6434365_result%next\, 
         \$18977_binop_int6434365_result%now\, \result4928%next\, 
         \result4928%now\, \$19366_compbranch6504391_result%next\, 
         \$19366_compbranch6504391_result%now\, 
         \$19333_compbranch6504388_result%next\, 
         \$19333_compbranch6504388_result%now\, 
         \$19135_binop_int6434374_result%next\, 
         \$19135_binop_int6434374_result%now\, 
         \$19373_compbranch6504392_result%next\, 
         \$19373_compbranch6504392_result%now\, 
         \$18795_offsetclosure_n639_result%next\, 
         \$18795_offsetclosure_n639_result%now\, 
         \$19401_compbranch6504396_result%next\, 
         \$19401_compbranch6504396_result%now\, 
         \$19190_binop_compare6454380_result%next\, 
         \$19190_binop_compare6454380_result%now\, 
         \$19072_binop_int6434370_result%next\, 
         \$19072_binop_int6434370_result%now\, 
         \$18958_binop_int6434364_result%next\, 
         \$18958_binop_int6434364_result%now\, 
         \$18797_branch_if648_result%next\, \$18797_branch_if648_result%now\, 
         \$18939_binop_int6434363_result%next\, 
         \$18939_binop_int6434363_result%now\, 
         \$19326_compbranch6504387_result%next\, 
         \$19326_compbranch6504387_result%now\ : value(0 to 121) := (others => '0');
  
  begin
    process (clk)
            begin
            if rising_edge(clk) then
                 if \$ram_write_request\ = '1' then
                    ram(\$ram_ptr_write\) <= \$ram_write\;
                 end if;
                 \$ram_value\ <= ram(\$ram_ptr\);
            end if;
        end process;
    
    process (clk)
            begin
            if rising_edge(clk) then
                 if \$global_end_write_request\ = '1' then
                    global_end(\$global_end_ptr_write\) <= \$global_end_write\;
                 end if;
                 \$global_end_value\ <= global_end(\$global_end_ptr\);
            end if;
        end process;
    
    process (clk)
            begin
            if rising_edge(clk) then
                 if \$code_write_request\ = '1' then
                    code(\$code_ptr_write\) <= \$code_write\;
                 end if;
                 \$code_value\ <= code(\$code_ptr\);
            end if;
        end process;
    
    process (reset,clk)
      begin
      if reset = '1' then
        \$18606%now\ <= (others => '0');
        \$19190_binop_compare6454380_arg%now\ <= (others => '0');
        \$v4743%now\ <= (others => '0');
        \$19072_binop_int6434370_arg%now\ <= (others => '0');
        \$18910_modulo6684349_id%now\ <= (others => '0');
        \$19299%now\ <= (others => '0');
        \$19069_modulo6684349_id%now\ <= (others => '0');
        \$v5526%now\ <= (others => '0');
        \$v4663%now\ <= (others => '0');
        \$v5913%now\ <= (others => '0');
        \$18602%now\ <= (others => '0');
        \$v5541%now\ <= (others => '0');
        \$18809%now\ <= (others => '0');
        \$18751%now\ <= (others => '0');
        \$19272%now\ <= (others => '0');
        \$v5486%now\ <= (others => '0');
        \$v5513%now\ <= (others => '0');
        \$18729%now\ <= (others => '0');
        \$v5507%now\ <= (others => '0');
        \$18801%now\ <= (others => '0');
        \$19779_loop666_id%now\ <= (others => '0');
        \$18775%now\ <= (others => '0');
        \$19874%now\ <= (others => '0');
        \$v5715%now\ <= (others => '0');
        \$18974_modulo6684349_id%now\ <= (others => '0');
        \$19828%now\ <= (others => '0');
        \$v4961%now\ <= (others => '0');
        \$v4499%now\ <= (others => '0');
        \$19326_compbranch6504387_result%now\ <= (others => '0');
        \$v5326%now\ <= (others => '0');
        \$v5484%now\ <= (others => '0');
        \$18504%now\ <= (others => '0');
        \$v5643%now\ <= (others => '0');
        \$18945_modulo6684356_result%now\ <= (others => '0');
        \$18933_modulo6684357_id%now\ <= (others => '0');
        \$19250%now\ <= (others => '0');
        \$18624%now\ <= (others => '0');
        \$v4650%now\ <= (others => '0');
        \$19553%now\ <= (others => '0');
        \$18637_w%now\ <= (others => '0');
        \$19380_compbranch6504393_id%now\ <= (others => '0');
        \$v5619%now\ <= (others => '0');
        \$18835%now\ <= (others => '0');
        \$19579%now\ <= (others => '0');
        \$19758%now\ <= (others => '0');
        \$19085_modulo6684357_result%now\ <= (others => '0');
        \$18776%now\ <= (others => '0');
        \$18875_v%now\ <= (others => '0');
        \$19132_modulo6684349_id%now\ <= (others => '0');
        \$18619%now\ <= (others => '0');
        \$19163_forever6704376_arg%now\ <= (others => '0');
        \$v4604%now\ <= (others => '0');
        \$v5699%now\ <= (others => '0');
        \$19292%now\ <= (others => '0');
        \$v5634%now\ <= (others => '0');
        \$19416_w36574398_result%now\ <= (others => '0');
        \$18993_modulo6684349_result%now\ <= (others => '0');
        \$18581%now\ <= (others => '0');
        \$19866_hd%now\ <= (others => '0');
        \$v5287%now\ <= (others => '0');
        \$v4467%now\ <= (others => '0');
        \$18900%now\ <= (others => '0');
        \$v4470%now\ <= (others => '0');
        \$v4325%now\ <= (others => '0');
        \$18696%now\ <= (others => '0');
        \$19245%now\ <= (others => '0');
        \$19024_modulo6684349_result%now\ <= (others => '0');
        \$18945_modulo6684356_arg%now\ <= (others => '0');
        \$19689%now\ <= (others => '0');
        \$v4577%now\ <= (others => '0');
        \$19140_r%now\ <= (others => '0');
        \$18802%now\ <= (others => '0');
        \$v5076%now\ <= (others => '0');
        \$19001_r%now\ <= (others => '0');
        \$v5532%now\ <= (others => '0');
        \$19501%now\ <= (others => '0');
        \$18769_hd%now\ <= (others => '0');
        \$v5152%now\ <= (others => '0');
        \$v4703%now\ <= (others => '0');
        \$19122_modulo6684356_result%now\ <= (others => '0');
        \$19499_aux664_id%now\ <= (others => '0');
        \$18483%now\ <= (others => '0');
        \$19290%now\ <= (others => '0');
        \$19273%now\ <= (others => '0');
        \$19104_modulo6684357_id%now\ <= (others => '0');
        \$v4710%now\ <= (others => '0');
        \$v4814%now\ <= (others => '0');
        \$19170_res%now\ <= (others => '0');
        \$18924_res%now\ <= (others => '0');
        \$19863%now\ <= (others => '0');
        \$18821_v%now\ <= (others => '0');
        \$19827%now\ <= (others => '0');
        \$19432%now\ <= (others => '0');
        \$19448_v%now\ <= (others => '0');
        \$18630%now\ <= (others => '0');
        \$19094_v%now\ <= (others => '0');
        \$v4535%now\ <= (others => '0');
        \$v5551%now\ <= (others => '0');
        \$19028_modulo6684357_result%now\ <= (others => '0');
        \$18939_binop_int6434363_result%now\ <= (others => '0');
        \$v5824%now\ <= (others => '0');
        \$18788%now\ <= (others => '0');
        \$v5226%now\ <= (others => '0');
        \$18582%now\ <= (others => '0');
        \$19081_modulo6684349_arg%now\ <= (others => '0');
        \$v5013%now\ <= (others => '0');
        \$18881_hd%now\ <= (others => '0');
        \$19525%now\ <= (others => '0');
        \$18509%now\ <= (others => '0');
        \$18793_make_block579_result%now\ <= (others => '0');
        \$18974_modulo6684349_arg%now\ <= (others => '0');
        \$19235_v%now\ <= (others => '0');
        \$v4515%now\ <= (others => '0');
        \$v5323%now\ <= (others => '0');
        \$18655%now\ <= (others => '0');
        \$19906%now\ <= (others => '0');
        \$v5592%now\ <= (others => '0');
        \$19194_res%now\ <= (others => '0');
        \$18990_modulo6684357_result%now\ <= (others => '0');
        \$19947%now\ <= (others => '0');
        \$19672%now\ <= (others => '0');
        \$v5692%now\ <= (others => '0');
        \$18474%now\ <= (others => '0');
        \$19641%now\ <= (others => '0');
        \$18855_next_env%now\ <= (others => '0');
        \$v5158%now\ <= (others => '0');
        \$19040_modulo6684356_id%now\ <= (others => '0');
        \$v5369%now\ <= (others => '0');
        \$v5733%now\ <= (others => '0');
        \$19661%now\ <= (others => '0');
        \$v5414%now\ <= (others => '0');
        \$v4443%now\ <= (others => '0');
        \$18876%now\ <= (others => '0');
        \$19653%now\ <= (others => '0');
        \$19508%now\ <= (others => '0');
        \$19358%now\ <= (others => '0');
        \$v5151%now\ <= (others => '0');
        \$v5594%now\ <= (others => '0');
        \$19043_modulo6684349_result%now\ <= (others => '0');
        \$18859%now\ <= (others => '0');
        \$v4830%now\ <= (others => '0');
        \$v5117%now\ <= (others => '0');
        \$19445%now\ <= (others => '0');
        \$18867%now\ <= (others => '0');
        \$v5752%now\ <= (others => '0');
        \$18865%now\ <= (others => '0');
        \$19890%now\ <= (others => '0');
        \$v4511%now\ <= (others => '0');
        \$18455%now\ <= (others => '0');
        \$18512%now\ <= (others => '0');
        \$v4590%now\ <= (others => '0');
        \$19427%now\ <= (others => '0');
        \$19934_hd%now\ <= (others => '0');
        \$18846%now\ <= (others => '0');
        \$18524_loop666_result%now\ <= (others => '0');
        \$v4472%now\ <= (others => '0');
        \$19723%now\ <= (others => '0');
        \$18778%now\ <= (others => '0');
        \$18694%now\ <= (others => '0');
        \$v5759%now\ <= (others => '0');
        \$19066_modulo6684357_result%now\ <= (others => '0');
        \$19850_w%now\ <= (others => '0');
        \$19419%now\ <= (others => '0');
        \$18961_v%now\ <= (others => '0');
        \$19201_v%now\ <= (others => '0');
        \$v5703%now\ <= (others => '0');
        \$19274_v%now\ <= (others => '0');
        \$19394_compbranch6504395_arg%now\ <= (others => '0');
        \$v5320%now\ <= (others => '0');
        \$19166_binop_compare6454377_arg%now\ <= (others => '0');
        \$v5212%now\ <= (others => '0');
        \$19704%now\ <= (others => '0');
        \$19930%now\ <= (others => '0');
        \$v5721%now\ <= (others => '0');
        \$19458%now\ <= (others => '0');
        \$19185_v%now\ <= (others => '0');
        \$v5586%now\ <= (others => '0');
        \$18738_next%now\ <= (others => '0');
        \$19364_v%now\ <= (others => '0');
        \$v5234%now\ <= (others => '0');
        \$v5760%now\ <= (others => '0');
        \$18974_modulo6684349_result%now\ <= (others => '0');
        \$19797_next%now\ <= (others => '0');
        \$18745_hd%now\ <= (others => '0');
        \$18797_branch_if648_result%now\ <= (others => '0');
        \$19589_copy_root_in_ram6634353_id%now\ <= (others => '0');
        \$v5766%now\ <= (others => '0');
        \$19478_v%now\ <= (others => '0');
        \$19752%now\ <= (others => '0');
        \$v4616%now\ <= (others => '0');
        \$19894%now\ <= (others => '0');
        \$19819%now\ <= (others => '0');
        \$19489%now\ <= (others => '0');
        \$v5776%now\ <= (others => '0');
        \$v5019%now\ <= (others => '0');
        \$18807%now\ <= (others => '0');
        \$19504%now\ <= (others => '0');
        \$18650%now\ <= (others => '0');
        \$18837%now\ <= (others => '0');
        \$18569%now\ <= (others => '0');
        \$19129_modulo6684357_id%now\ <= (others => '0');
        \$18805%now\ <= (others => '0');
        \$v5869%now\ <= (others => '0');
        \$19112%now\ <= (others => '0');
        \$19135_binop_int6434374_arg%now\ <= (others => '0');
        \$19002_modulo6684356_arg%now\ <= (others => '0');
        \$v5515%now\ <= (others => '0');
        \$19319%now\ <= (others => '0');
        \$v5646%now\ <= (others => '0');
        \$v4952%now\ <= (others => '0');
        \$v5610%now\ <= (others => '0');
        \$v5683%now\ <= (others => '0');
        \$18958_binop_int6434364_result%now\ <= (others => '0');
        \$19342%now\ <= (others => '0');
        \$19657%now\ <= (others => '0');
        \$19777%now\ <= (others => '0');
        \$19620%now\ <= (others => '0');
        \$18793_make_block579_id%now\ <= (others => '0');
        \$18521_loop666_arg%now\ <= (others => '0');
        \$19803%now\ <= (others => '0');
        \$19217%now\ <= (others => '0');
        \$v4949%now\ <= (others => '0');
        \$19486%now\ <= (others => '0');
        \$v5857%now\ <= (others => '0');
        \$18482%now\ <= (others => '0');
        \$v4692%now\ <= (others => '0');
        \$19309_v%now\ <= (others => '0');
        \$18529%now\ <= (others => '0');
        \$19916%now\ <= (others => '0');
        \$v5686%now\ <= (others => '0');
        \$v4854%now\ <= (others => '0');
        \$v4628%now\ <= (others => '0');
        \$18703%now\ <= (others => '0');
        \$v5506%now\ <= (others => '0');
        \$v4926%now\ <= (others => '0');
        \$19829%now\ <= (others => '0');
        \$v4523%now\ <= (others => '0');
        \$v4569%now\ <= (others => '0');
        \$v5749%now\ <= (others => '0');
        \$19209_v%now\ <= (others => '0');
        \$19482%now\ <= (others => '0');
        \$19611%now\ <= (others => '0');
        \$19811_copy_root_in_ram6634341_id%now\ <= (others => '0');
        \$19784%now\ <= (others => '0');
        \$18502%now\ <= (others => '0');
        \$v4770%now\ <= (others => '0');
        \$18667_w%now\ <= (others => '0');
        \$19434%now\ <= (others => '0');
        \$19333_compbranch6504388_arg%now\ <= (others => '0');
        \$19732%now\ <= (others => '0');
        \$19609%now\ <= (others => '0');
        \$19714_next%now\ <= (others => '0');
        \$18815%now\ <= (others => '0');
        \$v5210%now\ <= (others => '0');
        \$18565%now\ <= (others => '0');
        \$v4491%now\ <= (others => '0');
        \$19076_res%now\ <= (others => '0');
        \$v4727%now\ <= (others => '0');
        \$19015_binop_int6434367_id%now\ <= (others => '0');
        \$18986_modulo6684349_arg%now\ <= (others => '0');
        \$v4734%now\ <= (others => '0');
        \$19656%now\ <= (others => '0');
        \$19496_aux664_arg%now\ <= (others => '0');
        \$18480%now\ <= (others => '0');
        \$v5537%now\ <= (others => '0');
        \$18458%now\ <= (others => '0');
        \$18993_modulo6684349_arg%now\ <= (others => '0');
        \$v5655%now\ <= (others => '0');
        \$19294%now\ <= (others => '0');
        \$v5828%now\ <= (others => '0');
        \$19583%now\ <= (others => '0');
        \$v5838%now\ <= (others => '0');
        \$19163_forever6704376_id%now\ <= (others => '0');
        \$18723%now\ <= (others => '0');
        \$v4481%now\ <= (others => '0');
        \$v5640%now\ <= (others => '0');
        \$19314%now\ <= (others => '0');
        \$18762%now\ <= (others => '0');
        \$19034_binop_int6434368_arg%now\ <= (others => '0');
        \$v4728%now\ <= (others => '0');
        \$v4596%now\ <= (others => '0');
        \$19062_modulo6684349_result%now\ <= (others => '0');
        \$18914_modulo6684357_arg%now\ <= (others => '0');
        \$18590%now\ <= (others => '0');
        \$19902%now\ <= (others => '0');
        \$18670%now\ <= (others => '0');
        \$v5604%now\ <= (others => '0');
        \$19248%now\ <= (others => '0');
        \$19088_modulo6684349_result%now\ <= (others => '0');
        \$19464%now\ <= (others => '0');
        \$19072_binop_int6434370_result%now\ <= (others => '0');
        \$v4761%now\ <= (others => '0');
        \$19816%now\ <= (others => '0');
        \$19081_modulo6684349_result%now\ <= (others => '0');
        \$v4845%now\ <= (others => '0');
        \$v4631%now\ <= (others => '0');
        \$19326_compbranch6504387_arg%now\ <= (others => '0');
        \$v5035%now\ <= (others => '0');
        \$18685%now\ <= (others => '0');
        \$v5603%now\ <= (others => '0');
        \$19628_w%now\ <= (others => '0');
        \$v5582%now\ <= (others => '0');
        \$18948_modulo6684349_arg%now\ <= (others => '0');
        \$v5060%now\ <= (others => '0');
        \$18668_hd%now\ <= (others => '0');
        \$v4552%now\ <= (others => '0');
        \$19187_compare6444358_result%now\ <= (others => '0');
        \$v5378%now\ <= (others => '0');
        \$19623%now\ <= (others => '0');
        \$v5052%now\ <= (others => '0');
        \$v4946%now\ <= (others => '0');
        \$18664%now\ <= (others => '0');
        \$18646%now\ <= (others => '0');
        \$18852%now\ <= (others => '0');
        \$18485%now\ <= (others => '0');
        \$19190_binop_compare6454380_result%now\ <= (others => '0');
        \$19043_modulo6684349_arg%now\ <= (others => '0');
        \$v4936%now\ <= (others => '0');
        \$v4417%now\ <= (others => '0');
        \$18447%now\ <= (others => '0');
        \$v4992%now\ <= (others => '0');
        \$v5702%now\ <= (others => '0');
        \$18967_modulo6684349_arg%now\ <= (others => '0');
        \$v5481%now\ <= (others => '0');
        \$18952_modulo6684357_result%now\ <= (others => '0');
        \$18662%now\ <= (others => '0');
        \$18600%now\ <= (others => '0');
        \$v5244%now\ <= (others => '0');
        \$19600%now\ <= (others => '0');
        \$19838_copy_root_in_ram6634340_result%now\ <= (others => '0');
        \$19885%now\ <= (others => '0');
        \$19685%now\ <= (others => '0');
        \$19187_compare6444358_id%now\ <= (others => '0');
        \$18926_modulo6684356_id%now\ <= (others => '0');
        \$19720_w%now\ <= (others => '0');
        \$v5530%now\ <= (others => '0');
        \$18644%now\ <= (others => '0');
        \$18466_loop666_id%now\ <= (others => '0');
        \$18638_hd%now\ <= (others => '0');
        \$v4674%now\ <= (others => '0');
        \$v5250%now\ <= (others => '0');
        \$18563%now\ <= (others => '0');
        \$19062_modulo6684349_id%now\ <= (others => '0');
        \$18645%now\ <= (others => '0');
        \$19897%now\ <= (others => '0');
        \$19139_res%now\ <= (others => '0');
        \$19347_fill6534389_arg%now\ <= (others => '0');
        \$19495_loop665_arg%now\ <= (others => '0');
        \$v4695%now\ <= (others => '0');
        \$18576%now\ <= (others => '0');
        \$18578%now\ <= (others => '0');
        \$18440_make_block579_arg%now\ <= (others => '0');
        \$19157_forever6704375_id%now\ <= (others => '0');
        \$19246_v%now\ <= (others => '0');
        \$19495_loop665_id%now\ <= (others => '0');
        \$19515_next%now\ <= (others => '0');
        \$v4563%now\ <= (others => '0');
        \$v4908%now\ <= (others => '0');
        \$18635%now\ <= (others => '0');
        \$19251%now\ <= (others => '0');
        \$19648%now\ <= (others => '0');
        \$18613_copy_root_in_ram6634346_id%now\ <= (others => '0');
        \$19780_loop665_arg%now\ <= (others => '0');
        \$18571_copy_root_in_ram6634345_arg%now\ <= (others => '0');
        \$v5120%now\ <= (others => '0');
        \$19854%now\ <= (others => '0');
        \$v4988%now\ <= (others => '0');
        \$v5607%now\ <= (others => '0');
        \$19848%now\ <= (others => '0');
        \$19232%now\ <= (others => '0');
        \$19814%now\ <= (others => '0');
        \$v4680%now\ <= (others => '0');
        \$18906_r%now\ <= (others => '0');
        \$v5127%now\ <= (others => '0');
        \$18620%now\ <= (others => '0');
        \$19887%now\ <= (others => '0');
        \$19296_v%now\ <= (others => '0');
        \$18709%now\ <= (others => '0');
        \$v4805%now\ <= (others => '0');
        \$v5514%now\ <= (others => '0');
        \$18913_r%now\ <= (others => '0');
        \$18457%now\ <= (others => '0');
        \$19269%now\ <= (others => '0');
        \$19569%now\ <= (others => '0');
        \$v5823%now\ <= (others => '0');
        \$v5164%now\ <= (others => '0');
        \$19721_hd%now\ <= (others => '0');
        \$v5831%now\ <= (others => '0');
        \$v4740%now\ <= (others => '0');
        \$v5308%now\ <= (others => '0');
        \$v4995%now\ <= (others => '0');
        \$v4601%now\ <= (others => '0');
        \$18484%now\ <= (others => '0');
        \$18733%now\ <= (others => '0');
        \$v4660%now\ <= (others => '0');
        \$19408_argument3%now\ <= (others => '0');
        \$18828_v%now\ <= (others => '0');
        \$19390_b%now\ <= (others => '0');
        \$19727%now\ <= (others => '0');
        \$18510%now\ <= (others => '0');
        \$19662%now\ <= (others => '0');
        \$v5577%now\ <= (others => '0');
        \$19015_binop_int6434367_arg%now\ <= (others => '0');
        \$19413%now\ <= (others => '0');
        \$v4584%now\ <= (others => '0');
        \$19845%now\ <= (others => '0');
        \$19337_compare6444359_id%now\ <= (others => '0');
        \$19698%now\ <= (others => '0');
        \$18566%now\ <= (others => '0');
        \$18767%now\ <= (others => '0');
        \$19359%now\ <= (others => '0');
        \$18977_binop_int6434365_arg%now\ <= (others => '0');
        \$v4878%now\ <= (others => '0');
        \$19267_hd%now\ <= (others => '0');
        \$19679%now\ <= (others => '0');
        \$v5195%now\ <= (others => '0');
        \$v4433%now\ <= (others => '0');
        \$18864%now\ <= (others => '0');
        \$18996_binop_int6434366_arg%now\ <= (others => '0');
        \$19599%now\ <= (others => '0');
        \$19526_forever6704355_arg%now\ <= (others => '0');
        \$19578%now\ <= (others => '0');
        \$18605%now\ <= (others => '0');
        \$19558%now\ <= (others => '0');
        \$19280%now\ <= (others => '0');
        \$v5278%now\ <= (others => '0');
        \$v5557%now\ <= (others => '0');
        \$19817%now\ <= (others => '0');
        \$19238_w6514383_arg%now\ <= (others => '0');
        \$v5284%now\ <= (others => '0');
        \$v5905%now\ <= (others => '0');
        \$19488%now\ <= (others => '0');
        \$19474%now\ <= (others => '0');
        \$v5564%now\ <= (others => '0');
        \$18591%now\ <= (others => '0');
        \$v4568%now\ <= (others => '0');
        \$v5883%now\ <= (others => '0');
        \$v5555%now\ <= (others => '0');
        \$19726%now\ <= (others => '0');
        \$v4842%now\ <= (others => '0');
        \$18834_v%now\ <= (others => '0');
        \$19401_compbranch6504396_result%now\ <= (others => '0');
        \$18699%now\ <= (others => '0');
        \$18680%now\ <= (others => '0');
        \$19751%now\ <= (others => '0');
        \$19157_forever6704375_arg%now\ <= (others => '0');
        \$18584_hd%now\ <= (others => '0');
        \$19867%now\ <= (others => '0');
        \$v5465%now\ <= (others => '0');
        \$18999_v%now\ <= (others => '0');
        \$18623%now\ <= (others => '0');
        \$19754%now\ <= (others => '0');
        \$19825%now\ <= (others => '0');
        \$19312_v%now\ <= (others => '0');
        \$18936_modulo6684349_arg%now\ <= (others => '0');
        \$18460%now\ <= (others => '0');
        \$19596%now\ <= (others => '0');
        \$18795_offsetclosure_n639_result%now\ <= (others => '0');
        \$19918%now\ <= (others => '0');
        \$v4328%now\ <= (others => '0');
        \$19373_compbranch6504392_result%now\ <= (others => '0');
        \$v5247%now\ <= (others => '0');
        \$v4543%now\ <= (others => '0');
        \$v5420%now\ <= (others => '0');
        \$19505%now\ <= (others => '0');
        \$18570%now\ <= (others => '0');
        \$v5263%now\ <= (others => '0');
        \$19391_compare6444359_id%now\ <= (others => '0');
        \$v5835%now\ <= (others => '0');
        \$18962_res%now\ <= (others => '0');
        \$18822_v%now\ <= (others => '0');
        \$v5614%now\ <= (others => '0');
        \$v5027%now\ <= (others => '0');
        \$18610%now\ <= (others => '0');
        \$v5069%now\ <= (others => '0');
        \$18684%now\ <= (others => '0');
        \$19535_copy_root_in_ram6634354_id%now\ <= (others => '0');
        \$v5860%now\ <= (others => '0');
        \$v4414%now\ <= (others => '0');
        \$v5237%now\ <= (others => '0');
        \$19066_modulo6684357_arg%now\ <= (others => '0');
        \$19852%now\ <= (others => '0');
        \$18577%now\ <= (others => '0');
        \$v5533%now\ <= (others => '0');
        \$18553_forever6704348_arg%now\ <= (others => '0');
        \$19387_compbranch6504394_id%now\ <= (others => '0');
        \$18643%now\ <= (others => '0');
        \$18754%now\ <= (others => '0');
        \$18933_modulo6684357_arg%now\ <= (others => '0');
        \$19397_b%now\ <= (others => '0');
        \$19279_v%now\ <= (others => '0');
        \$18933_modulo6684357_result%now\ <= (others => '0');
        \$v5485%now\ <= (others => '0');
        \$19550%now\ <= (others => '0');
        \$18816%now\ <= (others => '0');
        \$19495_loop665_result%now\ <= (others => '0');
        \$v5516%now\ <= (others => '0');
        \$v5180%now\ <= (others => '0');
        \$18952_modulo6684357_arg%now\ <= (others => '0');
        \$19855%now\ <= (others => '0');
        \$v5426%now\ <= (others => '0');
        \$19313%now\ <= (others => '0');
        \$v5542%now\ <= (others => '0');
        \$19565%now\ <= (others => '0');
        \$v4863%now\ <= (others => '0');
        \$18980_v%now\ <= (others => '0');
        \$18521_loop666_id%now\ <= (others => '0');
        \$v5870%now\ <= (others => '0');
        \$19800_next%now\ <= (others => '0');
        \$19746%now\ <= (others => '0');
        \$19851_hd%now\ <= (others => '0');
        \$18488%now\ <= (others => '0');
        \$18746%now\ <= (others => '0');
        \$v5203%now\ <= (others => '0');
        \$19222%now\ <= (others => '0');
        \$v5290%now\ <= (others => '0');
        \$18796_make_block_n646_id%now\ <= (others => '0');
        \$19096_r%now\ <= (others => '0');
        \$19450_v%now\ <= (others => '0');
        \$19651%now\ <= (others => '0');
        \$v5130%now\ <= (others => '0');
        \$v5595%now\ <= (others => '0');
        \$v4699%now\ <= (others => '0');
        \$18559_copy_root_in_ram6634347_result%now\ <= (others => '0');
        \$18831%now\ <= (others => '0');
        \$v5123%now\ <= (others => '0');
        \$18829%now\ <= (others => '0');
        \$19761%now\ <= (others => '0');
        \$19547_copy_root_in_ram6634352_result%now\ <= (others => '0');
        \$v5737%now\ <= (others => '0');
        \$19676%now\ <= (others => '0');
        \$18450%now\ <= (others => '0');
        \$18982_r%now\ <= (others => '0');
        \$19179_compare6444358_arg%now\ <= (others => '0');
        \$v4462%now\ <= (others => '0');
        \$18717%now\ <= (others => '0');
        \$v5148%now\ <= (others => '0');
        \$18571_copy_root_in_ram6634345_id%now\ <= (others => '0');
        \$v5170%now\ <= (others => '0');
        \$19438%now\ <= (others => '0');
        \$19647%now\ <= (others => '0');
        \$19483%now\ <= (others => '0');
        \$19361_fill6544390_arg%now\ <= (others => '0');
        \$19861%now\ <= (others => '0');
        \$19211_compare6444358_id%now\ <= (others => '0');
        \$19786%now\ <= (others => '0');
        \$18725%now\ <= (others => '0');
        \$18459%now\ <= (others => '0');
        \$19135_binop_int6434374_result%now\ <= (others => '0');
        \$v5546%now\ <= (others => '0');
        \$19724%now\ <= (others => '0');
        \$18711_w%now\ <= (others => '0');
        \$18948_modulo6684349_result%now\ <= (others => '0');
        \$v5144%now\ <= (others => '0');
        \$19908%now\ <= (others => '0');
        \$19858%now\ <= (others => '0');
        \$18779%now\ <= (others => '0');
        \$v5272%now\ <= (others => '0');
        \$18612%now\ <= (others => '0');
        \$19303%now\ <= (others => '0');
        \$19551%now\ <= (others => '0');
        \$v5269%now\ <= (others => '0');
        \$19186_res%now\ <= (others => '0');
        \$18689%now\ <= (others => '0');
        \$19631%now\ <= (others => '0');
        \$18791_loop665_arg%now\ <= (others => '0');
        \$18905_res%now\ <= (others => '0');
        \$19694%now\ <= (others => '0');
        \$18755%now\ <= (others => '0');
        \$v5795%now\ <= (others => '0');
        \$v5202%now\ <= (others => '0');
        \$v5565%now\ <= (others => '0');
        \$v4923%now\ <= (others => '0');
        \$19835%now\ <= (others => '0');
        \$19588%now\ <= (others => '0');
        \$v4943%now\ <= (others => '0');
        \$19078_modulo6684356_id%now\ <= (others => '0');
        \$v5317%now\ <= (others => '0');
        \result4434%now\ <= (others => '0');
        \$v5512%now\ <= (others => '0');
        \$18465%now\ <= (others => '0');
        \$v4484%now\ <= (others => '0');
        \$18830_v%now\ <= (others => '0');
        \$19779_loop666_arg%now\ <= (others => '0');
        \$19616%now\ <= (others => '0');
        \$v4792%now\ <= (others => '0');
        \$19088_modulo6684349_arg%now\ <= (others => '0');
        \$19666%now\ <= (others => '0');
        \$19179_compare6444358_id%now\ <= (others => '0');
        \$19681_next%now\ <= (others => '0');
        \$18742%now\ <= (others => '0');
        \$18795_offsetclosure_n639_arg%now\ <= (others => '0');
        \$19384_compare6444359_id%now\ <= (others => '0');
        \$18993_modulo6684349_id%now\ <= (others => '0');
        \$19610%now\ <= (others => '0');
        \$18856_loop_push6494360_arg%now\ <= (others => '0');
        \$19909_w%now\ <= (others => '0');
        \$19686%now\ <= (others => '0');
        \$v4975%now\ <= (others => '0');
        \$19019_res%now\ <= (others => '0');
        \$v5534%now\ <= (others => '0');
        \$18479%now\ <= (others => '0');
        \$18525_loop665_result%now\ <= (others => '0');
        \$v5893%now\ <= (others => '0');
        \$19671%now\ <= (others => '0');
        \$v4475%now\ <= (others => '0');
        \$18734%now\ <= (others => '0');
        \$19128_r%now\ <= (others => '0');
        \$19750%now\ <= (others => '0');
        \$19499_aux664_arg%now\ <= (others => '0');
        \$19826%now\ <= (others => '0');
        \$18799_w1656_result%now\ <= (others => '0');
        \$18798_w652_result%now\ <= (others => '0');
        \$18467_loop665_arg%now\ <= (others => '0');
        \$19021_modulo6684356_id%now\ <= (others => '0');
        \$19088_modulo6684349_id%now\ <= (others => '0');
        \$19162%now\ <= (others => '0');
        \$v4851%now\ <= (others => '0');
        \$19357_v%now\ <= (others => '0');
        \$19097_modulo6684356_result%now\ <= (others => '0');
        \$v5580%now\ <= (others => '0');
        \$19012_modulo6684349_id%now\ <= (others => '0');
        \$18765%now\ <= (others => '0');
        \$v4893%now\ <= (others => '0');
        \$v5329%now\ <= (others => '0');
        \$19936%now\ <= (others => '0');
        \$19020_r%now\ <= (others => '0');
        \$19238_w6514383_result%now\ <= (others => '0');
        \$v5601%now\ <= (others => '0');
        \$18996_binop_int6434366_id%now\ <= (others => '0');
        \$v5511%now\ <= (others => '0');
        \$v4570%now\ <= (others => '0');
        \$19675%now\ <= (others => '0');
        \$18601%now\ <= (others => '0');
        \$v4565%now\ <= (others => '0');
        \$18552%now\ <= (others => '0');
        \$19077_r%now\ <= (others => '0');
        \$v5545%now\ <= (others => '0');
        \$v5031%now\ <= (others => '0');
        \$v5456%now\ <= (others => '0');
        \$v5161%now\ <= (others => '0');
        \$19075_v%now\ <= (others => '0');
        \$18791_loop665_result%now\ <= (others => '0');
        \$18750%now\ <= (others => '0');
        \$18718%now\ <= (others => '0');
        \$19849%now\ <= (others => '0');
        \$19059_modulo6684356_arg%now\ <= (others => '0');
        \$v4724%now\ <= (others => '0');
        \$19423_v%now\ <= (others => '0');
        \$19352%now\ <= (others => '0');
        \$19601_copy_root_in_ram6634352_result%now\ <= (others => '0');
        \$18789%now\ <= (others => '0');
        \$18977_binop_int6434365_id%now\ <= (others => '0');
        \$v5789%now\ <= (others => '0');
        \$v5450%now\ <= (others => '0');
        \$18681%now\ <= (others => '0');
        \$19206_binop_compare6454382_arg%now\ <= (others => '0');
        \$v5010%now\ <= (others => '0');
        \$19523%now\ <= (others => '0');
        \$18964_modulo6684356_id%now\ <= (others => '0');
        \$19923%now\ <= (others => '0');
        \$19361_fill6544390_result%now\ <= (others => '0');
        \$19535_copy_root_in_ram6634354_arg%now\ <= (others => '0');
        \$19564%now\ <= (others => '0');
        \$18770%now\ <= (others => '0');
        \$19790%now\ <= (others => '0');
        \$19509%now\ <= (others => '0');
        \$18598_w%now\ <= (others => '0');
        \$18462%now\ <= (others => '0');
        \$19873%now\ <= (others => '0');
        \$v5496%now\ <= (others => '0');
        \$v5573%now\ <= (others => '0');
        \$19177_v%now\ <= (others => '0');
        \$19320_forever6704386_arg%now\ <= (others => '0');
        \$19069_modulo6684349_arg%now\ <= (others => '0');
        \$v5225%now\ <= (others => '0');
        \$v5611%now\ <= (others => '0');
        \$v5063%now\ <= (others => '0');
        \$v5393%now\ <= (others => '0');
        \$19778%now\ <= (others => '0');
        \$19821%now\ <= (others => '0');
        \$v5174%now\ <= (others => '0');
        \$18494%now\ <= (others => '0');
        \$19333_compbranch6504388_result%now\ <= (others => '0');
        \$19441_arg%now\ <= (others => '0');
        \$18920_binop_int6434362_arg%now\ <= (others => '0');
        \$v5080%now\ <= (others => '0');
        \$18790_loop666_id%now\ <= (others => '0');
        \$v5763%now\ <= (others => '0');
        \$v5618%now\ <= (others => '0');
        \$18613_copy_root_in_ram6634346_result%now\ <= (others => '0');
        \$19498_loop665_arg%now\ <= (others => '0');
        \$19467_sp%now\ <= (others => '0');
        \$v4799%now\ <= (others => '0');
        \$19187_compare6444358_arg%now\ <= (others => '0');
        \$v4860%now\ <= (others => '0');
        \$18849%now\ <= (others => '0');
        \$18749%now\ <= (others => '0');
        \$18907_modulo6684356_id%now\ <= (others => '0');
        \$19794%now\ <= (others => '0');
        \$18863%now\ <= (others => '0');
        \$19910_hd%now\ <= (others => '0');
        \$18958_binop_int6434364_id%now\ <= (others => '0');
        \$v5135%now\ <= (others => '0');
        \$v4495%now\ <= (others => '0');
        \$19320_forever6704386_id%now\ <= (others => '0');
        \$19300%now\ <= (others => '0');
        \$19116_binop_int6434373_arg%now\ <= (others => '0');
        \$v5147%now\ <= (others => '0');
        \$v4899%now\ <= (others => '0');
        \$19333_compbranch6504388_id%now\ <= (others => '0');
        \$19880_w%now\ <= (others => '0');
        \$v5730%now\ <= (others => '0');
        \$19366_compbranch6504391_arg%now\ <= (others => '0');
        \$v5007%now\ <= (others => '0');
        \$19377_compare6444359_result%now\ <= (others => '0');
        \$19203_compare6444358_result%now\ <= (others => '0');
        \$v5570%now\ <= (others => '0');
        \$19664%now\ <= (others => '0');
        \$19637%now\ <= (others => '0');
        \$18926_modulo6684356_result%now\ <= (others => '0');
        \$v4431%now\ <= (others => '0');
        \$18854_sp%now\ <= (others => '0');
        \$19710%now\ <= (others => '0');
        \$19771%now\ <= (others => '0');
        \$19057_res%now\ <= (others => '0');
        \$18907_modulo6684356_arg%now\ <= (others => '0');
        \$18537%now\ <= (others => '0');
        \$19785%now\ <= (others => '0');
        \$18792_wait662_result%now\ <= (others => '0');
        \$18826%now\ <= (others => '0');
        \$19307_v%now\ <= (others => '0');
        \$19354_v%now\ <= (others => '0');
        \$19463%now\ <= (others => '0');
        \$19734%now\ <= (others => '0');
        \rdy4929%now\ <= (others => '0');
        \$18799_w1656_id%now\ <= (others => '0');
        \$19589_copy_root_in_ram6634353_result%now\ <= (others => '0');
        \$18472%now\ <= (others => '0');
        \$v4666%now\ <= (others => '0');
        \$19129_modulo6684357_arg%now\ <= (others => '0');
        \$v4458%now\ <= (others => '0');
        \$18873_v%now\ <= (others => '0');
        \$19038_res%now\ <= (others => '0');
        \$19595%now\ <= (others => '0');
        \$19883%now\ <= (others => '0');
        \$18677%now\ <= (others => '0');
        \$19249%now\ <= (others => '0');
        \$v5266%now\ <= (others => '0');
        \$19546%now\ <= (others => '0');
        \$v4767%now\ <= (others => '0');
        \$v5189%now\ <= (others => '0');
        \$v4442%now\ <= (others => '0');
        \$19891%now\ <= (others => '0');
        \$v5649%now\ <= (others => '0');
        \$v5199%now\ <= (others => '0');
        \$19559_w%now\ <= (others => '0');
        \$19920%now\ <= (others => '0');
        \$v4549%now\ <= (others => '0');
        \$18990_modulo6684357_id%now\ <= (others => '0');
        \$19107_modulo6684349_arg%now\ <= (others => '0');
        \$18520%now\ <= (others => '0');
        \$19420_w06554397_result%now\ <= (others => '0');
        \$18884_v%now\ <= (others => '0');
        \$18925_r%now\ <= (others => '0');
        \$19179_compare6444358_result%now\ <= (others => '0');
        \$19078_modulo6684356_arg%now\ <= (others => '0');
        \$v5103%now\ <= (others => '0');
        \$19522%now\ <= (others => '0');
        \$19544%now\ <= (others => '0');
        \$19243%now\ <= (others => '0');
        \$19718%now\ <= (others => '0');
        \$19148_modulo6684357_arg%now\ <= (others => '0');
        \$19538%now\ <= (others => '0');
        \$19255%now\ <= (others => '0');
        \$v4571%now\ <= (others => '0');
        \$19275%now\ <= (others => '0');
        \$19281%now\ <= (others => '0');
        \$18599_hd%now\ <= (others => '0');
        \$19836%now\ <= (others => '0');
        \$v4872%now\ <= (others => '0');
        \$19043_modulo6684349_id%now\ <= (others => '0');
        \$19884%now\ <= (others => '0');
        \$19871%now\ <= (others => '0');
        \$18851%now\ <= (others => '0');
        \$19557%now\ <= (others => '0');
        \$19517%now\ <= (others => '0');
        \$19532_forever6704350_id%now\ <= (others => '0');
        \$18782%now\ <= (others => '0');
        \$18526_aux664_id%now\ <= (others => '0');
        \$v4696%now\ <= (others => '0');
        \$19238_w6514383_id%now\ <= (others => '0');
        \$19582%now\ <= (others => '0');
        \$v5344%now\ <= (others => '0');
        \$19570%now\ <= (others => '0');
        \$v4619%now\ <= (others => '0');
        \$19888%now\ <= (others => '0');
        \$18794_apply638_id%now\ <= (others => '0');
        \$19497_loop666_id%now\ <= (others => '0');
        \$v4651%now\ <= (others => '0');
        \$18521_loop666_result%now\ <= (others => '0');
        \$19901%now\ <= (others => '0');
        \$18442_cy%now\ <= (others => '0');
        \$19444%now\ <= (others => '0');
        \$18549%now\ <= (others => '0');
        \$v5468%now\ <= (others => '0');
        \$18604%now\ <= (others => '0');
        \$18540%now\ <= (others => '0');
        \$18575%now\ <= (others => '0');
        \$19330_compare6444359_id%now\ <= (others => '0');
        \$19085_modulo6684357_arg%now\ <= (others => '0');
        \$19040_modulo6684356_result%now\ <= (others => '0');
        \$19324_f0%now\ <= (others => '0');
        \$v5083%now\ <= (others => '0');
        \$19540%now\ <= (others => '0');
        \$v5817%now\ <= (others => '0');
        \$19554%now\ <= (others => '0');
        \$19295%now\ <= (others => '0');
        \$19120_res%now\ <= (others => '0');
        \$18475%now\ <= (others => '0');
        \$18580%now\ <= (others => '0');
        \$v4612%now\ <= (others => '0');
        \$19005_modulo6684349_arg%now\ <= (others => '0');
        \$v4518%now\ <= (others => '0');
        \$v5637%now\ <= (others => '0');
        \$18848%now\ <= (others => '0');
        \$19801%now\ <= (others => '0');
        \$18893_v%now\ <= (others => '0');
        \$19913%now\ <= (others => '0');
        \$19262_forever6704385_id%now\ <= (others => '0');
        \$19210_res%now\ <= (others => '0');
        \$v5169%now\ <= (others => '0');
        \$18514%now\ <= (others => '0');
        \$18747%now\ <= (others => '0');
        \$v5402%now\ <= (others => '0');
        \$v5090%now\ <= (others => '0');
        \$v4408%now\ <= (others => '0');
        \$19304%now\ <= (others => '0');
        \$v5523%now\ <= (others => '0');
        \$18505%now\ <= (others => '0');
        \$18888_next_acc%now\ <= (others => '0');
        \$19376_b%now\ <= (others => '0');
        \$18688%now\ <= (others => '0');
        \$19100_modulo6684349_arg%now\ <= (others => '0');
        \$19412_sp%now\ <= (others => '0');
        \$v4407%now\ <= (others => '0');
        \$v5447%now\ <= (others => '0');
        \$19798%now\ <= (others => '0');
        \$v5003%now\ <= (others => '0');
        \$v5873%now\ <= (others => '0');
        \$19097_modulo6684356_arg%now\ <= (others => '0');
        \$v5550%now\ <= (others => '0');
        \$19626%now\ <= (others => '0');
        \$19471%now\ <= (others => '0');
        \$18721%now\ <= (others => '0');
        \$18971_modulo6684357_id%now\ <= (others => '0');
        \$18797_branch_if648_id%now\ <= (others => '0');
        \$v4704%now\ <= (others => '0');
        \$19288_v%now\ <= (others => '0');
        \$v5390%now\ <= (others => '0');
        \$19366_compbranch6504391_result%now\ <= (others => '0');
        \$v5462%now\ <= (others => '0');
        \$19914%now\ <= (others => '0');
        \$v5311%now\ <= (others => '0');
        \$18608%now\ <= (others => '0');
        \$19317%now\ <= (others => '0');
        \$19141_modulo6684356_result%now\ <= (others => '0');
        \$18511%now\ <= (others => '0');
        \$v4671%now\ <= (others => '0');
        \$19487%now\ <= (others => '0');
        \$18522_loop665_arg%now\ <= (others => '0');
        \$v4420%now\ <= (others => '0');
        \$19625%now\ <= (others => '0');
        \$v5576%now\ <= (others => '0');
        \$19886%now\ <= (others => '0');
        \$v5482%now\ <= (others => '0');
        \result4928%now\ <= (others => '0');
        \$19773%now\ <= (others => '0');
        \$v4424%now\ <= (others => '0');
        \$19787%now\ <= (others => '0');
        \$19104_modulo6684357_result%now\ <= (others => '0');
        \$v5769%now\ <= (others => '0');
        \$19496_aux664_result%now\ <= (others => '0');
        \$19717%now\ <= (others => '0');
        \$18647%now\ <= (others => '0');
        \$19155%now\ <= (others => '0');
        \$18661%now\ <= (others => '0');
        \$v4587%now\ <= (others => '0');
        \$19939%now\ <= (others => '0');
        \$18832_v%now\ <= (others => '0');
        \$19227%now\ <= (others => '0');
        \$19650%now\ <= (others => '0');
        \$18495%now\ <= (others => '0');
        \$18551%now\ <= (others => '0');
        \$v5658%now\ <= (others => '0');
        \$19276%now\ <= (others => '0');
        \$19859%now\ <= (others => '0');
        \$19325%now\ <= (others => '0');
        \$18977_binop_int6434365_result%now\ <= (others => '0');
        \$18944_r%now\ <= (others => '0');
        \$18527%now\ <= (others => '0');
        \$19119_v%now\ <= (others => '0');
        \$18648%now\ <= (others => '0');
        \$19793%now\ <= (others => '0');
        \$18877_v%now\ <= (others => '0');
        \$18939_binop_int6434363_id%now\ <= (others => '0');
        \$v5673%now\ <= (others => '0');
        \$19190_binop_compare6454380_id%now\ <= (others => '0');
        \$19842%now\ <= (others => '0');
        \$19144_modulo6684349_id%now\ <= (others => '0');
        \$v5536%now\ <= (others => '0');
        \$v5299%now\ <= (others => '0');
        \$19601_copy_root_in_ram6634352_arg%now\ <= (others => '0');
        \$18539%now\ <= (others => '0');
        \$18936_modulo6684349_id%now\ <= (others => '0');
        \$19015_binop_int6434367_result%now\ <= (others => '0');
        \$19171_compare6444358_id%now\ <= (others => '0');
        \$19597%now\ <= (others => '0');
        \$19581%now\ <= (others => '0');
        \$v4338%now\ <= (others => '0');
        \$19384_compare6444359_result%now\ <= (others => '0');
        \$19748%now\ <= (others => '0');
        \$18522_loop665_id%now\ <= (others => '0');
        \$18461%now\ <= (others => '0');
        \$19256_v%now\ <= (others => '0');
        \$v5206%now\ <= (others => '0');
        \$18824_v%now\ <= (others => '0');
        \$v5059%now\ <= (others => '0');
        \$18657%now\ <= (others => '0');
        \$v5026%now\ <= (others => '0');
        \$v4996%now\ <= (others => '0');
        \$v5036%now\ <= (others => '0');
        \$18825%now\ <= (others => '0');
        \$18806%now\ <= (others => '0');
        \$v4866%now\ <= (others => '0');
        \$v4647%now\ <= (others => '0');
        \$18891%now\ <= (others => '0');
        \$18843%now\ <= (others => '0');
        \$v4330%now\ <= (others => '0');
        \$19370_compare6444359_id%now\ <= (others => '0');
        \$19601_copy_root_in_ram6634352_id%now\ <= (others => '0');
        \$v5281%now\ <= (others => '0');
        \$v4546%now\ <= (others => '0');
        \$v4779%now\ <= (others => '0');
        \$v4636%now\ <= (others => '0');
        \$v4812%now\ <= (others => '0');
        \$v5574%now\ <= (others => '0');
        \$18526_aux664_arg%now\ <= (others => '0');
        \$19308_v%now\ <= (others => '0');
        \$18793_make_block579_arg%now\ <= (others => '0');
        \$18437_loop666_arg%now\ <= (others => '0');
        \$19206_binop_compare6454382_result%now\ <= (others => '0');
        \$18444%now\ <= (others => '0');
        \$19066_modulo6684357_id%now\ <= (others => '0');
        \$19046_r%now\ <= (others => '0');
        \$19837%now\ <= (others => '0');
        \$v5429%now\ <= (others => '0');
        \$19571%now\ <= (others => '0');
        \$v4978%now\ <= (others => '0');
        \$v4920%now\ <= (others => '0');
        \$v5799%now\ <= (others => '0');
        \$18524_loop666_arg%now\ <= (others => '0');
        \$18810%now\ <= (others => '0');
        \$19944%now\ <= (others => '0');
        \$18880%now\ <= (others => '0');
        \$18869%now\ <= (others => '0');
        \$v5490%now\ <= (others => '0');
        \$18659%now\ <= (others => '0');
        \$v5257%now\ <= (others => '0');
        \$18945_modulo6684356_id%now\ <= (others => '0');
        \$18683_hd%now\ <= (others => '0');
        \$v4428%now\ <= (others => '0');
        \$v5055%now\ <= (others => '0');
        \$19774%now\ <= (others => '0');
        \$v5522%now\ <= (others => '0');
        \$19783%now\ <= (others => '0');
        \$19125_modulo6684349_result%now\ <= (others => '0');
        \$19097_modulo6684356_id%now\ <= (others => '0');
        \$19507_next%now\ <= (others => '0');
        \rdy4400%now\ <= (others => '0');
        \$19542%now\ <= (others => '0');
        \$v5042%now\ <= (others => '0');
        \$18813%now\ <= (others => '0');
        \$19220%now\ <= (others => '0');
        \$v4667%now\ <= (others => '0');
        \$v4678%now\ <= (others => '0');
        \$19211_compare6444358_result%now\ <= (others => '0');
        \$18790_loop666_result%now\ <= (others => '0');
        \$19804%now\ <= (others => '0');
        \$18622%now\ <= (others => '0');
        \$v4519%now\ <= (others => '0');
        \$19667%now\ <= (others => '0');
        \$v4593%now\ <= (others => '0');
        \$19811_copy_root_in_ram6634341_arg%now\ <= (others => '0');
        \$18695%now\ <= (others => '0');
        \$19789_next%now\ <= (others => '0');
        \$19259%now\ <= (others => '0');
        \$18437_loop666_id%now\ <= (others => '0');
        \$19203_compare6444358_id%now\ <= (others => '0');
        \$19788%now\ <= (others => '0');
        \$19141_modulo6684356_arg%now\ <= (others => '0');
        \$18473%now\ <= (others => '0');
        \$v5134%now\ <= (others => '0');
        \$19144_modulo6684349_result%now\ <= (others => '0');
        \$19932%now\ <= (others => '0');
        \$18603%now\ <= (others => '0');
        \$v5365%now\ <= (others => '0');
        \$19701%now\ <= (others => '0');
        \$19543%now\ <= (others => '0');
        \$v5168%now\ <= (others => '0');
        \$v4529%now\ <= (others => '0');
        \$v4839%now\ <= (others => '0');
        \$v4679%now\ <= (others => '0');
        \$19796%now\ <= (others => '0');
        \$18845%now\ <= (others => '0');
        \$v5233%now\ <= (others => '0');
        \$18438_loop665_arg%now\ <= (others => '0');
        \$19337_compare6444359_arg%now\ <= (others => '0');
        \$v4632%now\ <= (others => '0');
        \$v4957%now\ <= (others => '0');
        \$19336_b%now\ <= (others => '0');
        \$19709%now\ <= (others => '0');
        \$19031_modulo6684349_result%now\ <= (others => '0');
        \$19824_hd%now\ <= (others => '0');
        \$19619%now\ <= (others => '0');
        \$18546%now\ <= (others => '0');
        \$v5872%now\ <= (others => '0');
        \$19818%now\ <= (others => '0');
        \$18971_modulo6684357_arg%now\ <= (others => '0');
        \$v4502%now\ <= (others => '0');
        \$19326_compbranch6504387_id%now\ <= (others => '0');
        \$18531%now\ <= (others => '0');
        \$v4802%now\ <= (others => '0');
        \$18841%now\ <= (others => '0');
        \$v4639%now\ <= (others => '0');
        \$19466_sp%now\ <= (others => '0');
        \$18567%now\ <= (others => '0');
        \$v4683%now\ <= (others => '0');
        \$19643_w%now\ <= (others => '0');
        \$18649%now\ <= (others => '0');
        \$18929_modulo6684349_arg%now\ <= (others => '0');
        \$v5184%now\ <= (others => '0');
        \$v4335%now\ <= (others => '0');
        \$v5915%now\ <= (others => '0');
        \$19169_v%now\ <= (others => '0');
        \$v5487%now\ <= (others => '0');
        \$v5552%now\ <= (others => '0');
        \$19361_fill6544390_id%now\ <= (others => '0');
        \$v5811%now\ <= (others => '0');
        \$19512%now\ <= (others => '0');
        \$v4471%now\ <= (others => '0');
        \$19725%now\ <= (others => '0');
        \$19844%now\ <= (others => '0');
        \$18732%now\ <= (others => '0');
        \$18618%now\ <= (others => '0');
        \$19387_compbranch6504394_arg%now\ <= (others => '0');
        \$19027_r%now\ <= (others => '0');
        \$v5471%now\ <= (others => '0');
        \$19659_hd%now\ <= (others => '0');
        \$19875%now\ <= (others => '0');
        \$19639%now\ <= (others => '0');
        \$18470%now\ <= (others => '0');
        \$19310%now\ <= (others => '0');
        \$19815%now\ <= (others => '0');
        \$v5696%now\ <= (others => '0');
        \$19350_v%now\ <= (others => '0');
        \$19503%now\ <= (others => '0');
        \$19182_binop_compare6454379_result%now\ <= (others => '0');
        \$18955_modulo6684349_result%now\ <= (others => '0');
        \$18476%now\ <= (others => '0');
        \$18443%now\ <= (others => '0');
        \$19230_v%now\ <= (others => '0');
        \$19018_v%now\ <= (others => '0');
        \$19713%now\ <= (others => '0');
        \$19218_v%now\ <= (others => '0');
        \$19009_modulo6684357_arg%now\ <= (others => '0');
        \$19498_loop665_result%now\ <= (others => '0');
        \$v5198%now\ <= (others => '0');
        \$19741%now\ <= (others => '0');
        \$v4581%now\ <= (others => '0');
        \$19161%now\ <= (others => '0');
        \$19156%now\ <= (others => '0');
        \$19104_modulo6684357_arg%now\ <= (others => '0');
        \$18492%now\ <= (others => '0');
        \$v5571%now\ <= (others => '0');
        \$v4615%now\ <= (others => '0');
        \$19937%now\ <= (others => '0');
        \$18917_modulo6684349_arg%now\ <= (others => '0');
        \$v5384%now\ <= (others => '0');
        \$18939_binop_int6434363_arg%now\ <= (others => '0');
        \$19572%now\ <= (others => '0');
        \$18898%now\ <= (others => '0');
        \$19391_compare6444359_result%now\ <= (others => '0');
        \$v5563%now\ <= (others => '0');
        \$18948_modulo6684349_id%now\ <= (others => '0');
        \$v5897%now\ <= (others => '0');
        \$19100_modulo6684349_id%now\ <= (others => '0');
        \$19409_sp%now\ <= (others => '0');
        \$18478%now\ <= (others => '0');
        \$19047_modulo6684357_result%now\ <= (others => '0');
        \$19009_modulo6684357_result%now\ <= (others => '0');
        \$v5072%now\ <= (others => '0');
        \$18895_v%now\ <= (others => '0');
        \$18559_copy_root_in_ram6634347_id%now\ <= (others => '0');
        \$18559_copy_root_in_ram6634347_arg%now\ <= (others => '0');
        \$19922%now\ <= (others => '0');
        \$19125_modulo6684349_id%now\ <= (others => '0');
        \$18629%now\ <= (others => '0');
        \$v4887%now\ <= (others => '0');
        \$v4556%now\ <= (others => '0');
        \$v5453%now\ <= (others => '0');
        \$19731%now\ <= (others => '0');
        \$19449%now\ <= (others => '0');
        \$18669%now\ <= (others => '0');
        \$18660%now\ <= (others => '0');
        \rdy4573%now\ <= (others => '0');
        \$18795_offsetclosure_n639_id%now\ <= (others => '0');
        \$19401_compbranch6504396_arg%now\ <= (others => '0');
        \$19878%now\ <= (others => '0');
        \$v5066%now\ <= (others => '0');
        \$18631%now\ <= (others => '0');
        \$v4327%now\ <= (others => '0');
        \$19234_sp%now\ <= (others => '0');
        \$18687%now\ <= (others => '0');
        \$19811_copy_root_in_ram6634341_result%now\ <= (others => '0');
        \rdy4608%now\ <= (others => '0');
        \$19728%now\ <= (others => '0');
        \$v5492%now\ <= (others => '0');
        \$19843%now\ <= (others => '0');
        \$19532_forever6704350_arg%now\ <= (others => '0');
        \$19028_modulo6684357_id%now\ <= (others => '0');
        \$18958_binop_int6434364_arg%now\ <= (others => '0');
        \$v4700%now\ <= (others => '0');
        \$19301_v%now\ <= (others => '0');
        \$v4940%now\ <= (others => '0');
        \$19012_modulo6684349_result%now\ <= (others => '0');
        \$19268%now\ <= (others => '0');
        \$19772%now\ <= (others => '0');
        \$19226%now\ <= (others => '0');
        \$v5727%now\ <= (others => '0');
        \$18889_v%now\ <= (others => '0');
        \$19882%now\ <= (others => '0');
        \$19877%now\ <= (others => '0');
        \$19091_binop_int6434371_id%now\ <= (others => '0');
        \$v4796%now\ <= (others => '0');
        \$18907_modulo6684356_result%now\ <= (others => '0');
        \$19561%now\ <= (others => '0');
        \$19282_v%now\ <= (others => '0');
        \$19806%now\ <= (others => '0');
        \$19257_v%now\ <= (others => '0');
        \$19660%now\ <= (others => '0');
        \$18583_w%now\ <= (others => '0');
        \$v4818%now\ <= (others => '0');
        \$v4750%now\ <= (others => '0');
        \$19492%now\ <= (others => '0');
        \$18525_loop665_id%now\ <= (others => '0');
        \$19311%now\ <= (others => '0');
        \$19743%now\ <= (others => '0');
        \$v4775%now\ <= (others => '0');
        \$v4713%now\ <= (others => '0');
        \$19519%now\ <= (others => '0');
        \$19870%now\ <= (others => '0');
        \$v4540%now\ <= (others => '0');
        \$19638%now\ <= (others => '0');
        \$v4821%now\ <= (others => '0');
        \$v5664%now\ <= (others => '0');
        \$19211_compare6444358_arg%now\ <= (others => '0');
        \$18500%now\ <= (others => '0');
        \$18545_next%now\ <= (others => '0');
        \$19078_modulo6684356_result%now\ <= (others => '0');
        \$19868%now\ <= (others => '0');
        \$19047_modulo6684357_id%now\ <= (others => '0');
        \$18663%now\ <= (others => '0');
        \$18679%now\ <= (others => '0');
        \$19053_binop_int6434369_result%now\ <= (others => '0');
        \$v4937%now\ <= (others => '0');
        \$v5305%now\ <= (others => '0');
        \$18986_modulo6684349_result%now\ <= (others => '0');
        \$19266%now\ <= (others => '0');
        \$19447_sp%now\ <= (others => '0');
        \$19084_r%now\ <= (others => '0');
        \$19779_loop666_result%now\ <= (others => '0');
        \$v5825%now\ <= (others => '0');
        \$18464_rdy%now\ <= (others => '0');
        \$19636%now\ <= (others => '0');
        \$19329_b%now\ <= (others => '0');
        \$v5596%now\ <= (others => '0');
        \$19031_modulo6684349_id%now\ <= (others => '0');
        \$19526_forever6704355_id%now\ <= (others => '0');
        \$19926%now\ <= (others => '0');
        \$19614_hd%now\ <= (others => '0');
        \$19594%now\ <= (others => '0');
        \$18542_next%now\ <= (others => '0');
        \$18553_forever6704348_id%now\ <= (others => '0');
        \$19521%now\ <= (others => '0');
        \$19832%now\ <= (others => '0');
        \$v4455%now\ <= (others => '0');
        \$v4640%now\ <= (others => '0');
        \$19053_binop_int6434369_arg%now\ <= (others => '0');
        \$18508%now\ <= (others => '0');
        \$19684%now\ <= (others => '0');
        \$19315%now\ <= (others => '0');
        \$19166_binop_compare6454377_id%now\ <= (others => '0');
        \$19110%now\ <= (others => '0');
        \$19678%now\ <= (others => '0');
        \$v5405%now\ <= (others => '0');
        \$v5622%now\ <= (others => '0');
        \$v5188%now\ <= (others => '0');
        \$v5138%now\ <= (others => '0');
        \$19198_binop_compare6454381_result%now\ <= (others => '0');
        \$v4972%now\ <= (others => '0');
        \$19872%now\ <= (others => '0');
        \$19031_modulo6684349_arg%now\ <= (others => '0');
        \$19405_compare6444359_arg%now\ <= (others => '0');
        \$v4754%now\ <= (others => '0');
        \$v5254%now\ <= (others => '0');
        \$v5275%now\ <= (others => '0');
        \$18642%now\ <= (others => '0');
        \$19892%now\ <= (others => '0');
        \$v4339%now\ <= (others => '0');
        \$v4532%now\ <= (others => '0');
        \$v5260%now\ <= (others => '0');
        \$19021_modulo6684356_arg%now\ <= (others => '0');
        \$18996_binop_int6434366_result%now\ <= (others => '0');
        \$19005_modulo6684349_id%now\ <= (others => '0');
        \$18522_loop665_result%now\ <= (others => '0');
        \$18682_w%now\ <= (others => '0');
        \$18914_modulo6684357_id%now\ <= (others => '0');
        \$18673%now\ <= (others => '0');
        \$19766%now\ <= (others => '0');
        \$v4558%now\ <= (others => '0');
        \$19214%now\ <= (others => '0');
        \$19566%now\ <= (others => '0');
        \$v4337%now\ <= (others => '0');
        \$v5096%now\ <= (others => '0');
        \$v5359%now\ <= (others => '0');
        \$19174_binop_compare6454378_result%now\ <= (others => '0');
        \$19563%now\ <= (others => '0');
        \$v4606%now\ <= (others => '0');
        \$v5141%now\ <= (others => '0');
        \$18639%now\ <= (others => '0');
        \$19154%now\ <= (others => '0');
        \$18562%now\ <= (others => '0');
        \$v4449%now\ <= (others => '0');
        \$v4605%now\ <= (others => '0');
        \$v4539%now\ <= (others => '0');
        \$18666%now\ <= (others => '0');
        \$19781_aux664_id%now\ <= (others => '0');
        \$18904_v%now\ <= (others => '0');
        \$18498%now\ <= (others => '0');
        \$v4562%now\ <= (others => '0');
        \$19497_loop666_arg%now\ <= (others => '0');
        \$18564%now\ <= (others => '0');
        \$v5335%now\ <= (others => '0');
        \$19834%now\ <= (others => '0');
        \$19700%now\ <= (others => '0');
        \$19769%now\ <= (others => '0');
        \$19907%now\ <= (others => '0');
        \$18724%now\ <= (others => '0');
        \$19425%now\ <= (others => '0');
        \$19293%now\ <= (others => '0');
        \$19147_r%now\ <= (others => '0');
        \$19950%now\ <= (others => '0');
        \$19355%now\ <= (others => '0');
        \$19024_modulo6684349_id%now\ <= (others => '0');
        \$19665%now\ <= (others => '0');
        \$19351%now\ <= (others => '0');
        \$19500%now\ <= (others => '0');
        \$v4833%now\ <= (others => '0');
        \$v4791%now\ <= (others => '0');
        \$v4746%now\ <= (others => '0');
        \$v5524%now\ <= (others => '0');
        \$19856%now\ <= (others => '0');
        \$18456%now\ <= (others => '0');
        \$19021_modulo6684356_result%now\ <= (others => '0');
        \$v5560%now\ <= (others => '0');
        \$v4751%now\ <= (others => '0');
        \$18487%now\ <= (others => '0');
        \$19755%now\ <= (others => '0');
        \$19233%now\ <= (others => '0');
        \$18654%now\ <= (others => '0');
        \$v4911%now\ <= (others => '0');
        \$v5743%now\ <= (others => '0');
        \$19414%now\ <= (others => '0');
        \$19649%now\ <= (others => '0');
        \$18702%now\ <= (others => '0');
        \$18897%now\ <= (others => '0');
        \$v4496%now\ <= (others => '0');
        \$18967_modulo6684349_result%now\ <= (others => '0');
        \$v5477%now\ <= (others => '0');
        \$v4675%now\ <= (others => '0');
        \$v5107%now\ <= (others => '0');
        \$19485%now\ <= (others => '0');
        \$v5597%now\ <= (others => '0');
        \$19132_modulo6684349_arg%now\ <= (others => '0');
        \$18781%now\ <= (others => '0');
        \$19252_forever6704384_id%now\ <= (others => '0');
        \$v4984%now\ <= (others => '0');
        \$v5753%now\ <= (others => '0');
        \$18896_v%now\ <= (others => '0');
        \$18737%now\ <= (others => '0');
        \$18439_wait662_result%now\ <= (others => '0');
        \$v5102%now\ <= (others => '0');
        \$v4813%now\ <= (others => '0');
        \$v5432%now\ <= (others => '0');
        \$19642%now\ <= (others => '0');
        \$18446_dur%now\ <= (others => '0');
        \$18625_copy_root_in_ram6634345_id%now\ <= (others => '0');
        \$v5314%now\ <= (others => '0');
        \$v5540%now\ <= (others => '0');
        \$19617%now\ <= (others => '0');
        \$19451%now\ <= (others => '0');
        \$18556_forever6704344_id%now\ <= (others => '0');
        \$19585%now\ <= (others => '0');
        \$18886%now\ <= (others => '0');
        \$18439_wait662_id%now\ <= (others => '0');
        \$v5441%now\ <= (others => '0');
        \$19737%now\ <= (others => '0');
        \$19879%now\ <= (others => '0');
        \$19072_binop_int6434370_id%now\ <= (others => '0');
        \$19462%now\ <= (others => '0');
        \$18516%now\ <= (others => '0');
        \$18838_v%now\ <= (others => '0');
        \$v5502%now\ <= (others => '0');
        \$v5814%now\ <= (others => '0');
        \$v5845%now\ <= (others => '0');
        \$18438_loop665_result%now\ <= (others => '0');
        \$19658_w%now\ <= (others => '0');
        \$19182_binop_compare6454379_arg%now\ <= (others => '0');
        \$18901_binop_int6434361_result%now\ <= (others => '0');
        \$18453%now\ <= (others => '0');
        \$19260%now\ <= (others => '0');
        \$v5605%now\ <= (others => '0');
        \$18971_modulo6684357_result%now\ <= (others => '0');
        \$19853%now\ <= (others => '0');
        \$v5131%now\ <= (others => '0');
        \$18820_v%now\ <= (others => '0');
        \$18571_copy_root_in_ram6634345_result%now\ <= (others => '0');
        \$18515%now\ <= (others => '0');
        \$v4689%now\ <= (others => '0');
        \$18914_modulo6684357_result%now\ <= (others => '0');
        \$v5497%now\ <= (others => '0');
        \$19951%now\ <= (others => '0');
        \$19807%now\ <= (others => '0');
        \$19241_v%now\ <= (others => '0');
        \$19242%now\ <= (others => '0');
        \$19539%now\ <= (others => '0');
        \$18752%now\ <= (others => '0');
        \$v5544%now\ <= (others => '0');
        \result4607%now\ <= (others => '0');
        \$19091_binop_int6434371_arg%now\ <= (others => '0');
        \$19345%now\ <= (others => '0');
        \$v5491%now\ <= (others => '0');
        \$18844%now\ <= (others => '0');
        \$18963_r%now\ <= (others => '0');
        \$v5652%now\ <= (others => '0');
        \$v5876%now\ <= (others => '0');
        \$19113_forever6704372_id%now\ <= (others => '0');
        \$19383_b%now\ <= (others => '0');
        \$19584%now\ <= (others => '0');
        \$19942%now\ <= (others => '0');
        \$19615%now\ <= (others => '0');
        \$18676%now\ <= (others => '0');
        \$v4514%now\ <= (others => '0');
        \$19316%now\ <= (others => '0');
        \$19148_modulo6684357_id%now\ <= (others => '0');
        \$v4492%now\ <= (others => '0');
        \$v5347%now\ <= (others => '0');
        \$v5411%now\ <= (others => '0');
        \$18756%now\ <= (others => '0');
        \$19865_w%now\ <= (others => '0');
        \$18533%now\ <= (others => '0');
        \$19297_v%now\ <= (others => '0');
        \$18497%now\ <= (others => '0');
        \$19062_modulo6684349_arg%now\ <= (others => '0');
        \$19456%now\ <= (others => '0');
        \$v5909%now\ <= (others => '0');
        \$v5356%now\ <= (others => '0');
        \$v5584%now\ <= (others => '0');
        \$v5023%now\ <= (others => '0');
        \$18766%now\ <= (others => '0');
        \$19770%now\ <= (others => '0');
        \$v4960%now\ <= (others => '0');
        \$18674%now\ <= (others => '0');
        \$18595%now\ <= (others => '0');
        \$19927%now\ <= (others => '0');
        \$v5293%now\ <= (others => '0');
        \$v5525%now\ <= (others => '0');
        \$18786%now\ <= (others => '0');
        \$19592%now\ <= (others => '0');
        \$18748%now\ <= (others => '0');
        \$18448_dis%now\ <= (others => '0');
        \$19398_compare6444359_result%now\ <= (others => '0');
        \$19202_res%now\ <= (others => '0');
        \$18951_r%now\ <= (others => '0');
        \$19040_modulo6684356_arg%now\ <= (others => '0');
        \$v5724%now\ <= (others => '0');
        \$18780%now\ <= (others => '0');
        \$18651%now\ <= (others => '0');
        \$19518_next%now\ <= (others => '0');
        \$19005_modulo6684349_result%now\ <= (others => '0');
        \$18808%now\ <= (others => '0');
        \$18715%now\ <= (others => '0');
        \$19799%now\ <= (others => '0');
        \$v5505%now\ <= (others => '0');
        \$v5867%now\ <= (others => '0');
        \$19646%now\ <= (others => '0');
        \$19833%now\ <= (others => '0');
        \$19182_binop_compare6454379_id%now\ <= (others => '0');
        \$v5000%now\ <= (others => '0');
        \$v5185%now\ <= (others => '0');
        \$v5034%now\ <= (others => '0');
        \$18467_loop665_result%now\ <= (others => '0');
        \$v5222%now\ <= (others => '0');
        \$v4782%now\ <= (others => '0');
        \$19547_copy_root_in_ram6634352_id%now\ <= (others => '0');
        \$19915%now\ <= (others => '0');
        \$19719%now\ <= (others => '0');
        \$18777%now\ <= (others => '0');
        \$18550%now\ <= (others => '0');
        \$18842%now\ <= (others => '0');
        \$18489%now\ <= (others => '0');
        \$18439_wait662_arg%now\ <= (others => '0');
        \$19100_modulo6684349_result%now\ <= (others => '0');
        \$19135_binop_int6434374_id%now\ <= (others => '0');
        \$18796_make_block_n646_arg%now\ <= (others => '0');
        \$v5084%now\ <= (others => '0');
        \$v4654%now\ <= (others => '0');
        \$19820%now\ <= (others => '0');
        \$18901_binop_int6434361_arg%now\ <= (others => '0');
        \$18701%now\ <= (others => '0');
        \$18768_w%now\ <= (others => '0');
        \$19586%now\ <= (others => '0');
        \$v5709%now\ <= (others => '0');
        \$18613_copy_root_in_ram6634346_arg%now\ <= (others => '0');
        \$19917%now\ <= (others => '0');
        \$19138_v%now\ <= (others => '0');
        \$19697%now\ <= (others => '0');
        \$v4423%now\ <= (others => '0');
        \result4963%now\ <= (others => '0');
        \$18794_apply638_arg%now\ <= (others => '0');
        \$18792_wait662_arg%now\ <= (others => '0');
        \$18741%now\ <= (others => '0');
        \$18735%now\ <= (others => '0');
        \$v5039%now\ <= (others => '0');
        \$19677%now\ <= (others => '0');
        \$v5296%now\ <= (others => '0');
        \$18714%now\ <= (others => '0');
        \$19231%now\ <= (others => '0');
        \$v5689%now\ <= (others => '0');
        \$v5251%now\ <= (others => '0');
        \$19876%now\ <= (others => '0');
        \$v5606%now\ <= (others => '0');
        \$v5670%now\ <= (others => '0');
        \$18794_apply638_result%now\ <= (others => '0');
        \$19921%now\ <= (others => '0');
        \$19420_w06554397_id%now\ <= (others => '0');
        \$v4719%now\ <= (others => '0');
        \$19059_modulo6684356_id%now\ <= (others => '0');
        \$19864%now\ <= (others => '0');
        \$19347_fill6534389_result%now\ <= (others => '0');
        \$v5099%now\ <= (others => '0');
        \$19860%now\ <= (others => '0');
        \$19781_aux664_arg%now\ <= (others => '0');
        \$v4827%now\ <= (others => '0');
        \$18964_modulo6684356_arg%now\ <= (others => '0');
        \$v5802%now\ <= (others => '0');
        \$v4917%now\ <= (others => '0');
        \$19302%now\ <= (others => '0');
        \$v5368%now\ <= (others => '0');
        \$19823_w%now\ <= (others => '0');
        \$v5494%now\ <= (others => '0');
        \$19668%now\ <= (others => '0');
        \$19398_compare6444359_id%now\ <= (others => '0');
        \$18574%now\ <= (others => '0');
        \$19228_v%now\ <= (others => '0');
        \$v5079%now\ <= (others => '0');
        \$19749%now\ <= (others => '0');
        \$19795%now\ <= (others => '0');
        \$19203_compare6444358_arg%now\ <= (others => '0');
        \$19768%now\ <= (others => '0');
        \$v4809%now\ <= (others => '0');
        \$19941%now\ <= (others => '0');
        \$v4902%now\ <= (others => '0');
        \$18899%now\ <= (others => '0');
        \$19605%now\ <= (others => '0');
        \$19514%now\ <= (others => '0');
        \$v4836%now\ <= (others => '0');
        \$18640%now\ <= (others => '0');
        \$v4716%now\ <= (others => '0');
        \$v5396%now\ <= (others => '0');
        \$19341%now\ <= (others => '0');
        \$18870_v%now\ <= (others => '0');
        \$19722%now\ <= (others => '0');
        \$19475%now\ <= (others => '0');
        \$v5353%now\ <= (others => '0');
        \$v4953%now\ <= (others => '0');
        \$19460%now\ <= (others => '0');
        \$19470%now\ <= (others => '0');
        \$19580%now\ <= (others => '0');
        \$19893%now\ <= (others => '0');
        \$v4597%now\ <= (others => '0');
        \$v5051%now\ <= (others => '0');
        \$v5679%now\ <= (others => '0');
        \$v5630%now\ <= (others => '0');
        \$19889%now\ <= (others => '0');
        \$18812%now\ <= (others => '0');
        \$v5543%now\ <= (others => '0');
        \$18955_modulo6684349_id%now\ <= (others => '0');
        \$19529_forever6704351_arg%now\ <= (others => '0');
        \$v5556%now\ <= (others => '0');
        \$19497_loop666_result%now\ <= (others => '0');
        \$18536%now\ <= (others => '0');
        \$19433%now\ <= (others => '0');
        \$v4857%now\ <= (others => '0');
        \$19286%now\ <= (others => '0');
        \$19621%now\ <= (others => '0');
        \$18758%now\ <= (others => '0');
        \$19261%now\ <= (others => '0');
        \$v5566%now\ <= (others => '0');
        \$v4881%now\ <= (others => '0');
        \$19148_modulo6684357_result%now\ <= (others => '0');
        \$v4795%now\ <= (others => '0');
        \$19945%now\ <= (others => '0');
        \$v4466%now\ <= (others => '0');
        \$v4824%now\ <= (others => '0');
        \$19747%now\ <= (others => '0');
        \$19081_modulo6684349_id%now\ <= (others => '0');
        \$19285%now\ <= (others => '0');
        \$v4884%now\ <= (others => '0');
        \$v5863%now\ <= (others => '0');
        \$19394_compbranch6504395_result%now\ <= (others => '0');
        \$19535_copy_root_in_ram6634354_result%now\ <= (others => '0');
        \$v4758%now\ <= (others => '0');
        \$v4488%now\ <= (others => '0');
        \$19012_modulo6684349_arg%now\ <= (others => '0');
        \$18607%now\ <= (others => '0');
        \$19753%now\ <= (others => '0');
        \$18785%now\ <= (others => '0');
        \$19394_compbranch6504395_id%now\ <= (others => '0');
        \$v5894%now\ <= (others => '0');
        \$18799_w1656_arg%now\ <= (others => '0');
        \$18856_loop_push6494360_id%now\ <= (others => '0');
        \$v4981%now\ <= (others => '0');
        \$19391_compare6444359_arg%now\ <= (others => '0');
        \$19366_compbranch6504391_id%now\ <= (others => '0');
        \$v4771%now\ <= (others => '0');
        \$19781_aux664_result%now\ <= (others => '0');
        \$19174_binop_compare6454378_id%now\ <= (others => '0');
        \$19416_w36574398_arg%now\ <= (others => '0');
        \$v5627%now\ <= (others => '0');
        \$19271%now\ <= (others => '0');
        \$v5126%now\ <= (others => '0');
        \$18708%now\ <= (others => '0');
        \$19780_loop665_id%now\ <= (others => '0');
        \$18827%now\ <= (others => '0');
        \$v5890%now\ <= (others => '0');
        \$18882_v%now\ <= (others => '0');
        \$18525_loop665_arg%now\ <= (others => '0');
        \$v5623%now\ <= (others => '0');
        \$19344%now\ <= (others => '0');
        \$19576%now\ <= (others => '0');
        \$19171_compare6444358_arg%now\ <= (others => '0');
        \$19838_copy_root_in_ram6634340_id%now\ <= (others => '0');
        \$v5387%now\ <= (others => '0');
        \$19373_compbranch6504392_arg%now\ <= (others => '0');
        \$v5602%now\ <= (others => '0');
        \$18544%now\ <= (others => '0');
        \$v5773%now\ <= (others => '0');
        \$18493%now\ <= (others => '0');
        \$18579%now\ <= (others => '0');
        \$v5444%now\ <= (others => '0');
        \$19524%now\ <= (others => '0');
        \$19247%now\ <= (others => '0');
        \$19122_modulo6684356_id%now\ <= (others => '0');
        \$v5585%now\ <= (others => '0');
        \$19494_loop666_result%now\ <= (others => '0');
        \$19284%now\ <= (others => '0');
        \$19373_compbranch6504392_id%now\ <= (others => '0');
        \$19287_v%now\ <= (others => '0');
        \$19808_forever6704342_id%now\ <= (others => '0');
        \$v5459%now\ <= (others => '0');
        \$19767%now\ <= (others => '0');
        \$v5181%now\ <= (others => '0');
        \$19494_loop666_id%now\ <= (others => '0');
        \$19529_forever6704351_id%now\ <= (others => '0');
        \$v5782%now\ <= (others => '0');
        \$19053_binop_int6434369_id%now\ <= (others => '0');
        \$v4478%now\ <= (others => '0');
        \$v5495%now\ <= (others => '0');
        \$v4505%now\ <= (others => '0');
        \$18621%now\ <= (others => '0');
        \$19598%now\ <= (others => '0');
        \$v4774%now\ <= (others => '0');
        \$18523_aux664_result%now\ <= (others => '0');
        \$v5919%now\ <= (others => '0');
        \$19298_v%now\ <= (others => '0');
        \$18872_v%now\ <= (others => '0');
        \$18817_v%now\ <= (others => '0');
        \$19762%now\ <= (others => '0');
        \$19002_modulo6684356_id%now\ <= (others => '0');
        \$v5695%now\ <= (others => '0');
        \$v5770%now\ <= (others => '0');
        \$19024_modulo6684349_arg%now\ <= (others => '0');
        \$18936_modulo6684349_result%now\ <= (others => '0');
        \$19428%now\ <= (others => '0');
        \$18890_v%now\ <= (others => '0');
        \$v5561%now\ <= (others => '0');
        \$18535%now\ <= (others => '0');
        \$19151_modulo6684349_arg%now\ <= (others => '0');
        \result4399%now\ <= (others => '0');
        \$19278%now\ <= (others => '0');
        \rdy4435%now\ <= (others => '0');
        \$19000_res%now\ <= (others => '0');
        \$18609%now\ <= (others => '0');
        \$18720%now\ <= (others => '0');
        \$19552%now\ <= (others => '0');
        \$18757%now\ <= (others => '0');
        \$v4459%now\ <= (others => '0');
        \$19305%now\ <= (others => '0');
        \$18874%now\ <= (others => '0');
        \$18800%now\ <= (others => '0');
        \$19607%now\ <= (others => '0');
        \$v4557%now\ <= (others => '0');
        \$19757%now\ <= (others => '0');
        \$v4536%now\ <= (others => '0');
        \$19933_w%now\ <= (others => '0');
        \$v4487%now\ <= (others => '0');
        \$19258%now\ <= (others => '0');
        \$v4720%now\ <= (others => '0');
        \$19151_modulo6684349_id%now\ <= (others => '0');
        \$19744_w%now\ <= (others => '0');
        \result4572%now\ <= (others => '0');
        \$19103_r%now\ <= (others => '0');
        \$v5562%now\ <= (others => '0');
        \$19178_res%now\ <= (others => '0');
        \$19160%now\ <= (others => '0');
        \$19663%now\ <= (others => '0');
        \$18871%now\ <= (others => '0');
        \$v5332%now\ <= (others => '0');
        \$v5045%now\ <= (others => '0');
        \$19193_v%now\ <= (others => '0');
        \$v4670%now\ <= (others => '0');
        \$v5880%now\ <= (others => '0');
        \$v5030%now\ <= (others => '0');
        \$18883_v%now\ <= (others => '0');
        \$v4333%now\ <= (others => '0');
        \$v5572%now\ <= (others => '0');
        \$18983_modulo6684356_result%now\ <= (others => '0');
        \$19493%now\ <= (others => '0');
        \$19095_res%now\ <= (others => '0');
        \$v5756%now\ <= (others => '0');
        \$18983_modulo6684356_arg%now\ <= (others => '0');
        \$v5114%now\ <= (others => '0');
        \$v5192%now\ <= (others => '0');
        \$19461%now\ <= (others => '0');
        \$19107_modulo6684349_result%now\ <= (others => '0');
        \$18839%now\ <= (others => '0');
        \$v5341%now\ <= (others => '0');
        \$v5626%now\ <= (others => '0');
        \$19050_modulo6684349_id%now\ <= (others => '0');
        \$18787%now\ <= (others => '0');
        \$18716%now\ <= (others => '0');
        \$19121_r%now\ <= (others => '0');
        \$19206_binop_compare6454382_id%now\ <= (others => '0');
        \$18885_v%now\ <= (others => '0');
        \$18658%now\ <= (others => '0');
        \$v5851%now\ <= (others => '0');
        \$19069_modulo6684349_result%now\ <= (others => '0');
        \$v5111%now\ <= (others => '0');
        \$18678%now\ <= (others => '0');
        \$19822%now\ <= (others => '0');
        \$v5510%now\ <= (others => '0');
        \$18753%now\ <= (others => '0');
        \$v5848%now\ <= (others => '0');
        \$19113_forever6704372_arg%now\ <= (others => '0');
        \$18840_v%now\ <= (others => '0');
        \$v5362%now\ <= (others => '0');
        \$v4905%now\ <= (others => '0');
        \$18596%now\ <= (others => '0');
        \$v4553%now\ <= (others => '0');
        \$v5218%now\ <= (others => '0');
        \$18440_make_block579_result%now\ <= (others => '0');
        \$19401_compbranch6504396_id%now\ <= (others => '0');
        \$19380_compbranch6504393_result%now\ <= (others => '0');
        \$19047_modulo6684357_arg%now\ <= (others => '0');
        \$18861%now\ <= (others => '0');
        \$19931%now\ <= (others => '0');
        \$19340_argument2%now\ <= (others => '0');
        \$v4991%now\ <= (others => '0');
        \$18983_modulo6684356_id%now\ <= (others => '0');
        \$v5591%now\ <= (others => '0');
        \$v5211%now\ <= (others => '0');
        \$18920_binop_int6434362_id%now\ <= (others => '0');
        \$v5531%now\ <= (others => '0');
        \$19002_modulo6684356_result%now\ <= (others => '0');
        \$v4890%now\ <= (others => '0');
        \$18589%now\ <= (others => '0');
        \$19144_modulo6684349_arg%now\ <= (others => '0');
        \$v4600%now\ <= (others => '0');
        \$19476_v%now\ <= (others => '0');
        \$19587%now\ <= (others => '0');
        \$19919%now\ <= (others => '0');
        \$19574_w%now\ <= (others => '0');
        \$19237_v%now\ <= (others => '0');
        \$19037_v%now\ <= (others => '0');
        \$v5483%now\ <= (others => '0');
        \$19634%now\ <= (others => '0');
        \$18585%now\ <= (others => '0');
        \$v4432%now\ <= (others => '0');
        \$19365%now\ <= (others => '0');
        \$v5736%now\ <= (others => '0');
        \$v4332%now\ <= (others => '0');
        \$19857%now\ <= (others => '0');
        \$v5868%now\ <= (others => '0');
        \$18803%now\ <= (others => '0');
        \$19346_sp%now\ <= (others => '0');
        \$18691%now\ <= (others => '0');
        \$19846%now\ <= (others => '0');
        \$v5841%now\ <= (others => '0');
        \$19695%now\ <= (others => '0');
        \$19494_loop666_arg%now\ <= (others => '0');
        \$v5177%now\ <= (others => '0');
        \$v4707%now\ <= (others => '0');
        \$19122_modulo6684356_arg%now\ <= (others => '0');
        \$v4737%now\ <= (others => '0');
        \$v5712%now\ <= (others => '0');
        \$19370_compare6444359_arg%now\ <= (others => '0');
        \$19622%now\ <= (others => '0');
        \$v4567%now\ <= (others => '0');
        \$v5500%now\ <= (others => '0');
        \$19899%now\ <= (others => '0');
        \$v5918%now\ <= (others => '0');
        \$v5408%now\ <= (others => '0');
        \$19039_r%now\ <= (others => '0');
        \$18814%now\ <= (others => '0');
        \$19738%now\ <= (others => '0');
        \$19670%now\ <= (others => '0');
        \$19457%now\ <= (others => '0');
        \$19377_compare6444359_id%now\ <= (others => '0');
        \$19556%now\ <= (others => '0');
        \$19711%now\ <= (others => '0');
        \$v5808%now\ <= (others => '0');
        \$19377_compare6444359_arg%now\ <= (others => '0');
        \$19405_compare6444359_result%now\ <= (others => '0');
        \$v5593%now\ <= (others => '0');
        \$19903_next%now\ <= (others => '0');
        \$18818_v%now\ <= (others => '0');
        \$18633%now\ <= (others => '0');
        \$18466_loop666_arg%now\ <= (others => '0');
        \$19459%now\ <= (others => '0');
        \$19705%now\ <= (others => '0');
        \$19629_hd%now\ <= (others => '0');
        \$18836_v%now\ <= (others => '0');
        \$19384_compare6444359_arg%now\ <= (others => '0');
        \$18736%now\ <= (others => '0');
        \$v5110%now\ <= (others => '0');
        \$18671%now\ <= (others => '0');
        \$18686%now\ <= (others => '0');
        \$v4526%now\ <= (others => '0');
        \$18990_modulo6684357_arg%now\ <= (others => '0');
        \$v5493%now\ <= (others => '0');
        \$19632%now\ <= (others => '0');
        \$v5871%now\ <= (others => '0');
        \$18823_v%now\ <= (others => '0');
        \$18593%now\ <= (others => '0');
        \$v5229%now\ <= (others => '0');
        \$v5302%now\ <= (others => '0');
        \$18652_w%now\ <= (others => '0');
        \$19506%now\ <= (others => '0');
        \$19337_compare6444359_result%now\ <= (others => '0');
        \$v4411%now\ <= (others => '0');
        \$19680%now\ <= (others => '0');
        \rdy4964%now\ <= (others => '0');
        \$18690%now\ <= (others => '0');
        \$v4755%now\ <= (others => '0');
        \$v5615%now\ <= (others => '0');
        \$19195_compare6444358_id%now\ <= (others => '0');
        \$19912%now\ <= (others => '0');
        \$18469_make_block579_arg%now\ <= (others => '0');
        \$18743%now\ <= (others => '0');
        \$19791%now\ <= (others => '0');
        \$19604%now\ <= (others => '0');
        \$v5805%now\ <= (others => '0');
        \$19510%now\ <= (others => '0');
        \$18728%now\ <= (others => '0');
        \$19869%now\ <= (others => '0');
        \$19900%now\ <= (others => '0');
        \$19898%now\ <= (others => '0');
        \$19111%now\ <= (others => '0');
        \$18586%now\ <= (others => '0');
        \$18986_modulo6684349_id%now\ <= (others => '0');
        \$18468_wait662_id%now\ <= (others => '0');
        \$19244_v%now\ <= (others => '0');
        \$19612%now\ <= (others => '0');
        \$v4785%now\ <= (others => '0');
        \$19847%now\ <= (others => '0');
        \$19398_compare6444359_arg%now\ <= (others => '0');
        \$v4987%now\ <= (others => '0');
        \$19830%now\ <= (others => '0');
        \$19034_binop_int6434368_id%now\ <= (others => '0');
        \$18856_loop_push6494360_result%now\ <= (others => '0');
        \$19687_w%now\ <= (others => '0');
        \$19745_hd%now\ <= (others => '0');
        \$18894_v%now\ <= (others => '0');
        \$v5887%now\ <= (others => '0');
        \$18672%now\ <= (others => '0');
        \$18617%now\ <= (others => '0');
        \$19938%now\ <= (others => '0');
        \$18892_v%now\ <= (others => '0');
        \$19437%now\ <= (others => '0');
        \$18636%now\ <= (others => '0');
        \$18611%now\ <= (others => '0');
        \$19225%now\ <= (others => '0');
        \$19420_w06554397_arg%now\ <= (others => '0');
        \$18713%now\ <= (others => '0');
        \$18616%now\ <= (others => '0');
        \$18771%now\ <= (others => '0');
        \$v4635%now\ <= (others => '0');
        \$v5792%now\ <= (others => '0');
        \$18868_v%now\ <= (others => '0');
        \$v5106%now\ <= (others => '0');
        \$18693%now\ <= (others => '0');
        \$18597%now\ <= (others => '0');
        \$18437_loop666_result%now\ <= (others => '0');
        \$19426%now\ <= (others => '0');
        \$19763%now\ <= (others => '0');
        \$v5575%now\ <= (others => '0');
        \$v4747%now\ <= (others => '0');
        \$v5381%now\ <= (others => '0');
        \$19151_modulo6684349_result%now\ <= (others => '0');
        \$v5474%now\ <= (others => '0');
        \$18850%now\ <= (others => '0');
        \$18445_x%now\ <= (others => '0');
        \$18798_w652_arg%now\ <= (others => '0');
        \$18878%now\ <= (others => '0');
        \$v5820%now\ <= (others => '0');
        \$v5022%now\ <= (others => '0');
        \$v4968%now\ <= (others => '0');
        \$v4686%now\ <= (others => '0');
        \$19472%now\ <= (others => '0');
        \$v5718%now\ <= (others => '0');
        \$19404_b%now\ <= (others => '0');
        \$v4446%now\ <= (others => '0');
        \$19624%now\ <= (others => '0');
        \$18587%now\ <= (others => '0');
        \$v5906%now\ <= (others => '0');
        \$18970_r%now\ <= (others => '0');
        \$19545%now\ <= (others => '0');
        \$18534_next%now\ <= (others => '0');
        \$19219%now\ <= (others => '0');
        \$18792_wait662_id%now\ <= (others => '0');
        \$19265_ofs%now\ <= (others => '0');
        \$19618%now\ <= (others => '0');
        \$19411%now\ <= (others => '0');
        \$19468_sp%now\ <= (others => '0');
        \$18547%now\ <= (others => '0');
        \$19116_binop_int6434373_id%now\ <= (others => '0');
        \$19065_r%now\ <= (others => '0');
        \$19645%now\ <= (others => '0');
        \$19129_modulo6684357_result%now\ <= (others => '0');
        \$v5155%now\ <= (others => '0');
        \$v5219%now\ <= (others => '0');
        \$19756%now\ <= (others => '0');
        \$18490%now\ <= (others => '0');
        \$18523_aux664_arg%now\ <= (others => '0');
        \$v5375%now\ <= (others => '0');
        \$19215_argument1%now\ <= (others => '0');
        \$18860%now\ <= (others => '0');
        \$v5898%now\ <= (others => '0');
        \$v4643%now\ <= (others => '0');
        \$19174_binop_compare6454378_arg%now\ <= (others => '0');
        \$v5581%now\ <= (others => '0');
        \$v4999%now\ <= (others => '0');
        \$18466_loop666_result%now\ <= (others => '0');
        \$18469_make_block579_result%now\ <= (others => '0');
        \$18625_copy_root_in_ram6634345_result%now\ <= (others => '0');
        \$19640%now\ <= (others => '0');
        \$v4657%now\ <= (others => '0');
        \$v5501%now\ <= (others => '0');
        \$19323%now\ <= (others => '0');
        \$v5631%now\ <= (others => '0');
        \$19270%now\ <= (others => '0');
        \$19473%now\ <= (others => '0');
        \$19318%now\ <= (others => '0');
        \$19132_modulo6684349_result%now\ <= (others => '0');
        \$18548%now\ <= (others => '0');
        \$18967_modulo6684349_id%now\ <= (others => '0');
        \$18772%now\ <= (others => '0');
        \$18628%now\ <= (others => '0');
        \$19562%now\ <= (others => '0');
        \$18538%now\ <= (others => '0');
        \$18819_v%now\ <= (others => '0');
        \$19198_binop_compare6454381_arg%now\ <= (others => '0');
        \$19465_sp%now\ <= (others => '0');
        \$18526_aux664_result%now\ <= (others => '0');
        \$19911%now\ <= (others => '0');
        \$v4914%now\ <= (others => '0');
        \$19446_sp%now\ <= (others => '0');
        \$18932_r%now\ <= (others => '0');
        \$v4463%now\ <= (others => '0');
        \$19946%now\ <= (others => '0');
        \$19943%now\ <= (others => '0');
        \$v5372%now\ <= (others => '0');
        \$19577%now\ <= (others => '0');
        \$18641%now\ <= (others => '0');
        \$18773%now\ <= (others => '0');
        \$v5740%now\ <= (others => '0');
        \$18524_loop666_id%now\ <= (others => '0');
        \$18964_modulo6684356_result%now\ <= (others => '0');
        \$v4427%now\ <= (others => '0');
        \$19655%now\ <= (others => '0');
        \$19028_modulo6684357_arg%now\ <= (others => '0');
        \$v4788%now\ <= (others => '0');
        \$19520%now\ <= (others => '0');
        \$v4875%now\ <= (others => '0');
        \$19306_v%now\ <= (others => '0');
        \$v5567%now\ <= (others => '0');
        \$v5521%now\ <= (others => '0');
        \$v4644%now\ <= (others => '0');
        \$19343_sp%now\ <= (others => '0');
        \$18722%now\ <= (others => '0');
        \$19935%now\ <= (others => '0');
        \$19056_v%now\ <= (others => '0');
        \$18513%now\ <= (others => '0');
        \$18989_r%now\ <= (others => '0');
        \$18879_v%now\ <= (others => '0');
        \$v4956%now\ <= (others => '0');
        \$19730%now\ <= (others => '0');
        \$18665%now\ <= (others => '0');
        \$v4452%now\ <= (others => '0');
        \$v5783%now\ <= (others => '0');
        \$18710%now\ <= (others => '0');
        \$v5676%now\ <= (others => '0');
        \$19009_modulo6684357_id%now\ <= (others => '0');
        \$19712%now\ <= (others => '0');
        \$19841%now\ <= (others => '0');
        \$18556_forever6704344_arg%now\ <= (others => '0');
        \$19780_loop665_result%now\ <= (others => '0');
        \$19236_v%now\ <= (others => '0');
        \$19330_compare6444359_result%now\ <= (others => '0');
        \$v5600%now\ <= (others => '0');
        \$19330_compare6444359_arg%now\ <= (others => '0');
        \$18592%now\ <= (others => '0');
        \$19289%now\ <= (others => '0');
        \$19589_copy_root_in_ram6634353_arg%now\ <= (others => '0');
        \$v4778%now\ <= (others => '0');
        \$19356%now\ <= (others => '0');
        \$19050_modulo6684349_arg%now\ <= (others => '0');
        \$v5241%now\ <= (others => '0');
        \$18594%now\ <= (others => '0');
        \$v5680%now\ <= (others => '0');
        \$18866_v%now\ <= (others => '0');
        \$v5877%now\ <= (others => '0');
        \$19424%now\ <= (others => '0');
        \$v5587%now\ <= (others => '0');
        \$19369_b%now\ <= (others => '0');
        \$18481%now\ <= (others => '0');
        \$19050_modulo6684349_result%now\ <= (others => '0');
        \$19691%now\ <= (others => '0');
        \$18471%now\ <= (others => '0');
        \$19058_r%now\ <= (others => '0');
        \$19560_hd%now\ <= (others => '0');
        \$19405_compare6444359_id%now\ <= (others => '0');
        \$v5901%now\ <= (others => '0');
        \$v5435%now\ <= (others => '0');
        \$19353%now\ <= (others => '0');
        \$19059_modulo6684356_result%now\ <= (others => '0');
        \$18910_modulo6684349_arg%now\ <= (others => '0');
        \$v5706%now\ <= (others => '0');
        \$18486%now\ <= (others => '0');
        \$18501%now\ <= (others => '0');
        \$18532%now\ <= (others => '0');
        \$v4764%now\ <= (others => '0');
        \$19216_v%now\ <= (others => '0');
        \$19613_w%now\ <= (others => '0');
        \$18528%now\ <= (others => '0');
        \$19283%now\ <= (others => '0');
        \$v5338%now\ <= (others => '0');
        \$19091_binop_int6434371_result%now\ <= (others => '0');
        \$v4962%now\ <= (others => '0');
        \$19654%now\ <= (others => '0');
        \$v5842%now\ <= (others => '0');
        \$v5527%now\ <= (others => '0');
        \$18920_binop_int6434362_result%now\ <= (others => '0');
        \$19195_compare6444358_arg%now\ <= (others => '0');
        \$v5910%now\ <= (others => '0');
        \$18705_next%now\ <= (others => '0');
        \$19511%now\ <= (others => '0');
        \$v5902%now\ <= (others => '0');
        \$19410%now\ <= (others => '0');
        \$18468_wait662_arg%now\ <= (others => '0');
        \$v5504%now\ <= (others => '0');
        \$v4522%now\ <= (others => '0');
        \$18797_branch_if648_arg%now\ <= (others => '0');
        \$19696%now\ <= (others => '0');
        \$18955_modulo6684349_arg%now\ <= (others => '0');
        \$19652%now\ <= (others => '0');
        \$19606%now\ <= (others => '0');
        \$19195_compare6444358_result%now\ <= (others => '0');
        \$v5006%now\ <= (others => '0');
        \$18804%now\ <= (others => '0');
        \$18910_modulo6684349_result%now\ <= (others => '0');
        \$19502%now\ <= (others => '0');
        \$v5583%now\ <= (others => '0');
        \$18853_hd%now\ <= (others => '0');
        \$v5746%now\ <= (others => '0');
        \$v5048%now\ <= (others => '0');
        \$19831%now\ <= (others => '0');
        \$19481%now\ <= (others => '0');
        \$18774%now\ <= (others => '0');
        \$19708%now\ <= (others => '0');
        \$18632%now\ <= (others => '0');
        \$18625_copy_root_in_ram6634345_arg%now\ <= (others => '0');
        \$v5834%now\ <= (others => '0');
        \$19568%now\ <= (others => '0');
        \$v4723%now\ <= (others => '0');
        \$18519%now\ <= (others => '0');
        \$v4580%now\ <= (others => '0');
        \$19547_copy_root_in_ram6634352_arg%now\ <= (others => '0');
        \$19477_v%now\ <= (others => '0');
        \$18704%now\ <= (others => '0');
        \$18503%now\ <= (others => '0');
        \$18790_loop666_arg%now\ <= (others => '0');
        \$v5854%now\ <= (others => '0');
        \$19690%now\ <= (others => '0');
        \$v5786%now\ <= (others => '0');
        \$19498_loop665_id%now\ <= (others => '0');
        \$v5864%now\ <= (others => '0');
        \$v5886%now\ <= (others => '0');
        \$18923_v%now\ <= (others => '0');
        \$v5914%now\ <= (others => '0');
        \$v5798%now\ <= (others => '0');
        \$v5016%now\ <= (others => '0');
        \$19499_aux664_result%now\ <= (others => '0');
        \$v5554%now\ <= (others => '0');
        \$18675%now\ <= (others => '0');
        \$18463%now\ <= (others => '0');
        \$19469%now\ <= (others => '0');
        \$18700%now\ <= (others => '0');
        \$18744_w%now\ <= (others => '0');
        \$v5087%now\ <= (others => '0');
        \$18530%now\ <= (others => '0');
        \$v5423%now\ <= (others => '0');
        \$v5215%now\ <= (others => '0');
        \$18929_modulo6684349_result%now\ <= (others => '0');
        \$19733%now\ <= (others => '0');
        \$18653_hd%now\ <= (others => '0');
        \$19429%now\ <= (others => '0');
        \$18833%now\ <= (others => '0');
        \$v5165%now\ <= (others => '0');
        \$18454%now\ <= (others => '0');
        \$18847%now\ <= (others => '0');
        \$v5553%now\ <= (others => '0');
        \$v5075%now\ <= (others => '0');
        \$18692%now\ <= (others => '0');
        \$18719%now\ <= (others => '0');
        \$19940%now\ <= (others => '0');
        \$18712_hd%now\ <= (others => '0');
        \$v5417%now\ <= (others => '0');
        \$19125_modulo6684349_arg%now\ <= (others => '0');
        \$18634%now\ <= (others => '0');
        \$19484%now\ <= (others => '0');
        \$18929_modulo6684349_id%now\ <= (others => '0');
        \$19198_binop_compare6454381_id%now\ <= (others => '0');
        \$19416_w36574398_id%now\ <= (others => '0');
        \$18798_w652_id%now\ <= (others => '0');
        \$v5056%now\ <= (others => '0');
        \$v4439%now\ <= (others => '0');
        \$v5503%now\ <= (others => '0');
        \$19608%now\ <= (others => '0');
        \$v5779%now\ <= (others => '0');
        \$19277%now\ <= (others => '0');
        \$19223%now\ <= (others => '0');
        \$18499%now\ <= (others => '0');
        \$18796_make_block_n646_result%now\ <= (others => '0');
        \$19085_modulo6684357_id%now\ <= (others => '0');
        \$v5399%now\ <= (others => '0');
        \$v4808%now\ <= (others => '0');
        \$18811%now\ <= (others => '0');
        \$19808_forever6704342_arg%now\ <= (others => '0');
        \$v4508%now\ <= (others => '0');
        \$v5207%now\ <= (others => '0');
        \$v5093%now\ <= (others => '0');
        \$19034_binop_int6434368_result%now\ <= (others => '0');
        \$19627%now\ <= (others => '0');
        \$19881_hd%now\ <= (others => '0');
        \$19291_v%now\ <= (others => '0');
        \$18901_binop_int6434361_id%now\ <= (others => '0');
        \$19387_compbranch6504394_result%now\ <= (others => '0');
        \$19644_hd%now\ <= (others => '0');
        \$19347_fill6534389_id%now\ <= (others => '0');
        \$v5917%now\ <= (others => '0');
        \$19792%now\ <= (others => '0');
        \$19541%now\ <= (others => '0');
        \$v5480%now\ <= (others => '0');
        \$19415_sp%now\ <= (others => '0');
        \$19262_forever6704385_arg%now\ <= (others => '0');
        \$18477%now\ <= (others => '0');
        \$19635%now\ <= (others => '0');
        \$v4933%now\ <= (others => '0');
        \$19633%now\ <= (others => '0');
        \$v4566%now\ <= (others => '0');
        \$18917_modulo6684349_id%now\ <= (others => '0');
        \$18451%now\ <= (others => '0');
        \$19802%now\ <= (others => '0');
        \$19221%now\ <= (others => '0');
        \$19224%now\ <= (others => '0');
        \$v5240%now\ <= (others => '0');
        \$19516%now\ <= (others => '0');
        \$18656%now\ <= (others => '0');
        \$19693%now\ <= (others => '0');
        \$18496%now\ <= (others => '0');
        \$18588%now\ <= (others => '0');
        \$18887_v%now\ <= (others => '0');
        \$19360_sp%now\ <= (others => '0');
        \$19171_compare6444358_result%now\ <= (others => '0');
        \$19688_hd%now\ <= (others => '0');
        \$18491%now\ <= (others => '0');
        \$18541%now\ <= (others => '0');
        \$19380_compbranch6504393_arg%now\ <= (others => '0');
        \$19782%now\ <= (others => '0');
        \$v5517%now\ <= (others => '0');
        \$19141_modulo6684356_id%now\ <= (others => '0');
        \$19107_modulo6684349_id%now\ <= (others => '0');
        \$v4971%now\ <= (others => '0');
        \$v4848%now\ <= (others => '0');
        \$19166_binop_compare6454377_result%now\ <= (others => '0');
        \$19593%now\ <= (others => '0');
        \$18568%now\ <= (others => '0');
        \$v4625%now\ <= (others => '0');
        \$18452%now\ <= (others => '0');
        \$19742%now\ <= (others => '0');
        \$v4869%now\ <= (others => '0');
        \$v5590%now\ <= (others => '0');
        \$18468_wait662_result%now\ <= (others => '0');
        \$19575_hd%now\ <= (others => '0');
        \$19229_v%now\ <= (others => '0');
        \$18981_res%now\ <= (others => '0');
        \$v4622%now\ <= (others => '0');
        \$18942_v%now\ <= (others => '0');
        \$18543%now\ <= (others => '0');
        \$19513%now\ <= (others => '0');
        \$19555%now\ <= (others => '0');
        \$19692%now\ <= (others => '0');
        \$19370_compare6444359_result%now\ <= (others => '0');
        \$v4896%now\ <= (others => '0');
        \$v5661%now\ <= (others => '0');
        \$v5520%now\ <= (others => '0');
        \$18917_modulo6684349_result%now\ <= (others => '0');
        \$19116_binop_int6434373_result%now\ <= (others => '0');
        \$v4404%now\ <= (others => '0');
        \$19862%now\ <= (others => '0');
        \$18449%now\ <= (others => '0');
        \$19573%now\ <= (others => '0');
        \$19729%now\ <= (others => '0');
        \$18952_modulo6684357_id%now\ <= (others => '0');
        \$19252_forever6704384_arg%now\ <= (others => '0');
        \$19805%now\ <= (others => '0');
        \$18943_res%now\ <= (others => '0');
        \$v4564%now\ <= (others => '0');
        \$18926_modulo6684356_arg%now\ <= (others => '0');
        \$v5438%now\ <= (others => '0');
        \$19567%now\ <= (others => '0');
        \$18761%now\ <= (others => '0');
        \$v5350%now\ <= (others => '0');
        \$v5230%now\ <= (others => '0');
        \$v4731%now\ <= (others => '0');
        \$19838_copy_root_in_ram6634340_arg%now\ <= (others => '0');
        \$v5667%now\ <= (others => '0');
        \$v5535%now\ <= (others => '0');
        \$19008_r%now\ <= (others => '0');
        \$v5547%now\ <= (others => '0');
        \$19669%now\ <= (others => '0');
        \$18862%now\ <= (others => '0');
        \$19699%now\ <= (others => '0');
        \$19630%now\ <= (others => '0');
        \$ram_lock%now\ <= (others => '0');
        \$global_end_lock%now\ <= (others => '0');
        \$code_lock%now\ <= (others => '0');
        \state%now\ <= idle4401;
        \state_var5924%now\ <= idle4436;
        \state_var5923%now\ <= idle4609;
        \state_var5922%now\ <= idle4574;
        \state_var5921%now\ <= idle4965;
        \state_var5920%now\ <= idle4930;
      elsif (rising_edge(clk)) then
        \$18606%now\ <= \$18606%next\;
        \$19190_binop_compare6454380_arg%now\ <= \$19190_binop_compare6454380_arg%next\;
        \$v4743%now\ <= \$v4743%next\;
        \$19072_binop_int6434370_arg%now\ <= \$19072_binop_int6434370_arg%next\;
        \$18910_modulo6684349_id%now\ <= \$18910_modulo6684349_id%next\;
        \$19299%now\ <= \$19299%next\;
        \$19069_modulo6684349_id%now\ <= \$19069_modulo6684349_id%next\;
        \$v5526%now\ <= \$v5526%next\;
        \$v4663%now\ <= \$v4663%next\;
        \$v5913%now\ <= \$v5913%next\;
        \$18602%now\ <= \$18602%next\;
        \$v5541%now\ <= \$v5541%next\;
        \$18809%now\ <= \$18809%next\;
        \$18751%now\ <= \$18751%next\;
        \$19272%now\ <= \$19272%next\;
        \$v5486%now\ <= \$v5486%next\;
        \$v5513%now\ <= \$v5513%next\;
        \$18729%now\ <= \$18729%next\;
        \$v5507%now\ <= \$v5507%next\;
        \$18801%now\ <= \$18801%next\;
        \$19779_loop666_id%now\ <= \$19779_loop666_id%next\;
        \$18775%now\ <= \$18775%next\;
        \$19874%now\ <= \$19874%next\;
        \$v5715%now\ <= \$v5715%next\;
        \$18974_modulo6684349_id%now\ <= \$18974_modulo6684349_id%next\;
        \$19828%now\ <= \$19828%next\;
        \$v4961%now\ <= \$v4961%next\;
        \$v4499%now\ <= \$v4499%next\;
        \$19326_compbranch6504387_result%now\ <= \$19326_compbranch6504387_result%next\;
        \$v5326%now\ <= \$v5326%next\;
        \$v5484%now\ <= \$v5484%next\;
        \$18504%now\ <= \$18504%next\;
        \$v5643%now\ <= \$v5643%next\;
        \$18945_modulo6684356_result%now\ <= \$18945_modulo6684356_result%next\;
        \$18933_modulo6684357_id%now\ <= \$18933_modulo6684357_id%next\;
        \$19250%now\ <= \$19250%next\;
        \$18624%now\ <= \$18624%next\;
        \$v4650%now\ <= \$v4650%next\;
        \$19553%now\ <= \$19553%next\;
        \$18637_w%now\ <= \$18637_w%next\;
        \$19380_compbranch6504393_id%now\ <= \$19380_compbranch6504393_id%next\;
        \$v5619%now\ <= \$v5619%next\;
        \$18835%now\ <= \$18835%next\;
        \$19579%now\ <= \$19579%next\;
        \$19758%now\ <= \$19758%next\;
        \$19085_modulo6684357_result%now\ <= \$19085_modulo6684357_result%next\;
        \$18776%now\ <= \$18776%next\;
        \$18875_v%now\ <= \$18875_v%next\;
        \$19132_modulo6684349_id%now\ <= \$19132_modulo6684349_id%next\;
        \$18619%now\ <= \$18619%next\;
        \$19163_forever6704376_arg%now\ <= \$19163_forever6704376_arg%next\;
        \$v4604%now\ <= \$v4604%next\;
        \$v5699%now\ <= \$v5699%next\;
        \$19292%now\ <= \$19292%next\;
        \$v5634%now\ <= \$v5634%next\;
        \$19416_w36574398_result%now\ <= \$19416_w36574398_result%next\;
        \$18993_modulo6684349_result%now\ <= \$18993_modulo6684349_result%next\;
        \$18581%now\ <= \$18581%next\;
        \$19866_hd%now\ <= \$19866_hd%next\;
        \$v5287%now\ <= \$v5287%next\;
        \$v4467%now\ <= \$v4467%next\;
        \$18900%now\ <= \$18900%next\;
        \$v4470%now\ <= \$v4470%next\;
        \$v4325%now\ <= \$v4325%next\;
        \$18696%now\ <= \$18696%next\;
        \$19245%now\ <= \$19245%next\;
        \$19024_modulo6684349_result%now\ <= \$19024_modulo6684349_result%next\;
        \$18945_modulo6684356_arg%now\ <= \$18945_modulo6684356_arg%next\;
        \$19689%now\ <= \$19689%next\;
        \$v4577%now\ <= \$v4577%next\;
        \$19140_r%now\ <= \$19140_r%next\;
        \$18802%now\ <= \$18802%next\;
        \$v5076%now\ <= \$v5076%next\;
        \$19001_r%now\ <= \$19001_r%next\;
        \$v5532%now\ <= \$v5532%next\;
        \$19501%now\ <= \$19501%next\;
        \$18769_hd%now\ <= \$18769_hd%next\;
        \$v5152%now\ <= \$v5152%next\;
        \$v4703%now\ <= \$v4703%next\;
        \$19122_modulo6684356_result%now\ <= \$19122_modulo6684356_result%next\;
        \$19499_aux664_id%now\ <= \$19499_aux664_id%next\;
        \$18483%now\ <= \$18483%next\;
        \$19290%now\ <= \$19290%next\;
        \$19273%now\ <= \$19273%next\;
        \$19104_modulo6684357_id%now\ <= \$19104_modulo6684357_id%next\;
        \$v4710%now\ <= \$v4710%next\;
        \$v4814%now\ <= \$v4814%next\;
        \$19170_res%now\ <= \$19170_res%next\;
        \$18924_res%now\ <= \$18924_res%next\;
        \$19863%now\ <= \$19863%next\;
        \$18821_v%now\ <= \$18821_v%next\;
        \$19827%now\ <= \$19827%next\;
        \$19432%now\ <= \$19432%next\;
        \$19448_v%now\ <= \$19448_v%next\;
        \$18630%now\ <= \$18630%next\;
        \$19094_v%now\ <= \$19094_v%next\;
        \$v4535%now\ <= \$v4535%next\;
        \$v5551%now\ <= \$v5551%next\;
        \$19028_modulo6684357_result%now\ <= \$19028_modulo6684357_result%next\;
        \$18939_binop_int6434363_result%now\ <= \$18939_binop_int6434363_result%next\;
        \$v5824%now\ <= \$v5824%next\;
        \$18788%now\ <= \$18788%next\;
        \$v5226%now\ <= \$v5226%next\;
        \$18582%now\ <= \$18582%next\;
        \$19081_modulo6684349_arg%now\ <= \$19081_modulo6684349_arg%next\;
        \$v5013%now\ <= \$v5013%next\;
        \$18881_hd%now\ <= \$18881_hd%next\;
        \$19525%now\ <= \$19525%next\;
        \$18509%now\ <= \$18509%next\;
        \$18793_make_block579_result%now\ <= \$18793_make_block579_result%next\;
        \$18974_modulo6684349_arg%now\ <= \$18974_modulo6684349_arg%next\;
        \$19235_v%now\ <= \$19235_v%next\;
        \$v4515%now\ <= \$v4515%next\;
        \$v5323%now\ <= \$v5323%next\;
        \$18655%now\ <= \$18655%next\;
        \$19906%now\ <= \$19906%next\;
        \$v5592%now\ <= \$v5592%next\;
        \$19194_res%now\ <= \$19194_res%next\;
        \$18990_modulo6684357_result%now\ <= \$18990_modulo6684357_result%next\;
        \$19947%now\ <= \$19947%next\;
        \$19672%now\ <= \$19672%next\;
        \$v5692%now\ <= \$v5692%next\;
        \$18474%now\ <= \$18474%next\;
        \$19641%now\ <= \$19641%next\;
        \$18855_next_env%now\ <= \$18855_next_env%next\;
        \$v5158%now\ <= \$v5158%next\;
        \$19040_modulo6684356_id%now\ <= \$19040_modulo6684356_id%next\;
        \$v5369%now\ <= \$v5369%next\;
        \$v5733%now\ <= \$v5733%next\;
        \$19661%now\ <= \$19661%next\;
        \$v5414%now\ <= \$v5414%next\;
        \$v4443%now\ <= \$v4443%next\;
        \$18876%now\ <= \$18876%next\;
        \$19653%now\ <= \$19653%next\;
        \$19508%now\ <= \$19508%next\;
        \$19358%now\ <= \$19358%next\;
        \$v5151%now\ <= \$v5151%next\;
        \$v5594%now\ <= \$v5594%next\;
        \$19043_modulo6684349_result%now\ <= \$19043_modulo6684349_result%next\;
        \$18859%now\ <= \$18859%next\;
        \$v4830%now\ <= \$v4830%next\;
        \$v5117%now\ <= \$v5117%next\;
        \$19445%now\ <= \$19445%next\;
        \$18867%now\ <= \$18867%next\;
        \$v5752%now\ <= \$v5752%next\;
        \$18865%now\ <= \$18865%next\;
        \$19890%now\ <= \$19890%next\;
        \$v4511%now\ <= \$v4511%next\;
        \$18455%now\ <= \$18455%next\;
        \$18512%now\ <= \$18512%next\;
        \$v4590%now\ <= \$v4590%next\;
        \$19427%now\ <= \$19427%next\;
        \$19934_hd%now\ <= \$19934_hd%next\;
        \$18846%now\ <= \$18846%next\;
        \$18524_loop666_result%now\ <= \$18524_loop666_result%next\;
        \$v4472%now\ <= \$v4472%next\;
        \$19723%now\ <= \$19723%next\;
        \$18778%now\ <= \$18778%next\;
        \$18694%now\ <= \$18694%next\;
        \$v5759%now\ <= \$v5759%next\;
        \$19066_modulo6684357_result%now\ <= \$19066_modulo6684357_result%next\;
        \$19850_w%now\ <= \$19850_w%next\;
        \$19419%now\ <= \$19419%next\;
        \$18961_v%now\ <= \$18961_v%next\;
        \$19201_v%now\ <= \$19201_v%next\;
        \$v5703%now\ <= \$v5703%next\;
        \$19274_v%now\ <= \$19274_v%next\;
        \$19394_compbranch6504395_arg%now\ <= \$19394_compbranch6504395_arg%next\;
        \$v5320%now\ <= \$v5320%next\;
        \$19166_binop_compare6454377_arg%now\ <= \$19166_binop_compare6454377_arg%next\;
        \$v5212%now\ <= \$v5212%next\;
        \$19704%now\ <= \$19704%next\;
        \$19930%now\ <= \$19930%next\;
        \$v5721%now\ <= \$v5721%next\;
        \$19458%now\ <= \$19458%next\;
        \$19185_v%now\ <= \$19185_v%next\;
        \$v5586%now\ <= \$v5586%next\;
        \$18738_next%now\ <= \$18738_next%next\;
        \$19364_v%now\ <= \$19364_v%next\;
        \$v5234%now\ <= \$v5234%next\;
        \$v5760%now\ <= \$v5760%next\;
        \$18974_modulo6684349_result%now\ <= \$18974_modulo6684349_result%next\;
        \$19797_next%now\ <= \$19797_next%next\;
        \$18745_hd%now\ <= \$18745_hd%next\;
        \$18797_branch_if648_result%now\ <= \$18797_branch_if648_result%next\;
        \$19589_copy_root_in_ram6634353_id%now\ <= \$19589_copy_root_in_ram6634353_id%next\;
        \$v5766%now\ <= \$v5766%next\;
        \$19478_v%now\ <= \$19478_v%next\;
        \$19752%now\ <= \$19752%next\;
        \$v4616%now\ <= \$v4616%next\;
        \$19894%now\ <= \$19894%next\;
        \$19819%now\ <= \$19819%next\;
        \$19489%now\ <= \$19489%next\;
        \$v5776%now\ <= \$v5776%next\;
        \$v5019%now\ <= \$v5019%next\;
        \$18807%now\ <= \$18807%next\;
        \$19504%now\ <= \$19504%next\;
        \$18650%now\ <= \$18650%next\;
        \$18837%now\ <= \$18837%next\;
        \$18569%now\ <= \$18569%next\;
        \$19129_modulo6684357_id%now\ <= \$19129_modulo6684357_id%next\;
        \$18805%now\ <= \$18805%next\;
        \$v5869%now\ <= \$v5869%next\;
        \$19112%now\ <= \$19112%next\;
        \$19135_binop_int6434374_arg%now\ <= \$19135_binop_int6434374_arg%next\;
        \$19002_modulo6684356_arg%now\ <= \$19002_modulo6684356_arg%next\;
        \$v5515%now\ <= \$v5515%next\;
        \$19319%now\ <= \$19319%next\;
        \$v5646%now\ <= \$v5646%next\;
        \$v4952%now\ <= \$v4952%next\;
        \$v5610%now\ <= \$v5610%next\;
        \$v5683%now\ <= \$v5683%next\;
        \$18958_binop_int6434364_result%now\ <= \$18958_binop_int6434364_result%next\;
        \$19342%now\ <= \$19342%next\;
        \$19657%now\ <= \$19657%next\;
        \$19777%now\ <= \$19777%next\;
        \$19620%now\ <= \$19620%next\;
        \$18793_make_block579_id%now\ <= \$18793_make_block579_id%next\;
        \$18521_loop666_arg%now\ <= \$18521_loop666_arg%next\;
        \$19803%now\ <= \$19803%next\;
        \$19217%now\ <= \$19217%next\;
        \$v4949%now\ <= \$v4949%next\;
        \$19486%now\ <= \$19486%next\;
        \$v5857%now\ <= \$v5857%next\;
        \$18482%now\ <= \$18482%next\;
        \$v4692%now\ <= \$v4692%next\;
        \$19309_v%now\ <= \$19309_v%next\;
        \$18529%now\ <= \$18529%next\;
        \$19916%now\ <= \$19916%next\;
        \$v5686%now\ <= \$v5686%next\;
        \$v4854%now\ <= \$v4854%next\;
        \$v4628%now\ <= \$v4628%next\;
        \$18703%now\ <= \$18703%next\;
        \$v5506%now\ <= \$v5506%next\;
        \$v4926%now\ <= \$v4926%next\;
        \$19829%now\ <= \$19829%next\;
        \$v4523%now\ <= \$v4523%next\;
        \$v4569%now\ <= \$v4569%next\;
        \$v5749%now\ <= \$v5749%next\;
        \$19209_v%now\ <= \$19209_v%next\;
        \$19482%now\ <= \$19482%next\;
        \$19611%now\ <= \$19611%next\;
        \$19811_copy_root_in_ram6634341_id%now\ <= \$19811_copy_root_in_ram6634341_id%next\;
        \$19784%now\ <= \$19784%next\;
        \$18502%now\ <= \$18502%next\;
        \$v4770%now\ <= \$v4770%next\;
        \$18667_w%now\ <= \$18667_w%next\;
        \$19434%now\ <= \$19434%next\;
        \$19333_compbranch6504388_arg%now\ <= \$19333_compbranch6504388_arg%next\;
        \$19732%now\ <= \$19732%next\;
        \$19609%now\ <= \$19609%next\;
        \$19714_next%now\ <= \$19714_next%next\;
        \$18815%now\ <= \$18815%next\;
        \$v5210%now\ <= \$v5210%next\;
        \$18565%now\ <= \$18565%next\;
        \$v4491%now\ <= \$v4491%next\;
        \$19076_res%now\ <= \$19076_res%next\;
        \$v4727%now\ <= \$v4727%next\;
        \$19015_binop_int6434367_id%now\ <= \$19015_binop_int6434367_id%next\;
        \$18986_modulo6684349_arg%now\ <= \$18986_modulo6684349_arg%next\;
        \$v4734%now\ <= \$v4734%next\;
        \$19656%now\ <= \$19656%next\;
        \$19496_aux664_arg%now\ <= \$19496_aux664_arg%next\;
        \$18480%now\ <= \$18480%next\;
        \$v5537%now\ <= \$v5537%next\;
        \$18458%now\ <= \$18458%next\;
        \$18993_modulo6684349_arg%now\ <= \$18993_modulo6684349_arg%next\;
        \$v5655%now\ <= \$v5655%next\;
        \$19294%now\ <= \$19294%next\;
        \$v5828%now\ <= \$v5828%next\;
        \$19583%now\ <= \$19583%next\;
        \$v5838%now\ <= \$v5838%next\;
        \$19163_forever6704376_id%now\ <= \$19163_forever6704376_id%next\;
        \$18723%now\ <= \$18723%next\;
        \$v4481%now\ <= \$v4481%next\;
        \$v5640%now\ <= \$v5640%next\;
        \$19314%now\ <= \$19314%next\;
        \$18762%now\ <= \$18762%next\;
        \$19034_binop_int6434368_arg%now\ <= \$19034_binop_int6434368_arg%next\;
        \$v4728%now\ <= \$v4728%next\;
        \$v4596%now\ <= \$v4596%next\;
        \$19062_modulo6684349_result%now\ <= \$19062_modulo6684349_result%next\;
        \$18914_modulo6684357_arg%now\ <= \$18914_modulo6684357_arg%next\;
        \$18590%now\ <= \$18590%next\;
        \$19902%now\ <= \$19902%next\;
        \$18670%now\ <= \$18670%next\;
        \$v5604%now\ <= \$v5604%next\;
        \$19248%now\ <= \$19248%next\;
        \$19088_modulo6684349_result%now\ <= \$19088_modulo6684349_result%next\;
        \$19464%now\ <= \$19464%next\;
        \$19072_binop_int6434370_result%now\ <= \$19072_binop_int6434370_result%next\;
        \$v4761%now\ <= \$v4761%next\;
        \$19816%now\ <= \$19816%next\;
        \$19081_modulo6684349_result%now\ <= \$19081_modulo6684349_result%next\;
        \$v4845%now\ <= \$v4845%next\;
        \$v4631%now\ <= \$v4631%next\;
        \$19326_compbranch6504387_arg%now\ <= \$19326_compbranch6504387_arg%next\;
        \$v5035%now\ <= \$v5035%next\;
        \$18685%now\ <= \$18685%next\;
        \$v5603%now\ <= \$v5603%next\;
        \$19628_w%now\ <= \$19628_w%next\;
        \$v5582%now\ <= \$v5582%next\;
        \$18948_modulo6684349_arg%now\ <= \$18948_modulo6684349_arg%next\;
        \$v5060%now\ <= \$v5060%next\;
        \$18668_hd%now\ <= \$18668_hd%next\;
        \$v4552%now\ <= \$v4552%next\;
        \$19187_compare6444358_result%now\ <= \$19187_compare6444358_result%next\;
        \$v5378%now\ <= \$v5378%next\;
        \$19623%now\ <= \$19623%next\;
        \$v5052%now\ <= \$v5052%next\;
        \$v4946%now\ <= \$v4946%next\;
        \$18664%now\ <= \$18664%next\;
        \$18646%now\ <= \$18646%next\;
        \$18852%now\ <= \$18852%next\;
        \$18485%now\ <= \$18485%next\;
        \$19190_binop_compare6454380_result%now\ <= \$19190_binop_compare6454380_result%next\;
        \$19043_modulo6684349_arg%now\ <= \$19043_modulo6684349_arg%next\;
        \$v4936%now\ <= \$v4936%next\;
        \$v4417%now\ <= \$v4417%next\;
        \$18447%now\ <= \$18447%next\;
        \$v4992%now\ <= \$v4992%next\;
        \$v5702%now\ <= \$v5702%next\;
        \$18967_modulo6684349_arg%now\ <= \$18967_modulo6684349_arg%next\;
        \$v5481%now\ <= \$v5481%next\;
        \$18952_modulo6684357_result%now\ <= \$18952_modulo6684357_result%next\;
        \$18662%now\ <= \$18662%next\;
        \$18600%now\ <= \$18600%next\;
        \$v5244%now\ <= \$v5244%next\;
        \$19600%now\ <= \$19600%next\;
        \$19838_copy_root_in_ram6634340_result%now\ <= \$19838_copy_root_in_ram6634340_result%next\;
        \$19885%now\ <= \$19885%next\;
        \$19685%now\ <= \$19685%next\;
        \$19187_compare6444358_id%now\ <= \$19187_compare6444358_id%next\;
        \$18926_modulo6684356_id%now\ <= \$18926_modulo6684356_id%next\;
        \$19720_w%now\ <= \$19720_w%next\;
        \$v5530%now\ <= \$v5530%next\;
        \$18644%now\ <= \$18644%next\;
        \$18466_loop666_id%now\ <= \$18466_loop666_id%next\;
        \$18638_hd%now\ <= \$18638_hd%next\;
        \$v4674%now\ <= \$v4674%next\;
        \$v5250%now\ <= \$v5250%next\;
        \$18563%now\ <= \$18563%next\;
        \$19062_modulo6684349_id%now\ <= \$19062_modulo6684349_id%next\;
        \$18645%now\ <= \$18645%next\;
        \$19897%now\ <= \$19897%next\;
        \$19139_res%now\ <= \$19139_res%next\;
        \$19347_fill6534389_arg%now\ <= \$19347_fill6534389_arg%next\;
        \$19495_loop665_arg%now\ <= \$19495_loop665_arg%next\;
        \$v4695%now\ <= \$v4695%next\;
        \$18576%now\ <= \$18576%next\;
        \$18578%now\ <= \$18578%next\;
        \$18440_make_block579_arg%now\ <= \$18440_make_block579_arg%next\;
        \$19157_forever6704375_id%now\ <= \$19157_forever6704375_id%next\;
        \$19246_v%now\ <= \$19246_v%next\;
        \$19495_loop665_id%now\ <= \$19495_loop665_id%next\;
        \$19515_next%now\ <= \$19515_next%next\;
        \$v4563%now\ <= \$v4563%next\;
        \$v4908%now\ <= \$v4908%next\;
        \$18635%now\ <= \$18635%next\;
        \$19251%now\ <= \$19251%next\;
        \$19648%now\ <= \$19648%next\;
        \$18613_copy_root_in_ram6634346_id%now\ <= \$18613_copy_root_in_ram6634346_id%next\;
        \$19780_loop665_arg%now\ <= \$19780_loop665_arg%next\;
        \$18571_copy_root_in_ram6634345_arg%now\ <= \$18571_copy_root_in_ram6634345_arg%next\;
        \$v5120%now\ <= \$v5120%next\;
        \$19854%now\ <= \$19854%next\;
        \$v4988%now\ <= \$v4988%next\;
        \$v5607%now\ <= \$v5607%next\;
        \$19848%now\ <= \$19848%next\;
        \$19232%now\ <= \$19232%next\;
        \$19814%now\ <= \$19814%next\;
        \$v4680%now\ <= \$v4680%next\;
        \$18906_r%now\ <= \$18906_r%next\;
        \$v5127%now\ <= \$v5127%next\;
        \$18620%now\ <= \$18620%next\;
        \$19887%now\ <= \$19887%next\;
        \$19296_v%now\ <= \$19296_v%next\;
        \$18709%now\ <= \$18709%next\;
        \$v4805%now\ <= \$v4805%next\;
        \$v5514%now\ <= \$v5514%next\;
        \$18913_r%now\ <= \$18913_r%next\;
        \$18457%now\ <= \$18457%next\;
        \$19269%now\ <= \$19269%next\;
        \$19569%now\ <= \$19569%next\;
        \$v5823%now\ <= \$v5823%next\;
        \$v5164%now\ <= \$v5164%next\;
        \$19721_hd%now\ <= \$19721_hd%next\;
        \$v5831%now\ <= \$v5831%next\;
        \$v4740%now\ <= \$v4740%next\;
        \$v5308%now\ <= \$v5308%next\;
        \$v4995%now\ <= \$v4995%next\;
        \$v4601%now\ <= \$v4601%next\;
        \$18484%now\ <= \$18484%next\;
        \$18733%now\ <= \$18733%next\;
        \$v4660%now\ <= \$v4660%next\;
        \$19408_argument3%now\ <= \$19408_argument3%next\;
        \$18828_v%now\ <= \$18828_v%next\;
        \$19390_b%now\ <= \$19390_b%next\;
        \$19727%now\ <= \$19727%next\;
        \$18510%now\ <= \$18510%next\;
        \$19662%now\ <= \$19662%next\;
        \$v5577%now\ <= \$v5577%next\;
        \$19015_binop_int6434367_arg%now\ <= \$19015_binop_int6434367_arg%next\;
        \$19413%now\ <= \$19413%next\;
        \$v4584%now\ <= \$v4584%next\;
        \$19845%now\ <= \$19845%next\;
        \$19337_compare6444359_id%now\ <= \$19337_compare6444359_id%next\;
        \$19698%now\ <= \$19698%next\;
        \$18566%now\ <= \$18566%next\;
        \$18767%now\ <= \$18767%next\;
        \$19359%now\ <= \$19359%next\;
        \$18977_binop_int6434365_arg%now\ <= \$18977_binop_int6434365_arg%next\;
        \$v4878%now\ <= \$v4878%next\;
        \$19267_hd%now\ <= \$19267_hd%next\;
        \$19679%now\ <= \$19679%next\;
        \$v5195%now\ <= \$v5195%next\;
        \$v4433%now\ <= \$v4433%next\;
        \$18864%now\ <= \$18864%next\;
        \$18996_binop_int6434366_arg%now\ <= \$18996_binop_int6434366_arg%next\;
        \$19599%now\ <= \$19599%next\;
        \$19526_forever6704355_arg%now\ <= \$19526_forever6704355_arg%next\;
        \$19578%now\ <= \$19578%next\;
        \$18605%now\ <= \$18605%next\;
        \$19558%now\ <= \$19558%next\;
        \$19280%now\ <= \$19280%next\;
        \$v5278%now\ <= \$v5278%next\;
        \$v5557%now\ <= \$v5557%next\;
        \$19817%now\ <= \$19817%next\;
        \$19238_w6514383_arg%now\ <= \$19238_w6514383_arg%next\;
        \$v5284%now\ <= \$v5284%next\;
        \$v5905%now\ <= \$v5905%next\;
        \$19488%now\ <= \$19488%next\;
        \$19474%now\ <= \$19474%next\;
        \$v5564%now\ <= \$v5564%next\;
        \$18591%now\ <= \$18591%next\;
        \$v4568%now\ <= \$v4568%next\;
        \$v5883%now\ <= \$v5883%next\;
        \$v5555%now\ <= \$v5555%next\;
        \$19726%now\ <= \$19726%next\;
        \$v4842%now\ <= \$v4842%next\;
        \$18834_v%now\ <= \$18834_v%next\;
        \$19401_compbranch6504396_result%now\ <= \$19401_compbranch6504396_result%next\;
        \$18699%now\ <= \$18699%next\;
        \$18680%now\ <= \$18680%next\;
        \$19751%now\ <= \$19751%next\;
        \$19157_forever6704375_arg%now\ <= \$19157_forever6704375_arg%next\;
        \$18584_hd%now\ <= \$18584_hd%next\;
        \$19867%now\ <= \$19867%next\;
        \$v5465%now\ <= \$v5465%next\;
        \$18999_v%now\ <= \$18999_v%next\;
        \$18623%now\ <= \$18623%next\;
        \$19754%now\ <= \$19754%next\;
        \$19825%now\ <= \$19825%next\;
        \$19312_v%now\ <= \$19312_v%next\;
        \$18936_modulo6684349_arg%now\ <= \$18936_modulo6684349_arg%next\;
        \$18460%now\ <= \$18460%next\;
        \$19596%now\ <= \$19596%next\;
        \$18795_offsetclosure_n639_result%now\ <= \$18795_offsetclosure_n639_result%next\;
        \$19918%now\ <= \$19918%next\;
        \$v4328%now\ <= \$v4328%next\;
        \$19373_compbranch6504392_result%now\ <= \$19373_compbranch6504392_result%next\;
        \$v5247%now\ <= \$v5247%next\;
        \$v4543%now\ <= \$v4543%next\;
        \$v5420%now\ <= \$v5420%next\;
        \$19505%now\ <= \$19505%next\;
        \$18570%now\ <= \$18570%next\;
        \$v5263%now\ <= \$v5263%next\;
        \$19391_compare6444359_id%now\ <= \$19391_compare6444359_id%next\;
        \$v5835%now\ <= \$v5835%next\;
        \$18962_res%now\ <= \$18962_res%next\;
        \$18822_v%now\ <= \$18822_v%next\;
        \$v5614%now\ <= \$v5614%next\;
        \$v5027%now\ <= \$v5027%next\;
        \$18610%now\ <= \$18610%next\;
        \$v5069%now\ <= \$v5069%next\;
        \$18684%now\ <= \$18684%next\;
        \$19535_copy_root_in_ram6634354_id%now\ <= \$19535_copy_root_in_ram6634354_id%next\;
        \$v5860%now\ <= \$v5860%next\;
        \$v4414%now\ <= \$v4414%next\;
        \$v5237%now\ <= \$v5237%next\;
        \$19066_modulo6684357_arg%now\ <= \$19066_modulo6684357_arg%next\;
        \$19852%now\ <= \$19852%next\;
        \$18577%now\ <= \$18577%next\;
        \$v5533%now\ <= \$v5533%next\;
        \$18553_forever6704348_arg%now\ <= \$18553_forever6704348_arg%next\;
        \$19387_compbranch6504394_id%now\ <= \$19387_compbranch6504394_id%next\;
        \$18643%now\ <= \$18643%next\;
        \$18754%now\ <= \$18754%next\;
        \$18933_modulo6684357_arg%now\ <= \$18933_modulo6684357_arg%next\;
        \$19397_b%now\ <= \$19397_b%next\;
        \$19279_v%now\ <= \$19279_v%next\;
        \$18933_modulo6684357_result%now\ <= \$18933_modulo6684357_result%next\;
        \$v5485%now\ <= \$v5485%next\;
        \$19550%now\ <= \$19550%next\;
        \$18816%now\ <= \$18816%next\;
        \$19495_loop665_result%now\ <= \$19495_loop665_result%next\;
        \$v5516%now\ <= \$v5516%next\;
        \$v5180%now\ <= \$v5180%next\;
        \$18952_modulo6684357_arg%now\ <= \$18952_modulo6684357_arg%next\;
        \$19855%now\ <= \$19855%next\;
        \$v5426%now\ <= \$v5426%next\;
        \$19313%now\ <= \$19313%next\;
        \$v5542%now\ <= \$v5542%next\;
        \$19565%now\ <= \$19565%next\;
        \$v4863%now\ <= \$v4863%next\;
        \$18980_v%now\ <= \$18980_v%next\;
        \$18521_loop666_id%now\ <= \$18521_loop666_id%next\;
        \$v5870%now\ <= \$v5870%next\;
        \$19800_next%now\ <= \$19800_next%next\;
        \$19746%now\ <= \$19746%next\;
        \$19851_hd%now\ <= \$19851_hd%next\;
        \$18488%now\ <= \$18488%next\;
        \$18746%now\ <= \$18746%next\;
        \$v5203%now\ <= \$v5203%next\;
        \$19222%now\ <= \$19222%next\;
        \$v5290%now\ <= \$v5290%next\;
        \$18796_make_block_n646_id%now\ <= \$18796_make_block_n646_id%next\;
        \$19096_r%now\ <= \$19096_r%next\;
        \$19450_v%now\ <= \$19450_v%next\;
        \$19651%now\ <= \$19651%next\;
        \$v5130%now\ <= \$v5130%next\;
        \$v5595%now\ <= \$v5595%next\;
        \$v4699%now\ <= \$v4699%next\;
        \$18559_copy_root_in_ram6634347_result%now\ <= \$18559_copy_root_in_ram6634347_result%next\;
        \$18831%now\ <= \$18831%next\;
        \$v5123%now\ <= \$v5123%next\;
        \$18829%now\ <= \$18829%next\;
        \$19761%now\ <= \$19761%next\;
        \$19547_copy_root_in_ram6634352_result%now\ <= \$19547_copy_root_in_ram6634352_result%next\;
        \$v5737%now\ <= \$v5737%next\;
        \$19676%now\ <= \$19676%next\;
        \$18450%now\ <= \$18450%next\;
        \$18982_r%now\ <= \$18982_r%next\;
        \$19179_compare6444358_arg%now\ <= \$19179_compare6444358_arg%next\;
        \$v4462%now\ <= \$v4462%next\;
        \$18717%now\ <= \$18717%next\;
        \$v5148%now\ <= \$v5148%next\;
        \$18571_copy_root_in_ram6634345_id%now\ <= \$18571_copy_root_in_ram6634345_id%next\;
        \$v5170%now\ <= \$v5170%next\;
        \$19438%now\ <= \$19438%next\;
        \$19647%now\ <= \$19647%next\;
        \$19483%now\ <= \$19483%next\;
        \$19361_fill6544390_arg%now\ <= \$19361_fill6544390_arg%next\;
        \$19861%now\ <= \$19861%next\;
        \$19211_compare6444358_id%now\ <= \$19211_compare6444358_id%next\;
        \$19786%now\ <= \$19786%next\;
        \$18725%now\ <= \$18725%next\;
        \$18459%now\ <= \$18459%next\;
        \$19135_binop_int6434374_result%now\ <= \$19135_binop_int6434374_result%next\;
        \$v5546%now\ <= \$v5546%next\;
        \$19724%now\ <= \$19724%next\;
        \$18711_w%now\ <= \$18711_w%next\;
        \$18948_modulo6684349_result%now\ <= \$18948_modulo6684349_result%next\;
        \$v5144%now\ <= \$v5144%next\;
        \$19908%now\ <= \$19908%next\;
        \$19858%now\ <= \$19858%next\;
        \$18779%now\ <= \$18779%next\;
        \$v5272%now\ <= \$v5272%next\;
        \$18612%now\ <= \$18612%next\;
        \$19303%now\ <= \$19303%next\;
        \$19551%now\ <= \$19551%next\;
        \$v5269%now\ <= \$v5269%next\;
        \$19186_res%now\ <= \$19186_res%next\;
        \$18689%now\ <= \$18689%next\;
        \$19631%now\ <= \$19631%next\;
        \$18791_loop665_arg%now\ <= \$18791_loop665_arg%next\;
        \$18905_res%now\ <= \$18905_res%next\;
        \$19694%now\ <= \$19694%next\;
        \$18755%now\ <= \$18755%next\;
        \$v5795%now\ <= \$v5795%next\;
        \$v5202%now\ <= \$v5202%next\;
        \$v5565%now\ <= \$v5565%next\;
        \$v4923%now\ <= \$v4923%next\;
        \$19835%now\ <= \$19835%next\;
        \$19588%now\ <= \$19588%next\;
        \$v4943%now\ <= \$v4943%next\;
        \$19078_modulo6684356_id%now\ <= \$19078_modulo6684356_id%next\;
        \$v5317%now\ <= \$v5317%next\;
        \result4434%now\ <= \result4434%next\;
        \$v5512%now\ <= \$v5512%next\;
        \$18465%now\ <= \$18465%next\;
        \$v4484%now\ <= \$v4484%next\;
        \$18830_v%now\ <= \$18830_v%next\;
        \$19779_loop666_arg%now\ <= \$19779_loop666_arg%next\;
        \$19616%now\ <= \$19616%next\;
        \$v4792%now\ <= \$v4792%next\;
        \$19088_modulo6684349_arg%now\ <= \$19088_modulo6684349_arg%next\;
        \$19666%now\ <= \$19666%next\;
        \$19179_compare6444358_id%now\ <= \$19179_compare6444358_id%next\;
        \$19681_next%now\ <= \$19681_next%next\;
        \$18742%now\ <= \$18742%next\;
        \$18795_offsetclosure_n639_arg%now\ <= \$18795_offsetclosure_n639_arg%next\;
        \$19384_compare6444359_id%now\ <= \$19384_compare6444359_id%next\;
        \$18993_modulo6684349_id%now\ <= \$18993_modulo6684349_id%next\;
        \$19610%now\ <= \$19610%next\;
        \$18856_loop_push6494360_arg%now\ <= \$18856_loop_push6494360_arg%next\;
        \$19909_w%now\ <= \$19909_w%next\;
        \$19686%now\ <= \$19686%next\;
        \$v4975%now\ <= \$v4975%next\;
        \$19019_res%now\ <= \$19019_res%next\;
        \$v5534%now\ <= \$v5534%next\;
        \$18479%now\ <= \$18479%next\;
        \$18525_loop665_result%now\ <= \$18525_loop665_result%next\;
        \$v5893%now\ <= \$v5893%next\;
        \$19671%now\ <= \$19671%next\;
        \$v4475%now\ <= \$v4475%next\;
        \$18734%now\ <= \$18734%next\;
        \$19128_r%now\ <= \$19128_r%next\;
        \$19750%now\ <= \$19750%next\;
        \$19499_aux664_arg%now\ <= \$19499_aux664_arg%next\;
        \$19826%now\ <= \$19826%next\;
        \$18799_w1656_result%now\ <= \$18799_w1656_result%next\;
        \$18798_w652_result%now\ <= \$18798_w652_result%next\;
        \$18467_loop665_arg%now\ <= \$18467_loop665_arg%next\;
        \$19021_modulo6684356_id%now\ <= \$19021_modulo6684356_id%next\;
        \$19088_modulo6684349_id%now\ <= \$19088_modulo6684349_id%next\;
        \$19162%now\ <= \$19162%next\;
        \$v4851%now\ <= \$v4851%next\;
        \$19357_v%now\ <= \$19357_v%next\;
        \$19097_modulo6684356_result%now\ <= \$19097_modulo6684356_result%next\;
        \$v5580%now\ <= \$v5580%next\;
        \$19012_modulo6684349_id%now\ <= \$19012_modulo6684349_id%next\;
        \$18765%now\ <= \$18765%next\;
        \$v4893%now\ <= \$v4893%next\;
        \$v5329%now\ <= \$v5329%next\;
        \$19936%now\ <= \$19936%next\;
        \$19020_r%now\ <= \$19020_r%next\;
        \$19238_w6514383_result%now\ <= \$19238_w6514383_result%next\;
        \$v5601%now\ <= \$v5601%next\;
        \$18996_binop_int6434366_id%now\ <= \$18996_binop_int6434366_id%next\;
        \$v5511%now\ <= \$v5511%next\;
        \$v4570%now\ <= \$v4570%next\;
        \$19675%now\ <= \$19675%next\;
        \$18601%now\ <= \$18601%next\;
        \$v4565%now\ <= \$v4565%next\;
        \$18552%now\ <= \$18552%next\;
        \$19077_r%now\ <= \$19077_r%next\;
        \$v5545%now\ <= \$v5545%next\;
        \$v5031%now\ <= \$v5031%next\;
        \$v5456%now\ <= \$v5456%next\;
        \$v5161%now\ <= \$v5161%next\;
        \$19075_v%now\ <= \$19075_v%next\;
        \$18791_loop665_result%now\ <= \$18791_loop665_result%next\;
        \$18750%now\ <= \$18750%next\;
        \$18718%now\ <= \$18718%next\;
        \$19849%now\ <= \$19849%next\;
        \$19059_modulo6684356_arg%now\ <= \$19059_modulo6684356_arg%next\;
        \$v4724%now\ <= \$v4724%next\;
        \$19423_v%now\ <= \$19423_v%next\;
        \$19352%now\ <= \$19352%next\;
        \$19601_copy_root_in_ram6634352_result%now\ <= \$19601_copy_root_in_ram6634352_result%next\;
        \$18789%now\ <= \$18789%next\;
        \$18977_binop_int6434365_id%now\ <= \$18977_binop_int6434365_id%next\;
        \$v5789%now\ <= \$v5789%next\;
        \$v5450%now\ <= \$v5450%next\;
        \$18681%now\ <= \$18681%next\;
        \$19206_binop_compare6454382_arg%now\ <= \$19206_binop_compare6454382_arg%next\;
        \$v5010%now\ <= \$v5010%next\;
        \$19523%now\ <= \$19523%next\;
        \$18964_modulo6684356_id%now\ <= \$18964_modulo6684356_id%next\;
        \$19923%now\ <= \$19923%next\;
        \$19361_fill6544390_result%now\ <= \$19361_fill6544390_result%next\;
        \$19535_copy_root_in_ram6634354_arg%now\ <= \$19535_copy_root_in_ram6634354_arg%next\;
        \$19564%now\ <= \$19564%next\;
        \$18770%now\ <= \$18770%next\;
        \$19790%now\ <= \$19790%next\;
        \$19509%now\ <= \$19509%next\;
        \$18598_w%now\ <= \$18598_w%next\;
        \$18462%now\ <= \$18462%next\;
        \$19873%now\ <= \$19873%next\;
        \$v5496%now\ <= \$v5496%next\;
        \$v5573%now\ <= \$v5573%next\;
        \$19177_v%now\ <= \$19177_v%next\;
        \$19320_forever6704386_arg%now\ <= \$19320_forever6704386_arg%next\;
        \$19069_modulo6684349_arg%now\ <= \$19069_modulo6684349_arg%next\;
        \$v5225%now\ <= \$v5225%next\;
        \$v5611%now\ <= \$v5611%next\;
        \$v5063%now\ <= \$v5063%next\;
        \$v5393%now\ <= \$v5393%next\;
        \$19778%now\ <= \$19778%next\;
        \$19821%now\ <= \$19821%next\;
        \$v5174%now\ <= \$v5174%next\;
        \$18494%now\ <= \$18494%next\;
        \$19333_compbranch6504388_result%now\ <= \$19333_compbranch6504388_result%next\;
        \$19441_arg%now\ <= \$19441_arg%next\;
        \$18920_binop_int6434362_arg%now\ <= \$18920_binop_int6434362_arg%next\;
        \$v5080%now\ <= \$v5080%next\;
        \$18790_loop666_id%now\ <= \$18790_loop666_id%next\;
        \$v5763%now\ <= \$v5763%next\;
        \$v5618%now\ <= \$v5618%next\;
        \$18613_copy_root_in_ram6634346_result%now\ <= \$18613_copy_root_in_ram6634346_result%next\;
        \$19498_loop665_arg%now\ <= \$19498_loop665_arg%next\;
        \$19467_sp%now\ <= \$19467_sp%next\;
        \$v4799%now\ <= \$v4799%next\;
        \$19187_compare6444358_arg%now\ <= \$19187_compare6444358_arg%next\;
        \$v4860%now\ <= \$v4860%next\;
        \$18849%now\ <= \$18849%next\;
        \$18749%now\ <= \$18749%next\;
        \$18907_modulo6684356_id%now\ <= \$18907_modulo6684356_id%next\;
        \$19794%now\ <= \$19794%next\;
        \$18863%now\ <= \$18863%next\;
        \$19910_hd%now\ <= \$19910_hd%next\;
        \$18958_binop_int6434364_id%now\ <= \$18958_binop_int6434364_id%next\;
        \$v5135%now\ <= \$v5135%next\;
        \$v4495%now\ <= \$v4495%next\;
        \$19320_forever6704386_id%now\ <= \$19320_forever6704386_id%next\;
        \$19300%now\ <= \$19300%next\;
        \$19116_binop_int6434373_arg%now\ <= \$19116_binop_int6434373_arg%next\;
        \$v5147%now\ <= \$v5147%next\;
        \$v4899%now\ <= \$v4899%next\;
        \$19333_compbranch6504388_id%now\ <= \$19333_compbranch6504388_id%next\;
        \$19880_w%now\ <= \$19880_w%next\;
        \$v5730%now\ <= \$v5730%next\;
        \$19366_compbranch6504391_arg%now\ <= \$19366_compbranch6504391_arg%next\;
        \$v5007%now\ <= \$v5007%next\;
        \$19377_compare6444359_result%now\ <= \$19377_compare6444359_result%next\;
        \$19203_compare6444358_result%now\ <= \$19203_compare6444358_result%next\;
        \$v5570%now\ <= \$v5570%next\;
        \$19664%now\ <= \$19664%next\;
        \$19637%now\ <= \$19637%next\;
        \$18926_modulo6684356_result%now\ <= \$18926_modulo6684356_result%next\;
        \$v4431%now\ <= \$v4431%next\;
        \$18854_sp%now\ <= \$18854_sp%next\;
        \$19710%now\ <= \$19710%next\;
        \$19771%now\ <= \$19771%next\;
        \$19057_res%now\ <= \$19057_res%next\;
        \$18907_modulo6684356_arg%now\ <= \$18907_modulo6684356_arg%next\;
        \$18537%now\ <= \$18537%next\;
        \$19785%now\ <= \$19785%next\;
        \$18792_wait662_result%now\ <= \$18792_wait662_result%next\;
        \$18826%now\ <= \$18826%next\;
        \$19307_v%now\ <= \$19307_v%next\;
        \$19354_v%now\ <= \$19354_v%next\;
        \$19463%now\ <= \$19463%next\;
        \$19734%now\ <= \$19734%next\;
        \rdy4929%now\ <= \rdy4929%next\;
        \$18799_w1656_id%now\ <= \$18799_w1656_id%next\;
        \$19589_copy_root_in_ram6634353_result%now\ <= \$19589_copy_root_in_ram6634353_result%next\;
        \$18472%now\ <= \$18472%next\;
        \$v4666%now\ <= \$v4666%next\;
        \$19129_modulo6684357_arg%now\ <= \$19129_modulo6684357_arg%next\;
        \$v4458%now\ <= \$v4458%next\;
        \$18873_v%now\ <= \$18873_v%next\;
        \$19038_res%now\ <= \$19038_res%next\;
        \$19595%now\ <= \$19595%next\;
        \$19883%now\ <= \$19883%next\;
        \$18677%now\ <= \$18677%next\;
        \$19249%now\ <= \$19249%next\;
        \$v5266%now\ <= \$v5266%next\;
        \$19546%now\ <= \$19546%next\;
        \$v4767%now\ <= \$v4767%next\;
        \$v5189%now\ <= \$v5189%next\;
        \$v4442%now\ <= \$v4442%next\;
        \$19891%now\ <= \$19891%next\;
        \$v5649%now\ <= \$v5649%next\;
        \$v5199%now\ <= \$v5199%next\;
        \$19559_w%now\ <= \$19559_w%next\;
        \$19920%now\ <= \$19920%next\;
        \$v4549%now\ <= \$v4549%next\;
        \$18990_modulo6684357_id%now\ <= \$18990_modulo6684357_id%next\;
        \$19107_modulo6684349_arg%now\ <= \$19107_modulo6684349_arg%next\;
        \$18520%now\ <= \$18520%next\;
        \$19420_w06554397_result%now\ <= \$19420_w06554397_result%next\;
        \$18884_v%now\ <= \$18884_v%next\;
        \$18925_r%now\ <= \$18925_r%next\;
        \$19179_compare6444358_result%now\ <= \$19179_compare6444358_result%next\;
        \$19078_modulo6684356_arg%now\ <= \$19078_modulo6684356_arg%next\;
        \$v5103%now\ <= \$v5103%next\;
        \$19522%now\ <= \$19522%next\;
        \$19544%now\ <= \$19544%next\;
        \$19243%now\ <= \$19243%next\;
        \$19718%now\ <= \$19718%next\;
        \$19148_modulo6684357_arg%now\ <= \$19148_modulo6684357_arg%next\;
        \$19538%now\ <= \$19538%next\;
        \$19255%now\ <= \$19255%next\;
        \$v4571%now\ <= \$v4571%next\;
        \$19275%now\ <= \$19275%next\;
        \$19281%now\ <= \$19281%next\;
        \$18599_hd%now\ <= \$18599_hd%next\;
        \$19836%now\ <= \$19836%next\;
        \$v4872%now\ <= \$v4872%next\;
        \$19043_modulo6684349_id%now\ <= \$19043_modulo6684349_id%next\;
        \$19884%now\ <= \$19884%next\;
        \$19871%now\ <= \$19871%next\;
        \$18851%now\ <= \$18851%next\;
        \$19557%now\ <= \$19557%next\;
        \$19517%now\ <= \$19517%next\;
        \$19532_forever6704350_id%now\ <= \$19532_forever6704350_id%next\;
        \$18782%now\ <= \$18782%next\;
        \$18526_aux664_id%now\ <= \$18526_aux664_id%next\;
        \$v4696%now\ <= \$v4696%next\;
        \$19238_w6514383_id%now\ <= \$19238_w6514383_id%next\;
        \$19582%now\ <= \$19582%next\;
        \$v5344%now\ <= \$v5344%next\;
        \$19570%now\ <= \$19570%next\;
        \$v4619%now\ <= \$v4619%next\;
        \$19888%now\ <= \$19888%next\;
        \$18794_apply638_id%now\ <= \$18794_apply638_id%next\;
        \$19497_loop666_id%now\ <= \$19497_loop666_id%next\;
        \$v4651%now\ <= \$v4651%next\;
        \$18521_loop666_result%now\ <= \$18521_loop666_result%next\;
        \$19901%now\ <= \$19901%next\;
        \$18442_cy%now\ <= \$18442_cy%next\;
        \$19444%now\ <= \$19444%next\;
        \$18549%now\ <= \$18549%next\;
        \$v5468%now\ <= \$v5468%next\;
        \$18604%now\ <= \$18604%next\;
        \$18540%now\ <= \$18540%next\;
        \$18575%now\ <= \$18575%next\;
        \$19330_compare6444359_id%now\ <= \$19330_compare6444359_id%next\;
        \$19085_modulo6684357_arg%now\ <= \$19085_modulo6684357_arg%next\;
        \$19040_modulo6684356_result%now\ <= \$19040_modulo6684356_result%next\;
        \$19324_f0%now\ <= \$19324_f0%next\;
        \$v5083%now\ <= \$v5083%next\;
        \$19540%now\ <= \$19540%next\;
        \$v5817%now\ <= \$v5817%next\;
        \$19554%now\ <= \$19554%next\;
        \$19295%now\ <= \$19295%next\;
        \$19120_res%now\ <= \$19120_res%next\;
        \$18475%now\ <= \$18475%next\;
        \$18580%now\ <= \$18580%next\;
        \$v4612%now\ <= \$v4612%next\;
        \$19005_modulo6684349_arg%now\ <= \$19005_modulo6684349_arg%next\;
        \$v4518%now\ <= \$v4518%next\;
        \$v5637%now\ <= \$v5637%next\;
        \$18848%now\ <= \$18848%next\;
        \$19801%now\ <= \$19801%next\;
        \$18893_v%now\ <= \$18893_v%next\;
        \$19913%now\ <= \$19913%next\;
        \$19262_forever6704385_id%now\ <= \$19262_forever6704385_id%next\;
        \$19210_res%now\ <= \$19210_res%next\;
        \$v5169%now\ <= \$v5169%next\;
        \$18514%now\ <= \$18514%next\;
        \$18747%now\ <= \$18747%next\;
        \$v5402%now\ <= \$v5402%next\;
        \$v5090%now\ <= \$v5090%next\;
        \$v4408%now\ <= \$v4408%next\;
        \$19304%now\ <= \$19304%next\;
        \$v5523%now\ <= \$v5523%next\;
        \$18505%now\ <= \$18505%next\;
        \$18888_next_acc%now\ <= \$18888_next_acc%next\;
        \$19376_b%now\ <= \$19376_b%next\;
        \$18688%now\ <= \$18688%next\;
        \$19100_modulo6684349_arg%now\ <= \$19100_modulo6684349_arg%next\;
        \$19412_sp%now\ <= \$19412_sp%next\;
        \$v4407%now\ <= \$v4407%next\;
        \$v5447%now\ <= \$v5447%next\;
        \$19798%now\ <= \$19798%next\;
        \$v5003%now\ <= \$v5003%next\;
        \$v5873%now\ <= \$v5873%next\;
        \$19097_modulo6684356_arg%now\ <= \$19097_modulo6684356_arg%next\;
        \$v5550%now\ <= \$v5550%next\;
        \$19626%now\ <= \$19626%next\;
        \$19471%now\ <= \$19471%next\;
        \$18721%now\ <= \$18721%next\;
        \$18971_modulo6684357_id%now\ <= \$18971_modulo6684357_id%next\;
        \$18797_branch_if648_id%now\ <= \$18797_branch_if648_id%next\;
        \$v4704%now\ <= \$v4704%next\;
        \$19288_v%now\ <= \$19288_v%next\;
        \$v5390%now\ <= \$v5390%next\;
        \$19366_compbranch6504391_result%now\ <= \$19366_compbranch6504391_result%next\;
        \$v5462%now\ <= \$v5462%next\;
        \$19914%now\ <= \$19914%next\;
        \$v5311%now\ <= \$v5311%next\;
        \$18608%now\ <= \$18608%next\;
        \$19317%now\ <= \$19317%next\;
        \$19141_modulo6684356_result%now\ <= \$19141_modulo6684356_result%next\;
        \$18511%now\ <= \$18511%next\;
        \$v4671%now\ <= \$v4671%next\;
        \$19487%now\ <= \$19487%next\;
        \$18522_loop665_arg%now\ <= \$18522_loop665_arg%next\;
        \$v4420%now\ <= \$v4420%next\;
        \$19625%now\ <= \$19625%next\;
        \$v5576%now\ <= \$v5576%next\;
        \$19886%now\ <= \$19886%next\;
        \$v5482%now\ <= \$v5482%next\;
        \result4928%now\ <= \result4928%next\;
        \$19773%now\ <= \$19773%next\;
        \$v4424%now\ <= \$v4424%next\;
        \$19787%now\ <= \$19787%next\;
        \$19104_modulo6684357_result%now\ <= \$19104_modulo6684357_result%next\;
        \$v5769%now\ <= \$v5769%next\;
        \$19496_aux664_result%now\ <= \$19496_aux664_result%next\;
        \$19717%now\ <= \$19717%next\;
        \$18647%now\ <= \$18647%next\;
        \$19155%now\ <= \$19155%next\;
        \$18661%now\ <= \$18661%next\;
        \$v4587%now\ <= \$v4587%next\;
        \$19939%now\ <= \$19939%next\;
        \$18832_v%now\ <= \$18832_v%next\;
        \$19227%now\ <= \$19227%next\;
        \$19650%now\ <= \$19650%next\;
        \$18495%now\ <= \$18495%next\;
        \$18551%now\ <= \$18551%next\;
        \$v5658%now\ <= \$v5658%next\;
        \$19276%now\ <= \$19276%next\;
        \$19859%now\ <= \$19859%next\;
        \$19325%now\ <= \$19325%next\;
        \$18977_binop_int6434365_result%now\ <= \$18977_binop_int6434365_result%next\;
        \$18944_r%now\ <= \$18944_r%next\;
        \$18527%now\ <= \$18527%next\;
        \$19119_v%now\ <= \$19119_v%next\;
        \$18648%now\ <= \$18648%next\;
        \$19793%now\ <= \$19793%next\;
        \$18877_v%now\ <= \$18877_v%next\;
        \$18939_binop_int6434363_id%now\ <= \$18939_binop_int6434363_id%next\;
        \$v5673%now\ <= \$v5673%next\;
        \$19190_binop_compare6454380_id%now\ <= \$19190_binop_compare6454380_id%next\;
        \$19842%now\ <= \$19842%next\;
        \$19144_modulo6684349_id%now\ <= \$19144_modulo6684349_id%next\;
        \$v5536%now\ <= \$v5536%next\;
        \$v5299%now\ <= \$v5299%next\;
        \$19601_copy_root_in_ram6634352_arg%now\ <= \$19601_copy_root_in_ram6634352_arg%next\;
        \$18539%now\ <= \$18539%next\;
        \$18936_modulo6684349_id%now\ <= \$18936_modulo6684349_id%next\;
        \$19015_binop_int6434367_result%now\ <= \$19015_binop_int6434367_result%next\;
        \$19171_compare6444358_id%now\ <= \$19171_compare6444358_id%next\;
        \$19597%now\ <= \$19597%next\;
        \$19581%now\ <= \$19581%next\;
        \$v4338%now\ <= \$v4338%next\;
        \$19384_compare6444359_result%now\ <= \$19384_compare6444359_result%next\;
        \$19748%now\ <= \$19748%next\;
        \$18522_loop665_id%now\ <= \$18522_loop665_id%next\;
        \$18461%now\ <= \$18461%next\;
        \$19256_v%now\ <= \$19256_v%next\;
        \$v5206%now\ <= \$v5206%next\;
        \$18824_v%now\ <= \$18824_v%next\;
        \$v5059%now\ <= \$v5059%next\;
        \$18657%now\ <= \$18657%next\;
        \$v5026%now\ <= \$v5026%next\;
        \$v4996%now\ <= \$v4996%next\;
        \$v5036%now\ <= \$v5036%next\;
        \$18825%now\ <= \$18825%next\;
        \$18806%now\ <= \$18806%next\;
        \$v4866%now\ <= \$v4866%next\;
        \$v4647%now\ <= \$v4647%next\;
        \$18891%now\ <= \$18891%next\;
        \$18843%now\ <= \$18843%next\;
        \$v4330%now\ <= \$v4330%next\;
        \$19370_compare6444359_id%now\ <= \$19370_compare6444359_id%next\;
        \$19601_copy_root_in_ram6634352_id%now\ <= \$19601_copy_root_in_ram6634352_id%next\;
        \$v5281%now\ <= \$v5281%next\;
        \$v4546%now\ <= \$v4546%next\;
        \$v4779%now\ <= \$v4779%next\;
        \$v4636%now\ <= \$v4636%next\;
        \$v4812%now\ <= \$v4812%next\;
        \$v5574%now\ <= \$v5574%next\;
        \$18526_aux664_arg%now\ <= \$18526_aux664_arg%next\;
        \$19308_v%now\ <= \$19308_v%next\;
        \$18793_make_block579_arg%now\ <= \$18793_make_block579_arg%next\;
        \$18437_loop666_arg%now\ <= \$18437_loop666_arg%next\;
        \$19206_binop_compare6454382_result%now\ <= \$19206_binop_compare6454382_result%next\;
        \$18444%now\ <= \$18444%next\;
        \$19066_modulo6684357_id%now\ <= \$19066_modulo6684357_id%next\;
        \$19046_r%now\ <= \$19046_r%next\;
        \$19837%now\ <= \$19837%next\;
        \$v5429%now\ <= \$v5429%next\;
        \$19571%now\ <= \$19571%next\;
        \$v4978%now\ <= \$v4978%next\;
        \$v4920%now\ <= \$v4920%next\;
        \$v5799%now\ <= \$v5799%next\;
        \$18524_loop666_arg%now\ <= \$18524_loop666_arg%next\;
        \$18810%now\ <= \$18810%next\;
        \$19944%now\ <= \$19944%next\;
        \$18880%now\ <= \$18880%next\;
        \$18869%now\ <= \$18869%next\;
        \$v5490%now\ <= \$v5490%next\;
        \$18659%now\ <= \$18659%next\;
        \$v5257%now\ <= \$v5257%next\;
        \$18945_modulo6684356_id%now\ <= \$18945_modulo6684356_id%next\;
        \$18683_hd%now\ <= \$18683_hd%next\;
        \$v4428%now\ <= \$v4428%next\;
        \$v5055%now\ <= \$v5055%next\;
        \$19774%now\ <= \$19774%next\;
        \$v5522%now\ <= \$v5522%next\;
        \$19783%now\ <= \$19783%next\;
        \$19125_modulo6684349_result%now\ <= \$19125_modulo6684349_result%next\;
        \$19097_modulo6684356_id%now\ <= \$19097_modulo6684356_id%next\;
        \$19507_next%now\ <= \$19507_next%next\;
        \rdy4400%now\ <= \rdy4400%next\;
        \$19542%now\ <= \$19542%next\;
        \$v5042%now\ <= \$v5042%next\;
        \$18813%now\ <= \$18813%next\;
        \$19220%now\ <= \$19220%next\;
        \$v4667%now\ <= \$v4667%next\;
        \$v4678%now\ <= \$v4678%next\;
        \$19211_compare6444358_result%now\ <= \$19211_compare6444358_result%next\;
        \$18790_loop666_result%now\ <= \$18790_loop666_result%next\;
        \$19804%now\ <= \$19804%next\;
        \$18622%now\ <= \$18622%next\;
        \$v4519%now\ <= \$v4519%next\;
        \$19667%now\ <= \$19667%next\;
        \$v4593%now\ <= \$v4593%next\;
        \$19811_copy_root_in_ram6634341_arg%now\ <= \$19811_copy_root_in_ram6634341_arg%next\;
        \$18695%now\ <= \$18695%next\;
        \$19789_next%now\ <= \$19789_next%next\;
        \$19259%now\ <= \$19259%next\;
        \$18437_loop666_id%now\ <= \$18437_loop666_id%next\;
        \$19203_compare6444358_id%now\ <= \$19203_compare6444358_id%next\;
        \$19788%now\ <= \$19788%next\;
        \$19141_modulo6684356_arg%now\ <= \$19141_modulo6684356_arg%next\;
        \$18473%now\ <= \$18473%next\;
        \$v5134%now\ <= \$v5134%next\;
        \$19144_modulo6684349_result%now\ <= \$19144_modulo6684349_result%next\;
        \$19932%now\ <= \$19932%next\;
        \$18603%now\ <= \$18603%next\;
        \$v5365%now\ <= \$v5365%next\;
        \$19701%now\ <= \$19701%next\;
        \$19543%now\ <= \$19543%next\;
        \$v5168%now\ <= \$v5168%next\;
        \$v4529%now\ <= \$v4529%next\;
        \$v4839%now\ <= \$v4839%next\;
        \$v4679%now\ <= \$v4679%next\;
        \$19796%now\ <= \$19796%next\;
        \$18845%now\ <= \$18845%next\;
        \$v5233%now\ <= \$v5233%next\;
        \$18438_loop665_arg%now\ <= \$18438_loop665_arg%next\;
        \$19337_compare6444359_arg%now\ <= \$19337_compare6444359_arg%next\;
        \$v4632%now\ <= \$v4632%next\;
        \$v4957%now\ <= \$v4957%next\;
        \$19336_b%now\ <= \$19336_b%next\;
        \$19709%now\ <= \$19709%next\;
        \$19031_modulo6684349_result%now\ <= \$19031_modulo6684349_result%next\;
        \$19824_hd%now\ <= \$19824_hd%next\;
        \$19619%now\ <= \$19619%next\;
        \$18546%now\ <= \$18546%next\;
        \$v5872%now\ <= \$v5872%next\;
        \$19818%now\ <= \$19818%next\;
        \$18971_modulo6684357_arg%now\ <= \$18971_modulo6684357_arg%next\;
        \$v4502%now\ <= \$v4502%next\;
        \$19326_compbranch6504387_id%now\ <= \$19326_compbranch6504387_id%next\;
        \$18531%now\ <= \$18531%next\;
        \$v4802%now\ <= \$v4802%next\;
        \$18841%now\ <= \$18841%next\;
        \$v4639%now\ <= \$v4639%next\;
        \$19466_sp%now\ <= \$19466_sp%next\;
        \$18567%now\ <= \$18567%next\;
        \$v4683%now\ <= \$v4683%next\;
        \$19643_w%now\ <= \$19643_w%next\;
        \$18649%now\ <= \$18649%next\;
        \$18929_modulo6684349_arg%now\ <= \$18929_modulo6684349_arg%next\;
        \$v5184%now\ <= \$v5184%next\;
        \$v4335%now\ <= \$v4335%next\;
        \$v5915%now\ <= \$v5915%next\;
        \$19169_v%now\ <= \$19169_v%next\;
        \$v5487%now\ <= \$v5487%next\;
        \$v5552%now\ <= \$v5552%next\;
        \$19361_fill6544390_id%now\ <= \$19361_fill6544390_id%next\;
        \$v5811%now\ <= \$v5811%next\;
        \$19512%now\ <= \$19512%next\;
        \$v4471%now\ <= \$v4471%next\;
        \$19725%now\ <= \$19725%next\;
        \$19844%now\ <= \$19844%next\;
        \$18732%now\ <= \$18732%next\;
        \$18618%now\ <= \$18618%next\;
        \$19387_compbranch6504394_arg%now\ <= \$19387_compbranch6504394_arg%next\;
        \$19027_r%now\ <= \$19027_r%next\;
        \$v5471%now\ <= \$v5471%next\;
        \$19659_hd%now\ <= \$19659_hd%next\;
        \$19875%now\ <= \$19875%next\;
        \$19639%now\ <= \$19639%next\;
        \$18470%now\ <= \$18470%next\;
        \$19310%now\ <= \$19310%next\;
        \$19815%now\ <= \$19815%next\;
        \$v5696%now\ <= \$v5696%next\;
        \$19350_v%now\ <= \$19350_v%next\;
        \$19503%now\ <= \$19503%next\;
        \$19182_binop_compare6454379_result%now\ <= \$19182_binop_compare6454379_result%next\;
        \$18955_modulo6684349_result%now\ <= \$18955_modulo6684349_result%next\;
        \$18476%now\ <= \$18476%next\;
        \$18443%now\ <= \$18443%next\;
        \$19230_v%now\ <= \$19230_v%next\;
        \$19018_v%now\ <= \$19018_v%next\;
        \$19713%now\ <= \$19713%next\;
        \$19218_v%now\ <= \$19218_v%next\;
        \$19009_modulo6684357_arg%now\ <= \$19009_modulo6684357_arg%next\;
        \$19498_loop665_result%now\ <= \$19498_loop665_result%next\;
        \$v5198%now\ <= \$v5198%next\;
        \$19741%now\ <= \$19741%next\;
        \$v4581%now\ <= \$v4581%next\;
        \$19161%now\ <= \$19161%next\;
        \$19156%now\ <= \$19156%next\;
        \$19104_modulo6684357_arg%now\ <= \$19104_modulo6684357_arg%next\;
        \$18492%now\ <= \$18492%next\;
        \$v5571%now\ <= \$v5571%next\;
        \$v4615%now\ <= \$v4615%next\;
        \$19937%now\ <= \$19937%next\;
        \$18917_modulo6684349_arg%now\ <= \$18917_modulo6684349_arg%next\;
        \$v5384%now\ <= \$v5384%next\;
        \$18939_binop_int6434363_arg%now\ <= \$18939_binop_int6434363_arg%next\;
        \$19572%now\ <= \$19572%next\;
        \$18898%now\ <= \$18898%next\;
        \$19391_compare6444359_result%now\ <= \$19391_compare6444359_result%next\;
        \$v5563%now\ <= \$v5563%next\;
        \$18948_modulo6684349_id%now\ <= \$18948_modulo6684349_id%next\;
        \$v5897%now\ <= \$v5897%next\;
        \$19100_modulo6684349_id%now\ <= \$19100_modulo6684349_id%next\;
        \$19409_sp%now\ <= \$19409_sp%next\;
        \$18478%now\ <= \$18478%next\;
        \$19047_modulo6684357_result%now\ <= \$19047_modulo6684357_result%next\;
        \$19009_modulo6684357_result%now\ <= \$19009_modulo6684357_result%next\;
        \$v5072%now\ <= \$v5072%next\;
        \$18895_v%now\ <= \$18895_v%next\;
        \$18559_copy_root_in_ram6634347_id%now\ <= \$18559_copy_root_in_ram6634347_id%next\;
        \$18559_copy_root_in_ram6634347_arg%now\ <= \$18559_copy_root_in_ram6634347_arg%next\;
        \$19922%now\ <= \$19922%next\;
        \$19125_modulo6684349_id%now\ <= \$19125_modulo6684349_id%next\;
        \$18629%now\ <= \$18629%next\;
        \$v4887%now\ <= \$v4887%next\;
        \$v4556%now\ <= \$v4556%next\;
        \$v5453%now\ <= \$v5453%next\;
        \$19731%now\ <= \$19731%next\;
        \$19449%now\ <= \$19449%next\;
        \$18669%now\ <= \$18669%next\;
        \$18660%now\ <= \$18660%next\;
        \rdy4573%now\ <= \rdy4573%next\;
        \$18795_offsetclosure_n639_id%now\ <= \$18795_offsetclosure_n639_id%next\;
        \$19401_compbranch6504396_arg%now\ <= \$19401_compbranch6504396_arg%next\;
        \$19878%now\ <= \$19878%next\;
        \$v5066%now\ <= \$v5066%next\;
        \$18631%now\ <= \$18631%next\;
        \$v4327%now\ <= \$v4327%next\;
        \$19234_sp%now\ <= \$19234_sp%next\;
        \$18687%now\ <= \$18687%next\;
        \$19811_copy_root_in_ram6634341_result%now\ <= \$19811_copy_root_in_ram6634341_result%next\;
        \rdy4608%now\ <= \rdy4608%next\;
        \$19728%now\ <= \$19728%next\;
        \$v5492%now\ <= \$v5492%next\;
        \$19843%now\ <= \$19843%next\;
        \$19532_forever6704350_arg%now\ <= \$19532_forever6704350_arg%next\;
        \$19028_modulo6684357_id%now\ <= \$19028_modulo6684357_id%next\;
        \$18958_binop_int6434364_arg%now\ <= \$18958_binop_int6434364_arg%next\;
        \$v4700%now\ <= \$v4700%next\;
        \$19301_v%now\ <= \$19301_v%next\;
        \$v4940%now\ <= \$v4940%next\;
        \$19012_modulo6684349_result%now\ <= \$19012_modulo6684349_result%next\;
        \$19268%now\ <= \$19268%next\;
        \$19772%now\ <= \$19772%next\;
        \$19226%now\ <= \$19226%next\;
        \$v5727%now\ <= \$v5727%next\;
        \$18889_v%now\ <= \$18889_v%next\;
        \$19882%now\ <= \$19882%next\;
        \$19877%now\ <= \$19877%next\;
        \$19091_binop_int6434371_id%now\ <= \$19091_binop_int6434371_id%next\;
        \$v4796%now\ <= \$v4796%next\;
        \$18907_modulo6684356_result%now\ <= \$18907_modulo6684356_result%next\;
        \$19561%now\ <= \$19561%next\;
        \$19282_v%now\ <= \$19282_v%next\;
        \$19806%now\ <= \$19806%next\;
        \$19257_v%now\ <= \$19257_v%next\;
        \$19660%now\ <= \$19660%next\;
        \$18583_w%now\ <= \$18583_w%next\;
        \$v4818%now\ <= \$v4818%next\;
        \$v4750%now\ <= \$v4750%next\;
        \$19492%now\ <= \$19492%next\;
        \$18525_loop665_id%now\ <= \$18525_loop665_id%next\;
        \$19311%now\ <= \$19311%next\;
        \$19743%now\ <= \$19743%next\;
        \$v4775%now\ <= \$v4775%next\;
        \$v4713%now\ <= \$v4713%next\;
        \$19519%now\ <= \$19519%next\;
        \$19870%now\ <= \$19870%next\;
        \$v4540%now\ <= \$v4540%next\;
        \$19638%now\ <= \$19638%next\;
        \$v4821%now\ <= \$v4821%next\;
        \$v5664%now\ <= \$v5664%next\;
        \$19211_compare6444358_arg%now\ <= \$19211_compare6444358_arg%next\;
        \$18500%now\ <= \$18500%next\;
        \$18545_next%now\ <= \$18545_next%next\;
        \$19078_modulo6684356_result%now\ <= \$19078_modulo6684356_result%next\;
        \$19868%now\ <= \$19868%next\;
        \$19047_modulo6684357_id%now\ <= \$19047_modulo6684357_id%next\;
        \$18663%now\ <= \$18663%next\;
        \$18679%now\ <= \$18679%next\;
        \$19053_binop_int6434369_result%now\ <= \$19053_binop_int6434369_result%next\;
        \$v4937%now\ <= \$v4937%next\;
        \$v5305%now\ <= \$v5305%next\;
        \$18986_modulo6684349_result%now\ <= \$18986_modulo6684349_result%next\;
        \$19266%now\ <= \$19266%next\;
        \$19447_sp%now\ <= \$19447_sp%next\;
        \$19084_r%now\ <= \$19084_r%next\;
        \$19779_loop666_result%now\ <= \$19779_loop666_result%next\;
        \$v5825%now\ <= \$v5825%next\;
        \$18464_rdy%now\ <= \$18464_rdy%next\;
        \$19636%now\ <= \$19636%next\;
        \$19329_b%now\ <= \$19329_b%next\;
        \$v5596%now\ <= \$v5596%next\;
        \$19031_modulo6684349_id%now\ <= \$19031_modulo6684349_id%next\;
        \$19526_forever6704355_id%now\ <= \$19526_forever6704355_id%next\;
        \$19926%now\ <= \$19926%next\;
        \$19614_hd%now\ <= \$19614_hd%next\;
        \$19594%now\ <= \$19594%next\;
        \$18542_next%now\ <= \$18542_next%next\;
        \$18553_forever6704348_id%now\ <= \$18553_forever6704348_id%next\;
        \$19521%now\ <= \$19521%next\;
        \$19832%now\ <= \$19832%next\;
        \$v4455%now\ <= \$v4455%next\;
        \$v4640%now\ <= \$v4640%next\;
        \$19053_binop_int6434369_arg%now\ <= \$19053_binop_int6434369_arg%next\;
        \$18508%now\ <= \$18508%next\;
        \$19684%now\ <= \$19684%next\;
        \$19315%now\ <= \$19315%next\;
        \$19166_binop_compare6454377_id%now\ <= \$19166_binop_compare6454377_id%next\;
        \$19110%now\ <= \$19110%next\;
        \$19678%now\ <= \$19678%next\;
        \$v5405%now\ <= \$v5405%next\;
        \$v5622%now\ <= \$v5622%next\;
        \$v5188%now\ <= \$v5188%next\;
        \$v5138%now\ <= \$v5138%next\;
        \$19198_binop_compare6454381_result%now\ <= \$19198_binop_compare6454381_result%next\;
        \$v4972%now\ <= \$v4972%next\;
        \$19872%now\ <= \$19872%next\;
        \$19031_modulo6684349_arg%now\ <= \$19031_modulo6684349_arg%next\;
        \$19405_compare6444359_arg%now\ <= \$19405_compare6444359_arg%next\;
        \$v4754%now\ <= \$v4754%next\;
        \$v5254%now\ <= \$v5254%next\;
        \$v5275%now\ <= \$v5275%next\;
        \$18642%now\ <= \$18642%next\;
        \$19892%now\ <= \$19892%next\;
        \$v4339%now\ <= \$v4339%next\;
        \$v4532%now\ <= \$v4532%next\;
        \$v5260%now\ <= \$v5260%next\;
        \$19021_modulo6684356_arg%now\ <= \$19021_modulo6684356_arg%next\;
        \$18996_binop_int6434366_result%now\ <= \$18996_binop_int6434366_result%next\;
        \$19005_modulo6684349_id%now\ <= \$19005_modulo6684349_id%next\;
        \$18522_loop665_result%now\ <= \$18522_loop665_result%next\;
        \$18682_w%now\ <= \$18682_w%next\;
        \$18914_modulo6684357_id%now\ <= \$18914_modulo6684357_id%next\;
        \$18673%now\ <= \$18673%next\;
        \$19766%now\ <= \$19766%next\;
        \$v4558%now\ <= \$v4558%next\;
        \$19214%now\ <= \$19214%next\;
        \$19566%now\ <= \$19566%next\;
        \$v4337%now\ <= \$v4337%next\;
        \$v5096%now\ <= \$v5096%next\;
        \$v5359%now\ <= \$v5359%next\;
        \$19174_binop_compare6454378_result%now\ <= \$19174_binop_compare6454378_result%next\;
        \$19563%now\ <= \$19563%next\;
        \$v4606%now\ <= \$v4606%next\;
        \$v5141%now\ <= \$v5141%next\;
        \$18639%now\ <= \$18639%next\;
        \$19154%now\ <= \$19154%next\;
        \$18562%now\ <= \$18562%next\;
        \$v4449%now\ <= \$v4449%next\;
        \$v4605%now\ <= \$v4605%next\;
        \$v4539%now\ <= \$v4539%next\;
        \$18666%now\ <= \$18666%next\;
        \$19781_aux664_id%now\ <= \$19781_aux664_id%next\;
        \$18904_v%now\ <= \$18904_v%next\;
        \$18498%now\ <= \$18498%next\;
        \$v4562%now\ <= \$v4562%next\;
        \$19497_loop666_arg%now\ <= \$19497_loop666_arg%next\;
        \$18564%now\ <= \$18564%next\;
        \$v5335%now\ <= \$v5335%next\;
        \$19834%now\ <= \$19834%next\;
        \$19700%now\ <= \$19700%next\;
        \$19769%now\ <= \$19769%next\;
        \$19907%now\ <= \$19907%next\;
        \$18724%now\ <= \$18724%next\;
        \$19425%now\ <= \$19425%next\;
        \$19293%now\ <= \$19293%next\;
        \$19147_r%now\ <= \$19147_r%next\;
        \$19950%now\ <= \$19950%next\;
        \$19355%now\ <= \$19355%next\;
        \$19024_modulo6684349_id%now\ <= \$19024_modulo6684349_id%next\;
        \$19665%now\ <= \$19665%next\;
        \$19351%now\ <= \$19351%next\;
        \$19500%now\ <= \$19500%next\;
        \$v4833%now\ <= \$v4833%next\;
        \$v4791%now\ <= \$v4791%next\;
        \$v4746%now\ <= \$v4746%next\;
        \$v5524%now\ <= \$v5524%next\;
        \$19856%now\ <= \$19856%next\;
        \$18456%now\ <= \$18456%next\;
        \$19021_modulo6684356_result%now\ <= \$19021_modulo6684356_result%next\;
        \$v5560%now\ <= \$v5560%next\;
        \$v4751%now\ <= \$v4751%next\;
        \$18487%now\ <= \$18487%next\;
        \$19755%now\ <= \$19755%next\;
        \$19233%now\ <= \$19233%next\;
        \$18654%now\ <= \$18654%next\;
        \$v4911%now\ <= \$v4911%next\;
        \$v5743%now\ <= \$v5743%next\;
        \$19414%now\ <= \$19414%next\;
        \$19649%now\ <= \$19649%next\;
        \$18702%now\ <= \$18702%next\;
        \$18897%now\ <= \$18897%next\;
        \$v4496%now\ <= \$v4496%next\;
        \$18967_modulo6684349_result%now\ <= \$18967_modulo6684349_result%next\;
        \$v5477%now\ <= \$v5477%next\;
        \$v4675%now\ <= \$v4675%next\;
        \$v5107%now\ <= \$v5107%next\;
        \$19485%now\ <= \$19485%next\;
        \$v5597%now\ <= \$v5597%next\;
        \$19132_modulo6684349_arg%now\ <= \$19132_modulo6684349_arg%next\;
        \$18781%now\ <= \$18781%next\;
        \$19252_forever6704384_id%now\ <= \$19252_forever6704384_id%next\;
        \$v4984%now\ <= \$v4984%next\;
        \$v5753%now\ <= \$v5753%next\;
        \$18896_v%now\ <= \$18896_v%next\;
        \$18737%now\ <= \$18737%next\;
        \$18439_wait662_result%now\ <= \$18439_wait662_result%next\;
        \$v5102%now\ <= \$v5102%next\;
        \$v4813%now\ <= \$v4813%next\;
        \$v5432%now\ <= \$v5432%next\;
        \$19642%now\ <= \$19642%next\;
        \$18446_dur%now\ <= \$18446_dur%next\;
        \$18625_copy_root_in_ram6634345_id%now\ <= \$18625_copy_root_in_ram6634345_id%next\;
        \$v5314%now\ <= \$v5314%next\;
        \$v5540%now\ <= \$v5540%next\;
        \$19617%now\ <= \$19617%next\;
        \$19451%now\ <= \$19451%next\;
        \$18556_forever6704344_id%now\ <= \$18556_forever6704344_id%next\;
        \$19585%now\ <= \$19585%next\;
        \$18886%now\ <= \$18886%next\;
        \$18439_wait662_id%now\ <= \$18439_wait662_id%next\;
        \$v5441%now\ <= \$v5441%next\;
        \$19737%now\ <= \$19737%next\;
        \$19879%now\ <= \$19879%next\;
        \$19072_binop_int6434370_id%now\ <= \$19072_binop_int6434370_id%next\;
        \$19462%now\ <= \$19462%next\;
        \$18516%now\ <= \$18516%next\;
        \$18838_v%now\ <= \$18838_v%next\;
        \$v5502%now\ <= \$v5502%next\;
        \$v5814%now\ <= \$v5814%next\;
        \$v5845%now\ <= \$v5845%next\;
        \$18438_loop665_result%now\ <= \$18438_loop665_result%next\;
        \$19658_w%now\ <= \$19658_w%next\;
        \$19182_binop_compare6454379_arg%now\ <= \$19182_binop_compare6454379_arg%next\;
        \$18901_binop_int6434361_result%now\ <= \$18901_binop_int6434361_result%next\;
        \$18453%now\ <= \$18453%next\;
        \$19260%now\ <= \$19260%next\;
        \$v5605%now\ <= \$v5605%next\;
        \$18971_modulo6684357_result%now\ <= \$18971_modulo6684357_result%next\;
        \$19853%now\ <= \$19853%next\;
        \$v5131%now\ <= \$v5131%next\;
        \$18820_v%now\ <= \$18820_v%next\;
        \$18571_copy_root_in_ram6634345_result%now\ <= \$18571_copy_root_in_ram6634345_result%next\;
        \$18515%now\ <= \$18515%next\;
        \$v4689%now\ <= \$v4689%next\;
        \$18914_modulo6684357_result%now\ <= \$18914_modulo6684357_result%next\;
        \$v5497%now\ <= \$v5497%next\;
        \$19951%now\ <= \$19951%next\;
        \$19807%now\ <= \$19807%next\;
        \$19241_v%now\ <= \$19241_v%next\;
        \$19242%now\ <= \$19242%next\;
        \$19539%now\ <= \$19539%next\;
        \$18752%now\ <= \$18752%next\;
        \$v5544%now\ <= \$v5544%next\;
        \result4607%now\ <= \result4607%next\;
        \$19091_binop_int6434371_arg%now\ <= \$19091_binop_int6434371_arg%next\;
        \$19345%now\ <= \$19345%next\;
        \$v5491%now\ <= \$v5491%next\;
        \$18844%now\ <= \$18844%next\;
        \$18963_r%now\ <= \$18963_r%next\;
        \$v5652%now\ <= \$v5652%next\;
        \$v5876%now\ <= \$v5876%next\;
        \$19113_forever6704372_id%now\ <= \$19113_forever6704372_id%next\;
        \$19383_b%now\ <= \$19383_b%next\;
        \$19584%now\ <= \$19584%next\;
        \$19942%now\ <= \$19942%next\;
        \$19615%now\ <= \$19615%next\;
        \$18676%now\ <= \$18676%next\;
        \$v4514%now\ <= \$v4514%next\;
        \$19316%now\ <= \$19316%next\;
        \$19148_modulo6684357_id%now\ <= \$19148_modulo6684357_id%next\;
        \$v4492%now\ <= \$v4492%next\;
        \$v5347%now\ <= \$v5347%next\;
        \$v5411%now\ <= \$v5411%next\;
        \$18756%now\ <= \$18756%next\;
        \$19865_w%now\ <= \$19865_w%next\;
        \$18533%now\ <= \$18533%next\;
        \$19297_v%now\ <= \$19297_v%next\;
        \$18497%now\ <= \$18497%next\;
        \$19062_modulo6684349_arg%now\ <= \$19062_modulo6684349_arg%next\;
        \$19456%now\ <= \$19456%next\;
        \$v5909%now\ <= \$v5909%next\;
        \$v5356%now\ <= \$v5356%next\;
        \$v5584%now\ <= \$v5584%next\;
        \$v5023%now\ <= \$v5023%next\;
        \$18766%now\ <= \$18766%next\;
        \$19770%now\ <= \$19770%next\;
        \$v4960%now\ <= \$v4960%next\;
        \$18674%now\ <= \$18674%next\;
        \$18595%now\ <= \$18595%next\;
        \$19927%now\ <= \$19927%next\;
        \$v5293%now\ <= \$v5293%next\;
        \$v5525%now\ <= \$v5525%next\;
        \$18786%now\ <= \$18786%next\;
        \$19592%now\ <= \$19592%next\;
        \$18748%now\ <= \$18748%next\;
        \$18448_dis%now\ <= \$18448_dis%next\;
        \$19398_compare6444359_result%now\ <= \$19398_compare6444359_result%next\;
        \$19202_res%now\ <= \$19202_res%next\;
        \$18951_r%now\ <= \$18951_r%next\;
        \$19040_modulo6684356_arg%now\ <= \$19040_modulo6684356_arg%next\;
        \$v5724%now\ <= \$v5724%next\;
        \$18780%now\ <= \$18780%next\;
        \$18651%now\ <= \$18651%next\;
        \$19518_next%now\ <= \$19518_next%next\;
        \$19005_modulo6684349_result%now\ <= \$19005_modulo6684349_result%next\;
        \$18808%now\ <= \$18808%next\;
        \$18715%now\ <= \$18715%next\;
        \$19799%now\ <= \$19799%next\;
        \$v5505%now\ <= \$v5505%next\;
        \$v5867%now\ <= \$v5867%next\;
        \$19646%now\ <= \$19646%next\;
        \$19833%now\ <= \$19833%next\;
        \$19182_binop_compare6454379_id%now\ <= \$19182_binop_compare6454379_id%next\;
        \$v5000%now\ <= \$v5000%next\;
        \$v5185%now\ <= \$v5185%next\;
        \$v5034%now\ <= \$v5034%next\;
        \$18467_loop665_result%now\ <= \$18467_loop665_result%next\;
        \$v5222%now\ <= \$v5222%next\;
        \$v4782%now\ <= \$v4782%next\;
        \$19547_copy_root_in_ram6634352_id%now\ <= \$19547_copy_root_in_ram6634352_id%next\;
        \$19915%now\ <= \$19915%next\;
        \$19719%now\ <= \$19719%next\;
        \$18777%now\ <= \$18777%next\;
        \$18550%now\ <= \$18550%next\;
        \$18842%now\ <= \$18842%next\;
        \$18489%now\ <= \$18489%next\;
        \$18439_wait662_arg%now\ <= \$18439_wait662_arg%next\;
        \$19100_modulo6684349_result%now\ <= \$19100_modulo6684349_result%next\;
        \$19135_binop_int6434374_id%now\ <= \$19135_binop_int6434374_id%next\;
        \$18796_make_block_n646_arg%now\ <= \$18796_make_block_n646_arg%next\;
        \$v5084%now\ <= \$v5084%next\;
        \$v4654%now\ <= \$v4654%next\;
        \$19820%now\ <= \$19820%next\;
        \$18901_binop_int6434361_arg%now\ <= \$18901_binop_int6434361_arg%next\;
        \$18701%now\ <= \$18701%next\;
        \$18768_w%now\ <= \$18768_w%next\;
        \$19586%now\ <= \$19586%next\;
        \$v5709%now\ <= \$v5709%next\;
        \$18613_copy_root_in_ram6634346_arg%now\ <= \$18613_copy_root_in_ram6634346_arg%next\;
        \$19917%now\ <= \$19917%next\;
        \$19138_v%now\ <= \$19138_v%next\;
        \$19697%now\ <= \$19697%next\;
        \$v4423%now\ <= \$v4423%next\;
        \result4963%now\ <= \result4963%next\;
        \$18794_apply638_arg%now\ <= \$18794_apply638_arg%next\;
        \$18792_wait662_arg%now\ <= \$18792_wait662_arg%next\;
        \$18741%now\ <= \$18741%next\;
        \$18735%now\ <= \$18735%next\;
        \$v5039%now\ <= \$v5039%next\;
        \$19677%now\ <= \$19677%next\;
        \$v5296%now\ <= \$v5296%next\;
        \$18714%now\ <= \$18714%next\;
        \$19231%now\ <= \$19231%next\;
        \$v5689%now\ <= \$v5689%next\;
        \$v5251%now\ <= \$v5251%next\;
        \$19876%now\ <= \$19876%next\;
        \$v5606%now\ <= \$v5606%next\;
        \$v5670%now\ <= \$v5670%next\;
        \$18794_apply638_result%now\ <= \$18794_apply638_result%next\;
        \$19921%now\ <= \$19921%next\;
        \$19420_w06554397_id%now\ <= \$19420_w06554397_id%next\;
        \$v4719%now\ <= \$v4719%next\;
        \$19059_modulo6684356_id%now\ <= \$19059_modulo6684356_id%next\;
        \$19864%now\ <= \$19864%next\;
        \$19347_fill6534389_result%now\ <= \$19347_fill6534389_result%next\;
        \$v5099%now\ <= \$v5099%next\;
        \$19860%now\ <= \$19860%next\;
        \$19781_aux664_arg%now\ <= \$19781_aux664_arg%next\;
        \$v4827%now\ <= \$v4827%next\;
        \$18964_modulo6684356_arg%now\ <= \$18964_modulo6684356_arg%next\;
        \$v5802%now\ <= \$v5802%next\;
        \$v4917%now\ <= \$v4917%next\;
        \$19302%now\ <= \$19302%next\;
        \$v5368%now\ <= \$v5368%next\;
        \$19823_w%now\ <= \$19823_w%next\;
        \$v5494%now\ <= \$v5494%next\;
        \$19668%now\ <= \$19668%next\;
        \$19398_compare6444359_id%now\ <= \$19398_compare6444359_id%next\;
        \$18574%now\ <= \$18574%next\;
        \$19228_v%now\ <= \$19228_v%next\;
        \$v5079%now\ <= \$v5079%next\;
        \$19749%now\ <= \$19749%next\;
        \$19795%now\ <= \$19795%next\;
        \$19203_compare6444358_arg%now\ <= \$19203_compare6444358_arg%next\;
        \$19768%now\ <= \$19768%next\;
        \$v4809%now\ <= \$v4809%next\;
        \$19941%now\ <= \$19941%next\;
        \$v4902%now\ <= \$v4902%next\;
        \$18899%now\ <= \$18899%next\;
        \$19605%now\ <= \$19605%next\;
        \$19514%now\ <= \$19514%next\;
        \$v4836%now\ <= \$v4836%next\;
        \$18640%now\ <= \$18640%next\;
        \$v4716%now\ <= \$v4716%next\;
        \$v5396%now\ <= \$v5396%next\;
        \$19341%now\ <= \$19341%next\;
        \$18870_v%now\ <= \$18870_v%next\;
        \$19722%now\ <= \$19722%next\;
        \$19475%now\ <= \$19475%next\;
        \$v5353%now\ <= \$v5353%next\;
        \$v4953%now\ <= \$v4953%next\;
        \$19460%now\ <= \$19460%next\;
        \$19470%now\ <= \$19470%next\;
        \$19580%now\ <= \$19580%next\;
        \$19893%now\ <= \$19893%next\;
        \$v4597%now\ <= \$v4597%next\;
        \$v5051%now\ <= \$v5051%next\;
        \$v5679%now\ <= \$v5679%next\;
        \$v5630%now\ <= \$v5630%next\;
        \$19889%now\ <= \$19889%next\;
        \$18812%now\ <= \$18812%next\;
        \$v5543%now\ <= \$v5543%next\;
        \$18955_modulo6684349_id%now\ <= \$18955_modulo6684349_id%next\;
        \$19529_forever6704351_arg%now\ <= \$19529_forever6704351_arg%next\;
        \$v5556%now\ <= \$v5556%next\;
        \$19497_loop666_result%now\ <= \$19497_loop666_result%next\;
        \$18536%now\ <= \$18536%next\;
        \$19433%now\ <= \$19433%next\;
        \$v4857%now\ <= \$v4857%next\;
        \$19286%now\ <= \$19286%next\;
        \$19621%now\ <= \$19621%next\;
        \$18758%now\ <= \$18758%next\;
        \$19261%now\ <= \$19261%next\;
        \$v5566%now\ <= \$v5566%next\;
        \$v4881%now\ <= \$v4881%next\;
        \$19148_modulo6684357_result%now\ <= \$19148_modulo6684357_result%next\;
        \$v4795%now\ <= \$v4795%next\;
        \$19945%now\ <= \$19945%next\;
        \$v4466%now\ <= \$v4466%next\;
        \$v4824%now\ <= \$v4824%next\;
        \$19747%now\ <= \$19747%next\;
        \$19081_modulo6684349_id%now\ <= \$19081_modulo6684349_id%next\;
        \$19285%now\ <= \$19285%next\;
        \$v4884%now\ <= \$v4884%next\;
        \$v5863%now\ <= \$v5863%next\;
        \$19394_compbranch6504395_result%now\ <= \$19394_compbranch6504395_result%next\;
        \$19535_copy_root_in_ram6634354_result%now\ <= \$19535_copy_root_in_ram6634354_result%next\;
        \$v4758%now\ <= \$v4758%next\;
        \$v4488%now\ <= \$v4488%next\;
        \$19012_modulo6684349_arg%now\ <= \$19012_modulo6684349_arg%next\;
        \$18607%now\ <= \$18607%next\;
        \$19753%now\ <= \$19753%next\;
        \$18785%now\ <= \$18785%next\;
        \$19394_compbranch6504395_id%now\ <= \$19394_compbranch6504395_id%next\;
        \$v5894%now\ <= \$v5894%next\;
        \$18799_w1656_arg%now\ <= \$18799_w1656_arg%next\;
        \$18856_loop_push6494360_id%now\ <= \$18856_loop_push6494360_id%next\;
        \$v4981%now\ <= \$v4981%next\;
        \$19391_compare6444359_arg%now\ <= \$19391_compare6444359_arg%next\;
        \$19366_compbranch6504391_id%now\ <= \$19366_compbranch6504391_id%next\;
        \$v4771%now\ <= \$v4771%next\;
        \$19781_aux664_result%now\ <= \$19781_aux664_result%next\;
        \$19174_binop_compare6454378_id%now\ <= \$19174_binop_compare6454378_id%next\;
        \$19416_w36574398_arg%now\ <= \$19416_w36574398_arg%next\;
        \$v5627%now\ <= \$v5627%next\;
        \$19271%now\ <= \$19271%next\;
        \$v5126%now\ <= \$v5126%next\;
        \$18708%now\ <= \$18708%next\;
        \$19780_loop665_id%now\ <= \$19780_loop665_id%next\;
        \$18827%now\ <= \$18827%next\;
        \$v5890%now\ <= \$v5890%next\;
        \$18882_v%now\ <= \$18882_v%next\;
        \$18525_loop665_arg%now\ <= \$18525_loop665_arg%next\;
        \$v5623%now\ <= \$v5623%next\;
        \$19344%now\ <= \$19344%next\;
        \$19576%now\ <= \$19576%next\;
        \$19171_compare6444358_arg%now\ <= \$19171_compare6444358_arg%next\;
        \$19838_copy_root_in_ram6634340_id%now\ <= \$19838_copy_root_in_ram6634340_id%next\;
        \$v5387%now\ <= \$v5387%next\;
        \$19373_compbranch6504392_arg%now\ <= \$19373_compbranch6504392_arg%next\;
        \$v5602%now\ <= \$v5602%next\;
        \$18544%now\ <= \$18544%next\;
        \$v5773%now\ <= \$v5773%next\;
        \$18493%now\ <= \$18493%next\;
        \$18579%now\ <= \$18579%next\;
        \$v5444%now\ <= \$v5444%next\;
        \$19524%now\ <= \$19524%next\;
        \$19247%now\ <= \$19247%next\;
        \$19122_modulo6684356_id%now\ <= \$19122_modulo6684356_id%next\;
        \$v5585%now\ <= \$v5585%next\;
        \$19494_loop666_result%now\ <= \$19494_loop666_result%next\;
        \$19284%now\ <= \$19284%next\;
        \$19373_compbranch6504392_id%now\ <= \$19373_compbranch6504392_id%next\;
        \$19287_v%now\ <= \$19287_v%next\;
        \$19808_forever6704342_id%now\ <= \$19808_forever6704342_id%next\;
        \$v5459%now\ <= \$v5459%next\;
        \$19767%now\ <= \$19767%next\;
        \$v5181%now\ <= \$v5181%next\;
        \$19494_loop666_id%now\ <= \$19494_loop666_id%next\;
        \$19529_forever6704351_id%now\ <= \$19529_forever6704351_id%next\;
        \$v5782%now\ <= \$v5782%next\;
        \$19053_binop_int6434369_id%now\ <= \$19053_binop_int6434369_id%next\;
        \$v4478%now\ <= \$v4478%next\;
        \$v5495%now\ <= \$v5495%next\;
        \$v4505%now\ <= \$v4505%next\;
        \$18621%now\ <= \$18621%next\;
        \$19598%now\ <= \$19598%next\;
        \$v4774%now\ <= \$v4774%next\;
        \$18523_aux664_result%now\ <= \$18523_aux664_result%next\;
        \$v5919%now\ <= \$v5919%next\;
        \$19298_v%now\ <= \$19298_v%next\;
        \$18872_v%now\ <= \$18872_v%next\;
        \$18817_v%now\ <= \$18817_v%next\;
        \$19762%now\ <= \$19762%next\;
        \$19002_modulo6684356_id%now\ <= \$19002_modulo6684356_id%next\;
        \$v5695%now\ <= \$v5695%next\;
        \$v5770%now\ <= \$v5770%next\;
        \$19024_modulo6684349_arg%now\ <= \$19024_modulo6684349_arg%next\;
        \$18936_modulo6684349_result%now\ <= \$18936_modulo6684349_result%next\;
        \$19428%now\ <= \$19428%next\;
        \$18890_v%now\ <= \$18890_v%next\;
        \$v5561%now\ <= \$v5561%next\;
        \$18535%now\ <= \$18535%next\;
        \$19151_modulo6684349_arg%now\ <= \$19151_modulo6684349_arg%next\;
        \result4399%now\ <= \result4399%next\;
        \$19278%now\ <= \$19278%next\;
        \rdy4435%now\ <= \rdy4435%next\;
        \$19000_res%now\ <= \$19000_res%next\;
        \$18609%now\ <= \$18609%next\;
        \$18720%now\ <= \$18720%next\;
        \$19552%now\ <= \$19552%next\;
        \$18757%now\ <= \$18757%next\;
        \$v4459%now\ <= \$v4459%next\;
        \$19305%now\ <= \$19305%next\;
        \$18874%now\ <= \$18874%next\;
        \$18800%now\ <= \$18800%next\;
        \$19607%now\ <= \$19607%next\;
        \$v4557%now\ <= \$v4557%next\;
        \$19757%now\ <= \$19757%next\;
        \$v4536%now\ <= \$v4536%next\;
        \$19933_w%now\ <= \$19933_w%next\;
        \$v4487%now\ <= \$v4487%next\;
        \$19258%now\ <= \$19258%next\;
        \$v4720%now\ <= \$v4720%next\;
        \$19151_modulo6684349_id%now\ <= \$19151_modulo6684349_id%next\;
        \$19744_w%now\ <= \$19744_w%next\;
        \result4572%now\ <= \result4572%next\;
        \$19103_r%now\ <= \$19103_r%next\;
        \$v5562%now\ <= \$v5562%next\;
        \$19178_res%now\ <= \$19178_res%next\;
        \$19160%now\ <= \$19160%next\;
        \$19663%now\ <= \$19663%next\;
        \$18871%now\ <= \$18871%next\;
        \$v5332%now\ <= \$v5332%next\;
        \$v5045%now\ <= \$v5045%next\;
        \$19193_v%now\ <= \$19193_v%next\;
        \$v4670%now\ <= \$v4670%next\;
        \$v5880%now\ <= \$v5880%next\;
        \$v5030%now\ <= \$v5030%next\;
        \$18883_v%now\ <= \$18883_v%next\;
        \$v4333%now\ <= \$v4333%next\;
        \$v5572%now\ <= \$v5572%next\;
        \$18983_modulo6684356_result%now\ <= \$18983_modulo6684356_result%next\;
        \$19493%now\ <= \$19493%next\;
        \$19095_res%now\ <= \$19095_res%next\;
        \$v5756%now\ <= \$v5756%next\;
        \$18983_modulo6684356_arg%now\ <= \$18983_modulo6684356_arg%next\;
        \$v5114%now\ <= \$v5114%next\;
        \$v5192%now\ <= \$v5192%next\;
        \$19461%now\ <= \$19461%next\;
        \$19107_modulo6684349_result%now\ <= \$19107_modulo6684349_result%next\;
        \$18839%now\ <= \$18839%next\;
        \$v5341%now\ <= \$v5341%next\;
        \$v5626%now\ <= \$v5626%next\;
        \$19050_modulo6684349_id%now\ <= \$19050_modulo6684349_id%next\;
        \$18787%now\ <= \$18787%next\;
        \$18716%now\ <= \$18716%next\;
        \$19121_r%now\ <= \$19121_r%next\;
        \$19206_binop_compare6454382_id%now\ <= \$19206_binop_compare6454382_id%next\;
        \$18885_v%now\ <= \$18885_v%next\;
        \$18658%now\ <= \$18658%next\;
        \$v5851%now\ <= \$v5851%next\;
        \$19069_modulo6684349_result%now\ <= \$19069_modulo6684349_result%next\;
        \$v5111%now\ <= \$v5111%next\;
        \$18678%now\ <= \$18678%next\;
        \$19822%now\ <= \$19822%next\;
        \$v5510%now\ <= \$v5510%next\;
        \$18753%now\ <= \$18753%next\;
        \$v5848%now\ <= \$v5848%next\;
        \$19113_forever6704372_arg%now\ <= \$19113_forever6704372_arg%next\;
        \$18840_v%now\ <= \$18840_v%next\;
        \$v5362%now\ <= \$v5362%next\;
        \$v4905%now\ <= \$v4905%next\;
        \$18596%now\ <= \$18596%next\;
        \$v4553%now\ <= \$v4553%next\;
        \$v5218%now\ <= \$v5218%next\;
        \$18440_make_block579_result%now\ <= \$18440_make_block579_result%next\;
        \$19401_compbranch6504396_id%now\ <= \$19401_compbranch6504396_id%next\;
        \$19380_compbranch6504393_result%now\ <= \$19380_compbranch6504393_result%next\;
        \$19047_modulo6684357_arg%now\ <= \$19047_modulo6684357_arg%next\;
        \$18861%now\ <= \$18861%next\;
        \$19931%now\ <= \$19931%next\;
        \$19340_argument2%now\ <= \$19340_argument2%next\;
        \$v4991%now\ <= \$v4991%next\;
        \$18983_modulo6684356_id%now\ <= \$18983_modulo6684356_id%next\;
        \$v5591%now\ <= \$v5591%next\;
        \$v5211%now\ <= \$v5211%next\;
        \$18920_binop_int6434362_id%now\ <= \$18920_binop_int6434362_id%next\;
        \$v5531%now\ <= \$v5531%next\;
        \$19002_modulo6684356_result%now\ <= \$19002_modulo6684356_result%next\;
        \$v4890%now\ <= \$v4890%next\;
        \$18589%now\ <= \$18589%next\;
        \$19144_modulo6684349_arg%now\ <= \$19144_modulo6684349_arg%next\;
        \$v4600%now\ <= \$v4600%next\;
        \$19476_v%now\ <= \$19476_v%next\;
        \$19587%now\ <= \$19587%next\;
        \$19919%now\ <= \$19919%next\;
        \$19574_w%now\ <= \$19574_w%next\;
        \$19237_v%now\ <= \$19237_v%next\;
        \$19037_v%now\ <= \$19037_v%next\;
        \$v5483%now\ <= \$v5483%next\;
        \$19634%now\ <= \$19634%next\;
        \$18585%now\ <= \$18585%next\;
        \$v4432%now\ <= \$v4432%next\;
        \$19365%now\ <= \$19365%next\;
        \$v5736%now\ <= \$v5736%next\;
        \$v4332%now\ <= \$v4332%next\;
        \$19857%now\ <= \$19857%next\;
        \$v5868%now\ <= \$v5868%next\;
        \$18803%now\ <= \$18803%next\;
        \$19346_sp%now\ <= \$19346_sp%next\;
        \$18691%now\ <= \$18691%next\;
        \$19846%now\ <= \$19846%next\;
        \$v5841%now\ <= \$v5841%next\;
        \$19695%now\ <= \$19695%next\;
        \$19494_loop666_arg%now\ <= \$19494_loop666_arg%next\;
        \$v5177%now\ <= \$v5177%next\;
        \$v4707%now\ <= \$v4707%next\;
        \$19122_modulo6684356_arg%now\ <= \$19122_modulo6684356_arg%next\;
        \$v4737%now\ <= \$v4737%next\;
        \$v5712%now\ <= \$v5712%next\;
        \$19370_compare6444359_arg%now\ <= \$19370_compare6444359_arg%next\;
        \$19622%now\ <= \$19622%next\;
        \$v4567%now\ <= \$v4567%next\;
        \$v5500%now\ <= \$v5500%next\;
        \$19899%now\ <= \$19899%next\;
        \$v5918%now\ <= \$v5918%next\;
        \$v5408%now\ <= \$v5408%next\;
        \$19039_r%now\ <= \$19039_r%next\;
        \$18814%now\ <= \$18814%next\;
        \$19738%now\ <= \$19738%next\;
        \$19670%now\ <= \$19670%next\;
        \$19457%now\ <= \$19457%next\;
        \$19377_compare6444359_id%now\ <= \$19377_compare6444359_id%next\;
        \$19556%now\ <= \$19556%next\;
        \$19711%now\ <= \$19711%next\;
        \$v5808%now\ <= \$v5808%next\;
        \$19377_compare6444359_arg%now\ <= \$19377_compare6444359_arg%next\;
        \$19405_compare6444359_result%now\ <= \$19405_compare6444359_result%next\;
        \$v5593%now\ <= \$v5593%next\;
        \$19903_next%now\ <= \$19903_next%next\;
        \$18818_v%now\ <= \$18818_v%next\;
        \$18633%now\ <= \$18633%next\;
        \$18466_loop666_arg%now\ <= \$18466_loop666_arg%next\;
        \$19459%now\ <= \$19459%next\;
        \$19705%now\ <= \$19705%next\;
        \$19629_hd%now\ <= \$19629_hd%next\;
        \$18836_v%now\ <= \$18836_v%next\;
        \$19384_compare6444359_arg%now\ <= \$19384_compare6444359_arg%next\;
        \$18736%now\ <= \$18736%next\;
        \$v5110%now\ <= \$v5110%next\;
        \$18671%now\ <= \$18671%next\;
        \$18686%now\ <= \$18686%next\;
        \$v4526%now\ <= \$v4526%next\;
        \$18990_modulo6684357_arg%now\ <= \$18990_modulo6684357_arg%next\;
        \$v5493%now\ <= \$v5493%next\;
        \$19632%now\ <= \$19632%next\;
        \$v5871%now\ <= \$v5871%next\;
        \$18823_v%now\ <= \$18823_v%next\;
        \$18593%now\ <= \$18593%next\;
        \$v5229%now\ <= \$v5229%next\;
        \$v5302%now\ <= \$v5302%next\;
        \$18652_w%now\ <= \$18652_w%next\;
        \$19506%now\ <= \$19506%next\;
        \$19337_compare6444359_result%now\ <= \$19337_compare6444359_result%next\;
        \$v4411%now\ <= \$v4411%next\;
        \$19680%now\ <= \$19680%next\;
        \rdy4964%now\ <= \rdy4964%next\;
        \$18690%now\ <= \$18690%next\;
        \$v4755%now\ <= \$v4755%next\;
        \$v5615%now\ <= \$v5615%next\;
        \$19195_compare6444358_id%now\ <= \$19195_compare6444358_id%next\;
        \$19912%now\ <= \$19912%next\;
        \$18469_make_block579_arg%now\ <= \$18469_make_block579_arg%next\;
        \$18743%now\ <= \$18743%next\;
        \$19791%now\ <= \$19791%next\;
        \$19604%now\ <= \$19604%next\;
        \$v5805%now\ <= \$v5805%next\;
        \$19510%now\ <= \$19510%next\;
        \$18728%now\ <= \$18728%next\;
        \$19869%now\ <= \$19869%next\;
        \$19900%now\ <= \$19900%next\;
        \$19898%now\ <= \$19898%next\;
        \$19111%now\ <= \$19111%next\;
        \$18586%now\ <= \$18586%next\;
        \$18986_modulo6684349_id%now\ <= \$18986_modulo6684349_id%next\;
        \$18468_wait662_id%now\ <= \$18468_wait662_id%next\;
        \$19244_v%now\ <= \$19244_v%next\;
        \$19612%now\ <= \$19612%next\;
        \$v4785%now\ <= \$v4785%next\;
        \$19847%now\ <= \$19847%next\;
        \$19398_compare6444359_arg%now\ <= \$19398_compare6444359_arg%next\;
        \$v4987%now\ <= \$v4987%next\;
        \$19830%now\ <= \$19830%next\;
        \$19034_binop_int6434368_id%now\ <= \$19034_binop_int6434368_id%next\;
        \$18856_loop_push6494360_result%now\ <= \$18856_loop_push6494360_result%next\;
        \$19687_w%now\ <= \$19687_w%next\;
        \$19745_hd%now\ <= \$19745_hd%next\;
        \$18894_v%now\ <= \$18894_v%next\;
        \$v5887%now\ <= \$v5887%next\;
        \$18672%now\ <= \$18672%next\;
        \$18617%now\ <= \$18617%next\;
        \$19938%now\ <= \$19938%next\;
        \$18892_v%now\ <= \$18892_v%next\;
        \$19437%now\ <= \$19437%next\;
        \$18636%now\ <= \$18636%next\;
        \$18611%now\ <= \$18611%next\;
        \$19225%now\ <= \$19225%next\;
        \$19420_w06554397_arg%now\ <= \$19420_w06554397_arg%next\;
        \$18713%now\ <= \$18713%next\;
        \$18616%now\ <= \$18616%next\;
        \$18771%now\ <= \$18771%next\;
        \$v4635%now\ <= \$v4635%next\;
        \$v5792%now\ <= \$v5792%next\;
        \$18868_v%now\ <= \$18868_v%next\;
        \$v5106%now\ <= \$v5106%next\;
        \$18693%now\ <= \$18693%next\;
        \$18597%now\ <= \$18597%next\;
        \$18437_loop666_result%now\ <= \$18437_loop666_result%next\;
        \$19426%now\ <= \$19426%next\;
        \$19763%now\ <= \$19763%next\;
        \$v5575%now\ <= \$v5575%next\;
        \$v4747%now\ <= \$v4747%next\;
        \$v5381%now\ <= \$v5381%next\;
        \$19151_modulo6684349_result%now\ <= \$19151_modulo6684349_result%next\;
        \$v5474%now\ <= \$v5474%next\;
        \$18850%now\ <= \$18850%next\;
        \$18445_x%now\ <= \$18445_x%next\;
        \$18798_w652_arg%now\ <= \$18798_w652_arg%next\;
        \$18878%now\ <= \$18878%next\;
        \$v5820%now\ <= \$v5820%next\;
        \$v5022%now\ <= \$v5022%next\;
        \$v4968%now\ <= \$v4968%next\;
        \$v4686%now\ <= \$v4686%next\;
        \$19472%now\ <= \$19472%next\;
        \$v5718%now\ <= \$v5718%next\;
        \$19404_b%now\ <= \$19404_b%next\;
        \$v4446%now\ <= \$v4446%next\;
        \$19624%now\ <= \$19624%next\;
        \$18587%now\ <= \$18587%next\;
        \$v5906%now\ <= \$v5906%next\;
        \$18970_r%now\ <= \$18970_r%next\;
        \$19545%now\ <= \$19545%next\;
        \$18534_next%now\ <= \$18534_next%next\;
        \$19219%now\ <= \$19219%next\;
        \$18792_wait662_id%now\ <= \$18792_wait662_id%next\;
        \$19265_ofs%now\ <= \$19265_ofs%next\;
        \$19618%now\ <= \$19618%next\;
        \$19411%now\ <= \$19411%next\;
        \$19468_sp%now\ <= \$19468_sp%next\;
        \$18547%now\ <= \$18547%next\;
        \$19116_binop_int6434373_id%now\ <= \$19116_binop_int6434373_id%next\;
        \$19065_r%now\ <= \$19065_r%next\;
        \$19645%now\ <= \$19645%next\;
        \$19129_modulo6684357_result%now\ <= \$19129_modulo6684357_result%next\;
        \$v5155%now\ <= \$v5155%next\;
        \$v5219%now\ <= \$v5219%next\;
        \$19756%now\ <= \$19756%next\;
        \$18490%now\ <= \$18490%next\;
        \$18523_aux664_arg%now\ <= \$18523_aux664_arg%next\;
        \$v5375%now\ <= \$v5375%next\;
        \$19215_argument1%now\ <= \$19215_argument1%next\;
        \$18860%now\ <= \$18860%next\;
        \$v5898%now\ <= \$v5898%next\;
        \$v4643%now\ <= \$v4643%next\;
        \$19174_binop_compare6454378_arg%now\ <= \$19174_binop_compare6454378_arg%next\;
        \$v5581%now\ <= \$v5581%next\;
        \$v4999%now\ <= \$v4999%next\;
        \$18466_loop666_result%now\ <= \$18466_loop666_result%next\;
        \$18469_make_block579_result%now\ <= \$18469_make_block579_result%next\;
        \$18625_copy_root_in_ram6634345_result%now\ <= \$18625_copy_root_in_ram6634345_result%next\;
        \$19640%now\ <= \$19640%next\;
        \$v4657%now\ <= \$v4657%next\;
        \$v5501%now\ <= \$v5501%next\;
        \$19323%now\ <= \$19323%next\;
        \$v5631%now\ <= \$v5631%next\;
        \$19270%now\ <= \$19270%next\;
        \$19473%now\ <= \$19473%next\;
        \$19318%now\ <= \$19318%next\;
        \$19132_modulo6684349_result%now\ <= \$19132_modulo6684349_result%next\;
        \$18548%now\ <= \$18548%next\;
        \$18967_modulo6684349_id%now\ <= \$18967_modulo6684349_id%next\;
        \$18772%now\ <= \$18772%next\;
        \$18628%now\ <= \$18628%next\;
        \$19562%now\ <= \$19562%next\;
        \$18538%now\ <= \$18538%next\;
        \$18819_v%now\ <= \$18819_v%next\;
        \$19198_binop_compare6454381_arg%now\ <= \$19198_binop_compare6454381_arg%next\;
        \$19465_sp%now\ <= \$19465_sp%next\;
        \$18526_aux664_result%now\ <= \$18526_aux664_result%next\;
        \$19911%now\ <= \$19911%next\;
        \$v4914%now\ <= \$v4914%next\;
        \$19446_sp%now\ <= \$19446_sp%next\;
        \$18932_r%now\ <= \$18932_r%next\;
        \$v4463%now\ <= \$v4463%next\;
        \$19946%now\ <= \$19946%next\;
        \$19943%now\ <= \$19943%next\;
        \$v5372%now\ <= \$v5372%next\;
        \$19577%now\ <= \$19577%next\;
        \$18641%now\ <= \$18641%next\;
        \$18773%now\ <= \$18773%next\;
        \$v5740%now\ <= \$v5740%next\;
        \$18524_loop666_id%now\ <= \$18524_loop666_id%next\;
        \$18964_modulo6684356_result%now\ <= \$18964_modulo6684356_result%next\;
        \$v4427%now\ <= \$v4427%next\;
        \$19655%now\ <= \$19655%next\;
        \$19028_modulo6684357_arg%now\ <= \$19028_modulo6684357_arg%next\;
        \$v4788%now\ <= \$v4788%next\;
        \$19520%now\ <= \$19520%next\;
        \$v4875%now\ <= \$v4875%next\;
        \$19306_v%now\ <= \$19306_v%next\;
        \$v5567%now\ <= \$v5567%next\;
        \$v5521%now\ <= \$v5521%next\;
        \$v4644%now\ <= \$v4644%next\;
        \$19343_sp%now\ <= \$19343_sp%next\;
        \$18722%now\ <= \$18722%next\;
        \$19935%now\ <= \$19935%next\;
        \$19056_v%now\ <= \$19056_v%next\;
        \$18513%now\ <= \$18513%next\;
        \$18989_r%now\ <= \$18989_r%next\;
        \$18879_v%now\ <= \$18879_v%next\;
        \$v4956%now\ <= \$v4956%next\;
        \$19730%now\ <= \$19730%next\;
        \$18665%now\ <= \$18665%next\;
        \$v4452%now\ <= \$v4452%next\;
        \$v5783%now\ <= \$v5783%next\;
        \$18710%now\ <= \$18710%next\;
        \$v5676%now\ <= \$v5676%next\;
        \$19009_modulo6684357_id%now\ <= \$19009_modulo6684357_id%next\;
        \$19712%now\ <= \$19712%next\;
        \$19841%now\ <= \$19841%next\;
        \$18556_forever6704344_arg%now\ <= \$18556_forever6704344_arg%next\;
        \$19780_loop665_result%now\ <= \$19780_loop665_result%next\;
        \$19236_v%now\ <= \$19236_v%next\;
        \$19330_compare6444359_result%now\ <= \$19330_compare6444359_result%next\;
        \$v5600%now\ <= \$v5600%next\;
        \$19330_compare6444359_arg%now\ <= \$19330_compare6444359_arg%next\;
        \$18592%now\ <= \$18592%next\;
        \$19289%now\ <= \$19289%next\;
        \$19589_copy_root_in_ram6634353_arg%now\ <= \$19589_copy_root_in_ram6634353_arg%next\;
        \$v4778%now\ <= \$v4778%next\;
        \$19356%now\ <= \$19356%next\;
        \$19050_modulo6684349_arg%now\ <= \$19050_modulo6684349_arg%next\;
        \$v5241%now\ <= \$v5241%next\;
        \$18594%now\ <= \$18594%next\;
        \$v5680%now\ <= \$v5680%next\;
        \$18866_v%now\ <= \$18866_v%next\;
        \$v5877%now\ <= \$v5877%next\;
        \$19424%now\ <= \$19424%next\;
        \$v5587%now\ <= \$v5587%next\;
        \$19369_b%now\ <= \$19369_b%next\;
        \$18481%now\ <= \$18481%next\;
        \$19050_modulo6684349_result%now\ <= \$19050_modulo6684349_result%next\;
        \$19691%now\ <= \$19691%next\;
        \$18471%now\ <= \$18471%next\;
        \$19058_r%now\ <= \$19058_r%next\;
        \$19560_hd%now\ <= \$19560_hd%next\;
        \$19405_compare6444359_id%now\ <= \$19405_compare6444359_id%next\;
        \$v5901%now\ <= \$v5901%next\;
        \$v5435%now\ <= \$v5435%next\;
        \$19353%now\ <= \$19353%next\;
        \$19059_modulo6684356_result%now\ <= \$19059_modulo6684356_result%next\;
        \$18910_modulo6684349_arg%now\ <= \$18910_modulo6684349_arg%next\;
        \$v5706%now\ <= \$v5706%next\;
        \$18486%now\ <= \$18486%next\;
        \$18501%now\ <= \$18501%next\;
        \$18532%now\ <= \$18532%next\;
        \$v4764%now\ <= \$v4764%next\;
        \$19216_v%now\ <= \$19216_v%next\;
        \$19613_w%now\ <= \$19613_w%next\;
        \$18528%now\ <= \$18528%next\;
        \$19283%now\ <= \$19283%next\;
        \$v5338%now\ <= \$v5338%next\;
        \$19091_binop_int6434371_result%now\ <= \$19091_binop_int6434371_result%next\;
        \$v4962%now\ <= \$v4962%next\;
        \$19654%now\ <= \$19654%next\;
        \$v5842%now\ <= \$v5842%next\;
        \$v5527%now\ <= \$v5527%next\;
        \$18920_binop_int6434362_result%now\ <= \$18920_binop_int6434362_result%next\;
        \$19195_compare6444358_arg%now\ <= \$19195_compare6444358_arg%next\;
        \$v5910%now\ <= \$v5910%next\;
        \$18705_next%now\ <= \$18705_next%next\;
        \$19511%now\ <= \$19511%next\;
        \$v5902%now\ <= \$v5902%next\;
        \$19410%now\ <= \$19410%next\;
        \$18468_wait662_arg%now\ <= \$18468_wait662_arg%next\;
        \$v5504%now\ <= \$v5504%next\;
        \$v4522%now\ <= \$v4522%next\;
        \$18797_branch_if648_arg%now\ <= \$18797_branch_if648_arg%next\;
        \$19696%now\ <= \$19696%next\;
        \$18955_modulo6684349_arg%now\ <= \$18955_modulo6684349_arg%next\;
        \$19652%now\ <= \$19652%next\;
        \$19606%now\ <= \$19606%next\;
        \$19195_compare6444358_result%now\ <= \$19195_compare6444358_result%next\;
        \$v5006%now\ <= \$v5006%next\;
        \$18804%now\ <= \$18804%next\;
        \$18910_modulo6684349_result%now\ <= \$18910_modulo6684349_result%next\;
        \$19502%now\ <= \$19502%next\;
        \$v5583%now\ <= \$v5583%next\;
        \$18853_hd%now\ <= \$18853_hd%next\;
        \$v5746%now\ <= \$v5746%next\;
        \$v5048%now\ <= \$v5048%next\;
        \$19831%now\ <= \$19831%next\;
        \$19481%now\ <= \$19481%next\;
        \$18774%now\ <= \$18774%next\;
        \$19708%now\ <= \$19708%next\;
        \$18632%now\ <= \$18632%next\;
        \$18625_copy_root_in_ram6634345_arg%now\ <= \$18625_copy_root_in_ram6634345_arg%next\;
        \$v5834%now\ <= \$v5834%next\;
        \$19568%now\ <= \$19568%next\;
        \$v4723%now\ <= \$v4723%next\;
        \$18519%now\ <= \$18519%next\;
        \$v4580%now\ <= \$v4580%next\;
        \$19547_copy_root_in_ram6634352_arg%now\ <= \$19547_copy_root_in_ram6634352_arg%next\;
        \$19477_v%now\ <= \$19477_v%next\;
        \$18704%now\ <= \$18704%next\;
        \$18503%now\ <= \$18503%next\;
        \$18790_loop666_arg%now\ <= \$18790_loop666_arg%next\;
        \$v5854%now\ <= \$v5854%next\;
        \$19690%now\ <= \$19690%next\;
        \$v5786%now\ <= \$v5786%next\;
        \$19498_loop665_id%now\ <= \$19498_loop665_id%next\;
        \$v5864%now\ <= \$v5864%next\;
        \$v5886%now\ <= \$v5886%next\;
        \$18923_v%now\ <= \$18923_v%next\;
        \$v5914%now\ <= \$v5914%next\;
        \$v5798%now\ <= \$v5798%next\;
        \$v5016%now\ <= \$v5016%next\;
        \$19499_aux664_result%now\ <= \$19499_aux664_result%next\;
        \$v5554%now\ <= \$v5554%next\;
        \$18675%now\ <= \$18675%next\;
        \$18463%now\ <= \$18463%next\;
        \$19469%now\ <= \$19469%next\;
        \$18700%now\ <= \$18700%next\;
        \$18744_w%now\ <= \$18744_w%next\;
        \$v5087%now\ <= \$v5087%next\;
        \$18530%now\ <= \$18530%next\;
        \$v5423%now\ <= \$v5423%next\;
        \$v5215%now\ <= \$v5215%next\;
        \$18929_modulo6684349_result%now\ <= \$18929_modulo6684349_result%next\;
        \$19733%now\ <= \$19733%next\;
        \$18653_hd%now\ <= \$18653_hd%next\;
        \$19429%now\ <= \$19429%next\;
        \$18833%now\ <= \$18833%next\;
        \$v5165%now\ <= \$v5165%next\;
        \$18454%now\ <= \$18454%next\;
        \$18847%now\ <= \$18847%next\;
        \$v5553%now\ <= \$v5553%next\;
        \$v5075%now\ <= \$v5075%next\;
        \$18692%now\ <= \$18692%next\;
        \$18719%now\ <= \$18719%next\;
        \$19940%now\ <= \$19940%next\;
        \$18712_hd%now\ <= \$18712_hd%next\;
        \$v5417%now\ <= \$v5417%next\;
        \$19125_modulo6684349_arg%now\ <= \$19125_modulo6684349_arg%next\;
        \$18634%now\ <= \$18634%next\;
        \$19484%now\ <= \$19484%next\;
        \$18929_modulo6684349_id%now\ <= \$18929_modulo6684349_id%next\;
        \$19198_binop_compare6454381_id%now\ <= \$19198_binop_compare6454381_id%next\;
        \$19416_w36574398_id%now\ <= \$19416_w36574398_id%next\;
        \$18798_w652_id%now\ <= \$18798_w652_id%next\;
        \$v5056%now\ <= \$v5056%next\;
        \$v4439%now\ <= \$v4439%next\;
        \$v5503%now\ <= \$v5503%next\;
        \$19608%now\ <= \$19608%next\;
        \$v5779%now\ <= \$v5779%next\;
        \$19277%now\ <= \$19277%next\;
        \$19223%now\ <= \$19223%next\;
        \$18499%now\ <= \$18499%next\;
        \$18796_make_block_n646_result%now\ <= \$18796_make_block_n646_result%next\;
        \$19085_modulo6684357_id%now\ <= \$19085_modulo6684357_id%next\;
        \$v5399%now\ <= \$v5399%next\;
        \$v4808%now\ <= \$v4808%next\;
        \$18811%now\ <= \$18811%next\;
        \$19808_forever6704342_arg%now\ <= \$19808_forever6704342_arg%next\;
        \$v4508%now\ <= \$v4508%next\;
        \$v5207%now\ <= \$v5207%next\;
        \$v5093%now\ <= \$v5093%next\;
        \$19034_binop_int6434368_result%now\ <= \$19034_binop_int6434368_result%next\;
        \$19627%now\ <= \$19627%next\;
        \$19881_hd%now\ <= \$19881_hd%next\;
        \$19291_v%now\ <= \$19291_v%next\;
        \$18901_binop_int6434361_id%now\ <= \$18901_binop_int6434361_id%next\;
        \$19387_compbranch6504394_result%now\ <= \$19387_compbranch6504394_result%next\;
        \$19644_hd%now\ <= \$19644_hd%next\;
        \$19347_fill6534389_id%now\ <= \$19347_fill6534389_id%next\;
        \$v5917%now\ <= \$v5917%next\;
        \$19792%now\ <= \$19792%next\;
        \$19541%now\ <= \$19541%next\;
        \$v5480%now\ <= \$v5480%next\;
        \$19415_sp%now\ <= \$19415_sp%next\;
        \$19262_forever6704385_arg%now\ <= \$19262_forever6704385_arg%next\;
        \$18477%now\ <= \$18477%next\;
        \$19635%now\ <= \$19635%next\;
        \$v4933%now\ <= \$v4933%next\;
        \$19633%now\ <= \$19633%next\;
        \$v4566%now\ <= \$v4566%next\;
        \$18917_modulo6684349_id%now\ <= \$18917_modulo6684349_id%next\;
        \$18451%now\ <= \$18451%next\;
        \$19802%now\ <= \$19802%next\;
        \$19221%now\ <= \$19221%next\;
        \$19224%now\ <= \$19224%next\;
        \$v5240%now\ <= \$v5240%next\;
        \$19516%now\ <= \$19516%next\;
        \$18656%now\ <= \$18656%next\;
        \$19693%now\ <= \$19693%next\;
        \$18496%now\ <= \$18496%next\;
        \$18588%now\ <= \$18588%next\;
        \$18887_v%now\ <= \$18887_v%next\;
        \$19360_sp%now\ <= \$19360_sp%next\;
        \$19171_compare6444358_result%now\ <= \$19171_compare6444358_result%next\;
        \$19688_hd%now\ <= \$19688_hd%next\;
        \$18491%now\ <= \$18491%next\;
        \$18541%now\ <= \$18541%next\;
        \$19380_compbranch6504393_arg%now\ <= \$19380_compbranch6504393_arg%next\;
        \$19782%now\ <= \$19782%next\;
        \$v5517%now\ <= \$v5517%next\;
        \$19141_modulo6684356_id%now\ <= \$19141_modulo6684356_id%next\;
        \$19107_modulo6684349_id%now\ <= \$19107_modulo6684349_id%next\;
        \$v4971%now\ <= \$v4971%next\;
        \$v4848%now\ <= \$v4848%next\;
        \$19166_binop_compare6454377_result%now\ <= \$19166_binop_compare6454377_result%next\;
        \$19593%now\ <= \$19593%next\;
        \$18568%now\ <= \$18568%next\;
        \$v4625%now\ <= \$v4625%next\;
        \$18452%now\ <= \$18452%next\;
        \$19742%now\ <= \$19742%next\;
        \$v4869%now\ <= \$v4869%next\;
        \$v5590%now\ <= \$v5590%next\;
        \$18468_wait662_result%now\ <= \$18468_wait662_result%next\;
        \$19575_hd%now\ <= \$19575_hd%next\;
        \$19229_v%now\ <= \$19229_v%next\;
        \$18981_res%now\ <= \$18981_res%next\;
        \$v4622%now\ <= \$v4622%next\;
        \$18942_v%now\ <= \$18942_v%next\;
        \$18543%now\ <= \$18543%next\;
        \$19513%now\ <= \$19513%next\;
        \$19555%now\ <= \$19555%next\;
        \$19692%now\ <= \$19692%next\;
        \$19370_compare6444359_result%now\ <= \$19370_compare6444359_result%next\;
        \$v4896%now\ <= \$v4896%next\;
        \$v5661%now\ <= \$v5661%next\;
        \$v5520%now\ <= \$v5520%next\;
        \$18917_modulo6684349_result%now\ <= \$18917_modulo6684349_result%next\;
        \$19116_binop_int6434373_result%now\ <= \$19116_binop_int6434373_result%next\;
        \$v4404%now\ <= \$v4404%next\;
        \$19862%now\ <= \$19862%next\;
        \$18449%now\ <= \$18449%next\;
        \$19573%now\ <= \$19573%next\;
        \$19729%now\ <= \$19729%next\;
        \$18952_modulo6684357_id%now\ <= \$18952_modulo6684357_id%next\;
        \$19252_forever6704384_arg%now\ <= \$19252_forever6704384_arg%next\;
        \$19805%now\ <= \$19805%next\;
        \$18943_res%now\ <= \$18943_res%next\;
        \$v4564%now\ <= \$v4564%next\;
        \$18926_modulo6684356_arg%now\ <= \$18926_modulo6684356_arg%next\;
        \$v5438%now\ <= \$v5438%next\;
        \$19567%now\ <= \$19567%next\;
        \$18761%now\ <= \$18761%next\;
        \$v5350%now\ <= \$v5350%next\;
        \$v5230%now\ <= \$v5230%next\;
        \$v4731%now\ <= \$v4731%next\;
        \$19838_copy_root_in_ram6634340_arg%now\ <= \$19838_copy_root_in_ram6634340_arg%next\;
        \$v5667%now\ <= \$v5667%next\;
        \$v5535%now\ <= \$v5535%next\;
        \$19008_r%now\ <= \$19008_r%next\;
        \$v5547%now\ <= \$v5547%next\;
        \$19669%now\ <= \$19669%next\;
        \$18862%now\ <= \$18862%next\;
        \$19699%now\ <= \$19699%next\;
        \$19630%now\ <= \$19630%next\;
        \$ram_lock%now\ <= \$ram_lock%next\;
        \$global_end_lock%now\ <= \$global_end_lock%next\;
        \$code_lock%now\ <= \$code_lock%next\;
        \state_var5924%now\ <= \state_var5924%next\;
        \state_var5923%now\ <= \state_var5923%next\;
        \state_var5922%now\ <= \state_var5922%next\;
        \state_var5921%now\ <= \state_var5921%next\;
        \state_var5920%now\ <= \state_var5920%next\;
        \state%now\ <= \state%next\;
      end if;
    end process;
      
      process(argument,\state%now\, clk,\state_var5924%now\,\state_var5923%now\,\state_var5922%now\,\state_var5921%now\,\state_var5920%now\, \$ram_value\, \$global_end_value\, \$code_value\, \$18606%now\, \$19190_binop_compare6454380_arg%now\, \$v4743%now\, \$19072_binop_int6434370_arg%now\, \$18910_modulo6684349_id%now\, \$19299%now\, \$19069_modulo6684349_id%now\, \$v5526%now\, \$v4663%now\, \$v5913%now\, \$18602%now\, \$v5541%now\, \$18809%now\, \$18751%now\, \$19272%now\, \$v5486%now\, \$v5513%now\, \$18729%now\, \$v5507%now\, \$18801%now\, \$19779_loop666_id%now\, \$18775%now\, \$19874%now\, \$v5715%now\, \$18974_modulo6684349_id%now\, \$19828%now\, \$v4961%now\, \$v4499%now\, \$19326_compbranch6504387_result%now\, \$v5326%now\, \$v5484%now\, \$18504%now\, \$v5643%now\, \$18945_modulo6684356_result%now\, \$18933_modulo6684357_id%now\, \$19250%now\, \$18624%now\, \$v4650%now\, \$19553%now\, \$18637_w%now\, \$19380_compbranch6504393_id%now\, \$v5619%now\, \$18835%now\, \$19579%now\, \$19758%now\, \$19085_modulo6684357_result%now\, \$18776%now\, \$18875_v%now\, \$19132_modulo6684349_id%now\, \$18619%now\, \$19163_forever6704376_arg%now\, \$v4604%now\, \$v5699%now\, \$19292%now\, \$v5634%now\, \$19416_w36574398_result%now\, \$18993_modulo6684349_result%now\, \$18581%now\, \$19866_hd%now\, \$v5287%now\, \$v4467%now\, \$18900%now\, \$v4470%now\, \$v4325%now\, \$18696%now\, \$19245%now\, \$19024_modulo6684349_result%now\, \$18945_modulo6684356_arg%now\, \$19689%now\, \$v4577%now\, \$19140_r%now\, \$18802%now\, \$v5076%now\, \$19001_r%now\, \$v5532%now\, \$19501%now\, \$18769_hd%now\, \$v5152%now\, \$v4703%now\, \$19122_modulo6684356_result%now\, \$19499_aux664_id%now\, \$18483%now\, \$19290%now\, \$19273%now\, \$19104_modulo6684357_id%now\, \$v4710%now\, \$v4814%now\, \$19170_res%now\, \$18924_res%now\, \$19863%now\, \$18821_v%now\, \$19827%now\, \$19432%now\, \$19448_v%now\, \$18630%now\, \$19094_v%now\, \$v4535%now\, \$v5551%now\, \$19028_modulo6684357_result%now\, \$18939_binop_int6434363_result%now\, \$v5824%now\, \$18788%now\, \$v5226%now\, \$18582%now\, \$19081_modulo6684349_arg%now\, \$v5013%now\, \$18881_hd%now\, \$19525%now\, \$18509%now\, \$18793_make_block579_result%now\, \$18974_modulo6684349_arg%now\, \$19235_v%now\, \$v4515%now\, \$v5323%now\, \$18655%now\, \$19906%now\, \$v5592%now\, \$19194_res%now\, \$18990_modulo6684357_result%now\, \$19947%now\, \$19672%now\, \$v5692%now\, \$18474%now\, \$19641%now\, \$18855_next_env%now\, \$v5158%now\, \$19040_modulo6684356_id%now\, \$v5369%now\, \$v5733%now\, \$19661%now\, \$v5414%now\, \$v4443%now\, \$18876%now\, \$19653%now\, \$19508%now\, \$19358%now\, \$v5151%now\, \$v5594%now\, \$19043_modulo6684349_result%now\, \$18859%now\, \$v4830%now\, \$v5117%now\, \$19445%now\, \$18867%now\, \$v5752%now\, \$18865%now\, \$19890%now\, \$v4511%now\, \$18455%now\, \$18512%now\, \$v4590%now\, \$19427%now\, \$19934_hd%now\, \$18846%now\, \$18524_loop666_result%now\, \$v4472%now\, \$19723%now\, \$18778%now\, \$18694%now\, \$v5759%now\, \$19066_modulo6684357_result%now\, \$19850_w%now\, \$19419%now\, \$18961_v%now\, \$19201_v%now\, \$v5703%now\, \$19274_v%now\, \$19394_compbranch6504395_arg%now\, \$v5320%now\, \$19166_binop_compare6454377_arg%now\, \$v5212%now\, \$19704%now\, \$19930%now\, \$v5721%now\, \$19458%now\, \$19185_v%now\, \$v5586%now\, \$18738_next%now\, \$19364_v%now\, \$v5234%now\, \$v5760%now\, \$18974_modulo6684349_result%now\, \$19797_next%now\, \$18745_hd%now\, \$18797_branch_if648_result%now\, \$19589_copy_root_in_ram6634353_id%now\, \$v5766%now\, \$19478_v%now\, \$19752%now\, \$v4616%now\, \$19894%now\, \$19819%now\, \$19489%now\, \$v5776%now\, \$v5019%now\, \$18807%now\, \$19504%now\, \$18650%now\, \$18837%now\, \$18569%now\, \$19129_modulo6684357_id%now\, \$18805%now\, \$v5869%now\, \$19112%now\, \$19135_binop_int6434374_arg%now\, \$19002_modulo6684356_arg%now\, \$v5515%now\, \$19319%now\, \$v5646%now\, \$v4952%now\, \$v5610%now\, \$v5683%now\, \$18958_binop_int6434364_result%now\, \$19342%now\, \$19657%now\, \$19777%now\, \$19620%now\, \$18793_make_block579_id%now\, \$18521_loop666_arg%now\, \$19803%now\, \$19217%now\, \$v4949%now\, \$19486%now\, \$v5857%now\, \$18482%now\, \$v4692%now\, \$19309_v%now\, \$18529%now\, \$19916%now\, \$v5686%now\, \$v4854%now\, \$v4628%now\, \$18703%now\, \$v5506%now\, \$v4926%now\, \$19829%now\, \$v4523%now\, \$v4569%now\, \$v5749%now\, \$19209_v%now\, \$19482%now\, \$19611%now\, \$19811_copy_root_in_ram6634341_id%now\, \$19784%now\, \$18502%now\, \$v4770%now\, \$18667_w%now\, \$19434%now\, \$19333_compbranch6504388_arg%now\, \$19732%now\, \$19609%now\, \$19714_next%now\, \$18815%now\, \$v5210%now\, \$18565%now\, \$v4491%now\, \$19076_res%now\, \$v4727%now\, \$19015_binop_int6434367_id%now\, \$18986_modulo6684349_arg%now\, \$v4734%now\, \$19656%now\, \$19496_aux664_arg%now\, \$18480%now\, \$v5537%now\, \$18458%now\, \$18993_modulo6684349_arg%now\, \$v5655%now\, \$19294%now\, \$v5828%now\, \$19583%now\, \$v5838%now\, \$19163_forever6704376_id%now\, \$18723%now\, \$v4481%now\, \$v5640%now\, \$19314%now\, \$18762%now\, \$19034_binop_int6434368_arg%now\, \$v4728%now\, \$v4596%now\, \$19062_modulo6684349_result%now\, \$18914_modulo6684357_arg%now\, \$18590%now\, \$19902%now\, \$18670%now\, \$v5604%now\, \$19248%now\, \$19088_modulo6684349_result%now\, \$19464%now\, \$19072_binop_int6434370_result%now\, \$v4761%now\, \$19816%now\, \$19081_modulo6684349_result%now\, \$v4845%now\, \$v4631%now\, \$19326_compbranch6504387_arg%now\, \$v5035%now\, \$18685%now\, \$v5603%now\, \$19628_w%now\, \$v5582%now\, \$18948_modulo6684349_arg%now\, \$v5060%now\, \$18668_hd%now\, \$v4552%now\, \$19187_compare6444358_result%now\, \$v5378%now\, \$19623%now\, \$v5052%now\, \$v4946%now\, \$18664%now\, \$18646%now\, \$18852%now\, \$18485%now\, \$19190_binop_compare6454380_result%now\, \$19043_modulo6684349_arg%now\, \$v4936%now\, \$v4417%now\, \$18447%now\, \$v4992%now\, \$v5702%now\, \$18967_modulo6684349_arg%now\, \$v5481%now\, \$18952_modulo6684357_result%now\, \$18662%now\, \$18600%now\, \$v5244%now\, \$19600%now\, \$19838_copy_root_in_ram6634340_result%now\, \$19885%now\, \$19685%now\, \$19187_compare6444358_id%now\, \$18926_modulo6684356_id%now\, \$19720_w%now\, \$v5530%now\, \$18644%now\, \$18466_loop666_id%now\, \$18638_hd%now\, \$v4674%now\, \$v5250%now\, \$18563%now\, \$19062_modulo6684349_id%now\, \$18645%now\, \$19897%now\, \$19139_res%now\, \$19347_fill6534389_arg%now\, \$19495_loop665_arg%now\, \$v4695%now\, \$18576%now\, \$18578%now\, \$18440_make_block579_arg%now\, \$19157_forever6704375_id%now\, \$19246_v%now\, \$19495_loop665_id%now\, \$19515_next%now\, \$v4563%now\, \$v4908%now\, \$18635%now\, \$19251%now\, \$19648%now\, \$18613_copy_root_in_ram6634346_id%now\, \$19780_loop665_arg%now\, \$18571_copy_root_in_ram6634345_arg%now\, \$v5120%now\, \$19854%now\, \$v4988%now\, \$v5607%now\, \$19848%now\, \$19232%now\, \$19814%now\, \$v4680%now\, \$18906_r%now\, \$v5127%now\, \$18620%now\, \$19887%now\, \$19296_v%now\, \$18709%now\, \$v4805%now\, \$v5514%now\, \$18913_r%now\, \$18457%now\, \$19269%now\, \$19569%now\, \$v5823%now\, \$v5164%now\, \$19721_hd%now\, \$v5831%now\, \$v4740%now\, \$v5308%now\, \$v4995%now\, \$v4601%now\, \$18484%now\, \$18733%now\, \$v4660%now\, \$19408_argument3%now\, \$18828_v%now\, \$19390_b%now\, \$19727%now\, \$18510%now\, \$19662%now\, \$v5577%now\, \$19015_binop_int6434367_arg%now\, \$19413%now\, \$v4584%now\, \$19845%now\, \$19337_compare6444359_id%now\, \$19698%now\, \$18566%now\, \$18767%now\, \$19359%now\, \$18977_binop_int6434365_arg%now\, \$v4878%now\, \$19267_hd%now\, \$19679%now\, \$v5195%now\, \$v4433%now\, \$18864%now\, \$18996_binop_int6434366_arg%now\, \$19599%now\, \$19526_forever6704355_arg%now\, \$19578%now\, \$18605%now\, \$19558%now\, \$19280%now\, \$v5278%now\, \$v5557%now\, \$19817%now\, \$19238_w6514383_arg%now\, \$v5284%now\, \$v5905%now\, \$19488%now\, \$19474%now\, \$v5564%now\, \$18591%now\, \$v4568%now\, \$v5883%now\, \$v5555%now\, \$19726%now\, \$v4842%now\, \$18834_v%now\, \$19401_compbranch6504396_result%now\, \$18699%now\, \$18680%now\, \$19751%now\, \$19157_forever6704375_arg%now\, \$18584_hd%now\, \$19867%now\, \$v5465%now\, \$18999_v%now\, \$18623%now\, \$19754%now\, \$19825%now\, \$19312_v%now\, \$18936_modulo6684349_arg%now\, \$18460%now\, \$19596%now\, \$18795_offsetclosure_n639_result%now\, \$19918%now\, \$v4328%now\, \$19373_compbranch6504392_result%now\, \$v5247%now\, \$v4543%now\, \$v5420%now\, \$19505%now\, \$18570%now\, \$v5263%now\, \$19391_compare6444359_id%now\, \$v5835%now\, \$18962_res%now\, \$18822_v%now\, \$v5614%now\, \$v5027%now\, \$18610%now\, \$v5069%now\, \$18684%now\, \$19535_copy_root_in_ram6634354_id%now\, \$v5860%now\, \$v4414%now\, \$v5237%now\, \$19066_modulo6684357_arg%now\, \$19852%now\, \$18577%now\, \$v5533%now\, \$18553_forever6704348_arg%now\, \$19387_compbranch6504394_id%now\, \$18643%now\, \$18754%now\, \$18933_modulo6684357_arg%now\, \$19397_b%now\, \$19279_v%now\, \$18933_modulo6684357_result%now\, \$v5485%now\, \$19550%now\, \$18816%now\, \$19495_loop665_result%now\, \$v5516%now\, \$v5180%now\, \$18952_modulo6684357_arg%now\, \$19855%now\, \$v5426%now\, \$19313%now\, \$v5542%now\, \$19565%now\, \$v4863%now\, \$18980_v%now\, \$18521_loop666_id%now\, \$v5870%now\, \$19800_next%now\, \$19746%now\, \$19851_hd%now\, \$18488%now\, \$18746%now\, \$v5203%now\, \$19222%now\, \$v5290%now\, \$18796_make_block_n646_id%now\, \$19096_r%now\, \$19450_v%now\, \$19651%now\, \$v5130%now\, \$v5595%now\, \$v4699%now\, \$18559_copy_root_in_ram6634347_result%now\, \$18831%now\, \$v5123%now\, \$18829%now\, \$19761%now\, \$19547_copy_root_in_ram6634352_result%now\, \$v5737%now\, \$19676%now\, \$18450%now\, \$18982_r%now\, \$19179_compare6444358_arg%now\, \$v4462%now\, \$18717%now\, \$v5148%now\, \$18571_copy_root_in_ram6634345_id%now\, \$v5170%now\, \$19438%now\, \$19647%now\, \$19483%now\, \$19361_fill6544390_arg%now\, \$19861%now\, \$19211_compare6444358_id%now\, \$19786%now\, \$18725%now\, \$18459%now\, \$19135_binop_int6434374_result%now\, \$v5546%now\, \$19724%now\, \$18711_w%now\, \$18948_modulo6684349_result%now\, \$v5144%now\, \$19908%now\, \$19858%now\, \$18779%now\, \$v5272%now\, \$18612%now\, \$19303%now\, \$19551%now\, \$v5269%now\, \$19186_res%now\, \$18689%now\, \$19631%now\, \$18791_loop665_arg%now\, \$18905_res%now\, \$19694%now\, \$18755%now\, \$v5795%now\, \$v5202%now\, \$v5565%now\, \$v4923%now\, \$19835%now\, \$19588%now\, \$v4943%now\, \$19078_modulo6684356_id%now\, \$v5317%now\, \result4434%now\, \$v5512%now\, \$18465%now\, \$v4484%now\, \$18830_v%now\, \$19779_loop666_arg%now\, \$19616%now\, \$v4792%now\, \$19088_modulo6684349_arg%now\, \$19666%now\, \$19179_compare6444358_id%now\, \$19681_next%now\, \$18742%now\, \$18795_offsetclosure_n639_arg%now\, \$19384_compare6444359_id%now\, \$18993_modulo6684349_id%now\, \$19610%now\, \$18856_loop_push6494360_arg%now\, \$19909_w%now\, \$19686%now\, \$v4975%now\, \$19019_res%now\, \$v5534%now\, \$18479%now\, \$18525_loop665_result%now\, \$v5893%now\, \$19671%now\, \$v4475%now\, \$18734%now\, \$19128_r%now\, \$19750%now\, \$19499_aux664_arg%now\, \$19826%now\, \$18799_w1656_result%now\, \$18798_w652_result%now\, \$18467_loop665_arg%now\, \$19021_modulo6684356_id%now\, \$19088_modulo6684349_id%now\, \$19162%now\, \$v4851%now\, \$19357_v%now\, \$19097_modulo6684356_result%now\, \$v5580%now\, \$19012_modulo6684349_id%now\, \$18765%now\, \$v4893%now\, \$v5329%now\, \$19936%now\, \$19020_r%now\, \$19238_w6514383_result%now\, \$v5601%now\, \$18996_binop_int6434366_id%now\, \$v5511%now\, \$v4570%now\, \$19675%now\, \$18601%now\, \$v4565%now\, \$18552%now\, \$19077_r%now\, \$v5545%now\, \$v5031%now\, \$v5456%now\, \$v5161%now\, \$19075_v%now\, \$18791_loop665_result%now\, \$18750%now\, \$18718%now\, \$19849%now\, \$19059_modulo6684356_arg%now\, \$v4724%now\, \$19423_v%now\, \$19352%now\, \$19601_copy_root_in_ram6634352_result%now\, \$18789%now\, \$18977_binop_int6434365_id%now\, \$v5789%now\, \$v5450%now\, \$18681%now\, \$19206_binop_compare6454382_arg%now\, \$v5010%now\, \$19523%now\, \$18964_modulo6684356_id%now\, \$19923%now\, \$19361_fill6544390_result%now\, \$19535_copy_root_in_ram6634354_arg%now\, \$19564%now\, \$18770%now\, \$19790%now\, \$19509%now\, \$18598_w%now\, \$18462%now\, \$19873%now\, \$v5496%now\, \$v5573%now\, \$19177_v%now\, \$19320_forever6704386_arg%now\, \$19069_modulo6684349_arg%now\, \$v5225%now\, \$v5611%now\, \$v5063%now\, \$v5393%now\, \$19778%now\, \$19821%now\, \$v5174%now\, \$18494%now\, \$19333_compbranch6504388_result%now\, \$19441_arg%now\, \$18920_binop_int6434362_arg%now\, \$v5080%now\, \$18790_loop666_id%now\, \$v5763%now\, \$v5618%now\, \$18613_copy_root_in_ram6634346_result%now\, \$19498_loop665_arg%now\, \$19467_sp%now\, \$v4799%now\, \$19187_compare6444358_arg%now\, \$v4860%now\, \$18849%now\, \$18749%now\, \$18907_modulo6684356_id%now\, \$19794%now\, \$18863%now\, \$19910_hd%now\, \$18958_binop_int6434364_id%now\, \$v5135%now\, \$v4495%now\, \$19320_forever6704386_id%now\, \$19300%now\, \$19116_binop_int6434373_arg%now\, \$v5147%now\, \$v4899%now\, \$19333_compbranch6504388_id%now\, \$19880_w%now\, \$v5730%now\, \$19366_compbranch6504391_arg%now\, \$v5007%now\, \$19377_compare6444359_result%now\, \$19203_compare6444358_result%now\, \$v5570%now\, \$19664%now\, \$19637%now\, \$18926_modulo6684356_result%now\, \$v4431%now\, \$18854_sp%now\, \$19710%now\, \$19771%now\, \$19057_res%now\, \$18907_modulo6684356_arg%now\, \$18537%now\, \$19785%now\, \$18792_wait662_result%now\, \$18826%now\, \$19307_v%now\, \$19354_v%now\, \$19463%now\, \$19734%now\, \rdy4929%now\, \$18799_w1656_id%now\, \$19589_copy_root_in_ram6634353_result%now\, \$18472%now\, \$v4666%now\, \$19129_modulo6684357_arg%now\, \$v4458%now\, \$18873_v%now\, \$19038_res%now\, \$19595%now\, \$19883%now\, \$18677%now\, \$19249%now\, \$v5266%now\, \$19546%now\, \$v4767%now\, \$v5189%now\, \$v4442%now\, \$19891%now\, \$v5649%now\, \$v5199%now\, \$19559_w%now\, \$19920%now\, \$v4549%now\, \$18990_modulo6684357_id%now\, \$19107_modulo6684349_arg%now\, \$18520%now\, \$19420_w06554397_result%now\, \$18884_v%now\, \$18925_r%now\, \$19179_compare6444358_result%now\, \$19078_modulo6684356_arg%now\, \$v5103%now\, \$19522%now\, \$19544%now\, \$19243%now\, \$19718%now\, \$19148_modulo6684357_arg%now\, \$19538%now\, \$19255%now\, \$v4571%now\, \$19275%now\, \$19281%now\, \$18599_hd%now\, \$19836%now\, \$v4872%now\, \$19043_modulo6684349_id%now\, \$19884%now\, \$19871%now\, \$18851%now\, \$19557%now\, \$19517%now\, \$19532_forever6704350_id%now\, \$18782%now\, \$18526_aux664_id%now\, \$v4696%now\, \$19238_w6514383_id%now\, \$19582%now\, \$v5344%now\, \$19570%now\, \$v4619%now\, \$19888%now\, \$18794_apply638_id%now\, \$19497_loop666_id%now\, \$v4651%now\, \$18521_loop666_result%now\, \$19901%now\, \$18442_cy%now\, \$19444%now\, \$18549%now\, \$v5468%now\, \$18604%now\, \$18540%now\, \$18575%now\, \$19330_compare6444359_id%now\, \$19085_modulo6684357_arg%now\, \$19040_modulo6684356_result%now\, \$19324_f0%now\, \$v5083%now\, \$19540%now\, \$v5817%now\, \$19554%now\, \$19295%now\, \$19120_res%now\, \$18475%now\, \$18580%now\, \$v4612%now\, \$19005_modulo6684349_arg%now\, \$v4518%now\, \$v5637%now\, \$18848%now\, \$19801%now\, \$18893_v%now\, \$19913%now\, \$19262_forever6704385_id%now\, \$19210_res%now\, \$v5169%now\, \$18514%now\, \$18747%now\, \$v5402%now\, \$v5090%now\, \$v4408%now\, \$19304%now\, \$v5523%now\, \$18505%now\, \$18888_next_acc%now\, \$19376_b%now\, \$18688%now\, \$19100_modulo6684349_arg%now\, \$19412_sp%now\, \$v4407%now\, \$v5447%now\, \$19798%now\, \$v5003%now\, \$v5873%now\, \$19097_modulo6684356_arg%now\, \$v5550%now\, \$19626%now\, \$19471%now\, \$18721%now\, \$18971_modulo6684357_id%now\, \$18797_branch_if648_id%now\, \$v4704%now\, \$19288_v%now\, \$v5390%now\, \$19366_compbranch6504391_result%now\, \$v5462%now\, \$19914%now\, \$v5311%now\, \$18608%now\, \$19317%now\, \$19141_modulo6684356_result%now\, \$18511%now\, \$v4671%now\, \$19487%now\, \$18522_loop665_arg%now\, \$v4420%now\, \$19625%now\, \$v5576%now\, \$19886%now\, \$v5482%now\, \result4928%now\, \$19773%now\, \$v4424%now\, \$19787%now\, \$19104_modulo6684357_result%now\, \$v5769%now\, \$19496_aux664_result%now\, \$19717%now\, \$18647%now\, \$19155%now\, \$18661%now\, \$v4587%now\, \$19939%now\, \$18832_v%now\, \$19227%now\, \$19650%now\, \$18495%now\, \$18551%now\, \$v5658%now\, \$19276%now\, \$19859%now\, \$19325%now\, \$18977_binop_int6434365_result%now\, \$18944_r%now\, \$18527%now\, \$19119_v%now\, \$18648%now\, \$19793%now\, \$18877_v%now\, \$18939_binop_int6434363_id%now\, \$v5673%now\, \$19190_binop_compare6454380_id%now\, \$19842%now\, \$19144_modulo6684349_id%now\, \$v5536%now\, \$v5299%now\, \$19601_copy_root_in_ram6634352_arg%now\, \$18539%now\, \$18936_modulo6684349_id%now\, \$19015_binop_int6434367_result%now\, \$19171_compare6444358_id%now\, \$19597%now\, \$19581%now\, \$v4338%now\, \$19384_compare6444359_result%now\, \$19748%now\, \$18522_loop665_id%now\, \$18461%now\, \$19256_v%now\, \$v5206%now\, \$18824_v%now\, \$v5059%now\, \$18657%now\, \$v5026%now\, \$v4996%now\, \$v5036%now\, \$18825%now\, \$18806%now\, \$v4866%now\, \$v4647%now\, \$18891%now\, \$18843%now\, \$v4330%now\, \$19370_compare6444359_id%now\, \$19601_copy_root_in_ram6634352_id%now\, \$v5281%now\, \$v4546%now\, \$v4779%now\, \$v4636%now\, \$v4812%now\, \$v5574%now\, \$18526_aux664_arg%now\, \$19308_v%now\, \$18793_make_block579_arg%now\, \$18437_loop666_arg%now\, \$19206_binop_compare6454382_result%now\, \$18444%now\, \$19066_modulo6684357_id%now\, \$19046_r%now\, \$19837%now\, \$v5429%now\, \$19571%now\, \$v4978%now\, \$v4920%now\, \$v5799%now\, \$18524_loop666_arg%now\, \$18810%now\, \$19944%now\, \$18880%now\, \$18869%now\, \$v5490%now\, \$18659%now\, \$v5257%now\, \$18945_modulo6684356_id%now\, \$18683_hd%now\, \$v4428%now\, \$v5055%now\, \$19774%now\, \$v5522%now\, \$19783%now\, \$19125_modulo6684349_result%now\, \$19097_modulo6684356_id%now\, \$19507_next%now\, \rdy4400%now\, \$19542%now\, \$v5042%now\, \$18813%now\, \$19220%now\, \$v4667%now\, \$v4678%now\, \$19211_compare6444358_result%now\, \$18790_loop666_result%now\, \$19804%now\, \$18622%now\, \$v4519%now\, \$19667%now\, \$v4593%now\, \$19811_copy_root_in_ram6634341_arg%now\, \$18695%now\, \$19789_next%now\, \$19259%now\, \$18437_loop666_id%now\, \$19203_compare6444358_id%now\, \$19788%now\, \$19141_modulo6684356_arg%now\, \$18473%now\, \$v5134%now\, \$19144_modulo6684349_result%now\, \$19932%now\, \$18603%now\, \$v5365%now\, \$19701%now\, \$19543%now\, \$v5168%now\, \$v4529%now\, \$v4839%now\, \$v4679%now\, \$19796%now\, \$18845%now\, \$v5233%now\, \$18438_loop665_arg%now\, \$19337_compare6444359_arg%now\, \$v4632%now\, \$v4957%now\, \$19336_b%now\, \$19709%now\, \$19031_modulo6684349_result%now\, \$19824_hd%now\, \$19619%now\, \$18546%now\, \$v5872%now\, \$19818%now\, \$18971_modulo6684357_arg%now\, \$v4502%now\, \$19326_compbranch6504387_id%now\, \$18531%now\, \$v4802%now\, \$18841%now\, \$v4639%now\, \$19466_sp%now\, \$18567%now\, \$v4683%now\, \$19643_w%now\, \$18649%now\, \$18929_modulo6684349_arg%now\, \$v5184%now\, \$v4335%now\, \$v5915%now\, \$19169_v%now\, \$v5487%now\, \$v5552%now\, \$19361_fill6544390_id%now\, \$v5811%now\, \$19512%now\, \$v4471%now\, \$19725%now\, \$19844%now\, \$18732%now\, \$18618%now\, \$19387_compbranch6504394_arg%now\, \$19027_r%now\, \$v5471%now\, \$19659_hd%now\, \$19875%now\, \$19639%now\, \$18470%now\, \$19310%now\, \$19815%now\, \$v5696%now\, \$19350_v%now\, \$19503%now\, \$19182_binop_compare6454379_result%now\, \$18955_modulo6684349_result%now\, \$18476%now\, \$18443%now\, \$19230_v%now\, \$19018_v%now\, \$19713%now\, \$19218_v%now\, \$19009_modulo6684357_arg%now\, \$19498_loop665_result%now\, \$v5198%now\, \$19741%now\, \$v4581%now\, \$19161%now\, \$19156%now\, \$19104_modulo6684357_arg%now\, \$18492%now\, \$v5571%now\, \$v4615%now\, \$19937%now\, \$18917_modulo6684349_arg%now\, \$v5384%now\, \$18939_binop_int6434363_arg%now\, \$19572%now\, \$18898%now\, \$19391_compare6444359_result%now\, \$v5563%now\, \$18948_modulo6684349_id%now\, \$v5897%now\, \$19100_modulo6684349_id%now\, \$19409_sp%now\, \$18478%now\, \$19047_modulo6684357_result%now\, \$19009_modulo6684357_result%now\, \$v5072%now\, \$18895_v%now\, \$18559_copy_root_in_ram6634347_id%now\, \$18559_copy_root_in_ram6634347_arg%now\, \$19922%now\, \$19125_modulo6684349_id%now\, \$18629%now\, \$v4887%now\, \$v4556%now\, \$v5453%now\, \$19731%now\, \$19449%now\, \$18669%now\, \$18660%now\, \rdy4573%now\, \$18795_offsetclosure_n639_id%now\, \$19401_compbranch6504396_arg%now\, \$19878%now\, \$v5066%now\, \$18631%now\, \$v4327%now\, \$19234_sp%now\, \$18687%now\, \$19811_copy_root_in_ram6634341_result%now\, \rdy4608%now\, \$19728%now\, \$v5492%now\, \$19843%now\, \$19532_forever6704350_arg%now\, \$19028_modulo6684357_id%now\, \$18958_binop_int6434364_arg%now\, \$v4700%now\, \$19301_v%now\, \$v4940%now\, \$19012_modulo6684349_result%now\, \$19268%now\, \$19772%now\, \$19226%now\, \$v5727%now\, \$18889_v%now\, \$19882%now\, \$19877%now\, \$19091_binop_int6434371_id%now\, \$v4796%now\, \$18907_modulo6684356_result%now\, \$19561%now\, \$19282_v%now\, \$19806%now\, \$19257_v%now\, \$19660%now\, \$18583_w%now\, \$v4818%now\, \$v4750%now\, \$19492%now\, \$18525_loop665_id%now\, \$19311%now\, \$19743%now\, \$v4775%now\, \$v4713%now\, \$19519%now\, \$19870%now\, \$v4540%now\, \$19638%now\, \$v4821%now\, \$v5664%now\, \$19211_compare6444358_arg%now\, \$18500%now\, \$18545_next%now\, \$19078_modulo6684356_result%now\, \$19868%now\, \$19047_modulo6684357_id%now\, \$18663%now\, \$18679%now\, \$19053_binop_int6434369_result%now\, \$v4937%now\, \$v5305%now\, \$18986_modulo6684349_result%now\, \$19266%now\, \$19447_sp%now\, \$19084_r%now\, \$19779_loop666_result%now\, \$v5825%now\, \$18464_rdy%now\, \$19636%now\, \$19329_b%now\, \$v5596%now\, \$19031_modulo6684349_id%now\, \$19526_forever6704355_id%now\, \$19926%now\, \$19614_hd%now\, \$19594%now\, \$18542_next%now\, \$18553_forever6704348_id%now\, \$19521%now\, \$19832%now\, \$v4455%now\, \$v4640%now\, \$19053_binop_int6434369_arg%now\, \$18508%now\, \$19684%now\, \$19315%now\, \$19166_binop_compare6454377_id%now\, \$19110%now\, \$19678%now\, \$v5405%now\, \$v5622%now\, \$v5188%now\, \$v5138%now\, \$19198_binop_compare6454381_result%now\, \$v4972%now\, \$19872%now\, \$19031_modulo6684349_arg%now\, \$19405_compare6444359_arg%now\, \$v4754%now\, \$v5254%now\, \$v5275%now\, \$18642%now\, \$19892%now\, \$v4339%now\, \$v4532%now\, \$v5260%now\, \$19021_modulo6684356_arg%now\, \$18996_binop_int6434366_result%now\, \$19005_modulo6684349_id%now\, \$18522_loop665_result%now\, \$18682_w%now\, \$18914_modulo6684357_id%now\, \$18673%now\, \$19766%now\, \$v4558%now\, \$19214%now\, \$19566%now\, \$v4337%now\, \$v5096%now\, \$v5359%now\, \$19174_binop_compare6454378_result%now\, \$19563%now\, \$v4606%now\, \$v5141%now\, \$18639%now\, \$19154%now\, \$18562%now\, \$v4449%now\, \$v4605%now\, \$v4539%now\, \$18666%now\, \$19781_aux664_id%now\, \$18904_v%now\, \$18498%now\, \$v4562%now\, \$19497_loop666_arg%now\, \$18564%now\, \$v5335%now\, \$19834%now\, \$19700%now\, \$19769%now\, \$19907%now\, \$18724%now\, \$19425%now\, \$19293%now\, \$19147_r%now\, \$19950%now\, \$19355%now\, \$19024_modulo6684349_id%now\, \$19665%now\, \$19351%now\, \$19500%now\, \$v4833%now\, \$v4791%now\, \$v4746%now\, \$v5524%now\, \$19856%now\, \$18456%now\, \$19021_modulo6684356_result%now\, \$v5560%now\, \$v4751%now\, \$18487%now\, \$19755%now\, \$19233%now\, \$18654%now\, \$v4911%now\, \$v5743%now\, \$19414%now\, \$19649%now\, \$18702%now\, \$18897%now\, \$v4496%now\, \$18967_modulo6684349_result%now\, \$v5477%now\, \$v4675%now\, \$v5107%now\, \$19485%now\, \$v5597%now\, \$19132_modulo6684349_arg%now\, \$18781%now\, \$19252_forever6704384_id%now\, \$v4984%now\, \$v5753%now\, \$18896_v%now\, \$18737%now\, \$18439_wait662_result%now\, \$v5102%now\, \$v4813%now\, \$v5432%now\, \$19642%now\, \$18446_dur%now\, \$18625_copy_root_in_ram6634345_id%now\, \$v5314%now\, \$v5540%now\, \$19617%now\, \$19451%now\, \$18556_forever6704344_id%now\, \$19585%now\, \$18886%now\, \$18439_wait662_id%now\, \$v5441%now\, \$19737%now\, \$19879%now\, \$19072_binop_int6434370_id%now\, \$19462%now\, \$18516%now\, \$18838_v%now\, \$v5502%now\, \$v5814%now\, \$v5845%now\, \$18438_loop665_result%now\, \$19658_w%now\, \$19182_binop_compare6454379_arg%now\, \$18901_binop_int6434361_result%now\, \$18453%now\, \$19260%now\, \$v5605%now\, \$18971_modulo6684357_result%now\, \$19853%now\, \$v5131%now\, \$18820_v%now\, \$18571_copy_root_in_ram6634345_result%now\, \$18515%now\, \$v4689%now\, \$18914_modulo6684357_result%now\, \$v5497%now\, \$19951%now\, \$19807%now\, \$19241_v%now\, \$19242%now\, \$19539%now\, \$18752%now\, \$v5544%now\, \result4607%now\, \$19091_binop_int6434371_arg%now\, \$19345%now\, \$v5491%now\, \$18844%now\, \$18963_r%now\, \$v5652%now\, \$v5876%now\, \$19113_forever6704372_id%now\, \$19383_b%now\, \$19584%now\, \$19942%now\, \$19615%now\, \$18676%now\, \$v4514%now\, \$19316%now\, \$19148_modulo6684357_id%now\, \$v4492%now\, \$v5347%now\, \$v5411%now\, \$18756%now\, \$19865_w%now\, \$18533%now\, \$19297_v%now\, \$18497%now\, \$19062_modulo6684349_arg%now\, \$19456%now\, \$v5909%now\, \$v5356%now\, \$v5584%now\, \$v5023%now\, \$18766%now\, \$19770%now\, \$v4960%now\, \$18674%now\, \$18595%now\, \$19927%now\, \$v5293%now\, \$v5525%now\, \$18786%now\, \$19592%now\, \$18748%now\, \$18448_dis%now\, \$19398_compare6444359_result%now\, \$19202_res%now\, \$18951_r%now\, \$19040_modulo6684356_arg%now\, \$v5724%now\, \$18780%now\, \$18651%now\, \$19518_next%now\, \$19005_modulo6684349_result%now\, \$18808%now\, \$18715%now\, \$19799%now\, \$v5505%now\, \$v5867%now\, \$19646%now\, \$19833%now\, \$19182_binop_compare6454379_id%now\, \$v5000%now\, \$v5185%now\, \$v5034%now\, \$18467_loop665_result%now\, \$v5222%now\, \$v4782%now\, \$19547_copy_root_in_ram6634352_id%now\, \$19915%now\, \$19719%now\, \$18777%now\, \$18550%now\, \$18842%now\, \$18489%now\, \$18439_wait662_arg%now\, \$19100_modulo6684349_result%now\, \$19135_binop_int6434374_id%now\, \$18796_make_block_n646_arg%now\, \$v5084%now\, \$v4654%now\, \$19820%now\, \$18901_binop_int6434361_arg%now\, \$18701%now\, \$18768_w%now\, \$19586%now\, \$v5709%now\, \$18613_copy_root_in_ram6634346_arg%now\, \$19917%now\, \$19138_v%now\, \$19697%now\, \$v4423%now\, \result4963%now\, \$18794_apply638_arg%now\, \$18792_wait662_arg%now\, \$18741%now\, \$18735%now\, \$v5039%now\, \$19677%now\, \$v5296%now\, \$18714%now\, \$19231%now\, \$v5689%now\, \$v5251%now\, \$19876%now\, \$v5606%now\, \$v5670%now\, \$18794_apply638_result%now\, \$19921%now\, \$19420_w06554397_id%now\, \$v4719%now\, \$19059_modulo6684356_id%now\, \$19864%now\, \$19347_fill6534389_result%now\, \$v5099%now\, \$19860%now\, \$19781_aux664_arg%now\, \$v4827%now\, \$18964_modulo6684356_arg%now\, \$v5802%now\, \$v4917%now\, \$19302%now\, \$v5368%now\, \$19823_w%now\, \$v5494%now\, \$19668%now\, \$19398_compare6444359_id%now\, \$18574%now\, \$19228_v%now\, \$v5079%now\, \$19749%now\, \$19795%now\, \$19203_compare6444358_arg%now\, \$19768%now\, \$v4809%now\, \$19941%now\, \$v4902%now\, \$18899%now\, \$19605%now\, \$19514%now\, \$v4836%now\, \$18640%now\, \$v4716%now\, \$v5396%now\, \$19341%now\, \$18870_v%now\, \$19722%now\, \$19475%now\, \$v5353%now\, \$v4953%now\, \$19460%now\, \$19470%now\, \$19580%now\, \$19893%now\, \$v4597%now\, \$v5051%now\, \$v5679%now\, \$v5630%now\, \$19889%now\, \$18812%now\, \$v5543%now\, \$18955_modulo6684349_id%now\, \$19529_forever6704351_arg%now\, \$v5556%now\, \$19497_loop666_result%now\, \$18536%now\, \$19433%now\, \$v4857%now\, \$19286%now\, \$19621%now\, \$18758%now\, \$19261%now\, \$v5566%now\, \$v4881%now\, \$19148_modulo6684357_result%now\, \$v4795%now\, \$19945%now\, \$v4466%now\, \$v4824%now\, \$19747%now\, \$19081_modulo6684349_id%now\, \$19285%now\, \$v4884%now\, \$v5863%now\, \$19394_compbranch6504395_result%now\, \$19535_copy_root_in_ram6634354_result%now\, \$v4758%now\, \$v4488%now\, \$19012_modulo6684349_arg%now\, \$18607%now\, \$19753%now\, \$18785%now\, \$19394_compbranch6504395_id%now\, \$v5894%now\, \$18799_w1656_arg%now\, \$18856_loop_push6494360_id%now\, \$v4981%now\, \$19391_compare6444359_arg%now\, \$19366_compbranch6504391_id%now\, \$v4771%now\, \$19781_aux664_result%now\, \$19174_binop_compare6454378_id%now\, \$19416_w36574398_arg%now\, \$v5627%now\, \$19271%now\, \$v5126%now\, \$18708%now\, \$19780_loop665_id%now\, \$18827%now\, \$v5890%now\, \$18882_v%now\, \$18525_loop665_arg%now\, \$v5623%now\, \$19344%now\, \$19576%now\, \$19171_compare6444358_arg%now\, \$19838_copy_root_in_ram6634340_id%now\, \$v5387%now\, \$19373_compbranch6504392_arg%now\, \$v5602%now\, \$18544%now\, \$v5773%now\, \$18493%now\, \$18579%now\, \$v5444%now\, \$19524%now\, \$19247%now\, \$19122_modulo6684356_id%now\, \$v5585%now\, \$19494_loop666_result%now\, \$19284%now\, \$19373_compbranch6504392_id%now\, \$19287_v%now\, \$19808_forever6704342_id%now\, \$v5459%now\, \$19767%now\, \$v5181%now\, \$19494_loop666_id%now\, \$19529_forever6704351_id%now\, \$v5782%now\, \$19053_binop_int6434369_id%now\, \$v4478%now\, \$v5495%now\, \$v4505%now\, \$18621%now\, \$19598%now\, \$v4774%now\, \$18523_aux664_result%now\, \$v5919%now\, \$19298_v%now\, \$18872_v%now\, \$18817_v%now\, \$19762%now\, \$19002_modulo6684356_id%now\, \$v5695%now\, \$v5770%now\, \$19024_modulo6684349_arg%now\, \$18936_modulo6684349_result%now\, \$19428%now\, \$18890_v%now\, \$v5561%now\, \$18535%now\, \$19151_modulo6684349_arg%now\, \result4399%now\, \$19278%now\, \rdy4435%now\, \$19000_res%now\, \$18609%now\, \$18720%now\, \$19552%now\, \$18757%now\, \$v4459%now\, \$19305%now\, \$18874%now\, \$18800%now\, \$19607%now\, \$v4557%now\, \$19757%now\, \$v4536%now\, \$19933_w%now\, \$v4487%now\, \$19258%now\, \$v4720%now\, \$19151_modulo6684349_id%now\, \$19744_w%now\, \result4572%now\, \$19103_r%now\, \$v5562%now\, \$19178_res%now\, \$19160%now\, \$19663%now\, \$18871%now\, \$v5332%now\, \$v5045%now\, \$19193_v%now\, \$v4670%now\, \$v5880%now\, \$v5030%now\, \$18883_v%now\, \$v4333%now\, \$v5572%now\, \$18983_modulo6684356_result%now\, \$19493%now\, \$19095_res%now\, \$v5756%now\, \$18983_modulo6684356_arg%now\, \$v5114%now\, \$v5192%now\, \$19461%now\, \$19107_modulo6684349_result%now\, \$18839%now\, \$v5341%now\, \$v5626%now\, \$19050_modulo6684349_id%now\, \$18787%now\, \$18716%now\, \$19121_r%now\, \$19206_binop_compare6454382_id%now\, \$18885_v%now\, \$18658%now\, \$v5851%now\, \$19069_modulo6684349_result%now\, \$v5111%now\, \$18678%now\, \$19822%now\, \$v5510%now\, \$18753%now\, \$v5848%now\, \$19113_forever6704372_arg%now\, \$18840_v%now\, \$v5362%now\, \$v4905%now\, \$18596%now\, \$v4553%now\, \$v5218%now\, \$18440_make_block579_result%now\, \$19401_compbranch6504396_id%now\, \$19380_compbranch6504393_result%now\, \$19047_modulo6684357_arg%now\, \$18861%now\, \$19931%now\, \$19340_argument2%now\, \$v4991%now\, \$18983_modulo6684356_id%now\, \$v5591%now\, \$v5211%now\, \$18920_binop_int6434362_id%now\, \$v5531%now\, \$19002_modulo6684356_result%now\, \$v4890%now\, \$18589%now\, \$19144_modulo6684349_arg%now\, \$v4600%now\, \$19476_v%now\, \$19587%now\, \$19919%now\, \$19574_w%now\, \$19237_v%now\, \$19037_v%now\, \$v5483%now\, \$19634%now\, \$18585%now\, \$v4432%now\, \$19365%now\, \$v5736%now\, \$v4332%now\, \$19857%now\, \$v5868%now\, \$18803%now\, \$19346_sp%now\, \$18691%now\, \$19846%now\, \$v5841%now\, \$19695%now\, \$19494_loop666_arg%now\, \$v5177%now\, \$v4707%now\, \$19122_modulo6684356_arg%now\, \$v4737%now\, \$v5712%now\, \$19370_compare6444359_arg%now\, \$19622%now\, \$v4567%now\, \$v5500%now\, \$19899%now\, \$v5918%now\, \$v5408%now\, \$19039_r%now\, \$18814%now\, \$19738%now\, \$19670%now\, \$19457%now\, \$19377_compare6444359_id%now\, \$19556%now\, \$19711%now\, \$v5808%now\, \$19377_compare6444359_arg%now\, \$19405_compare6444359_result%now\, \$v5593%now\, \$19903_next%now\, \$18818_v%now\, \$18633%now\, \$18466_loop666_arg%now\, \$19459%now\, \$19705%now\, \$19629_hd%now\, \$18836_v%now\, \$19384_compare6444359_arg%now\, \$18736%now\, \$v5110%now\, \$18671%now\, \$18686%now\, \$v4526%now\, \$18990_modulo6684357_arg%now\, \$v5493%now\, \$19632%now\, \$v5871%now\, \$18823_v%now\, \$18593%now\, \$v5229%now\, \$v5302%now\, \$18652_w%now\, \$19506%now\, \$19337_compare6444359_result%now\, \$v4411%now\, \$19680%now\, \rdy4964%now\, \$18690%now\, \$v4755%now\, \$v5615%now\, \$19195_compare6444358_id%now\, \$19912%now\, \$18469_make_block579_arg%now\, \$18743%now\, \$19791%now\, \$19604%now\, \$v5805%now\, \$19510%now\, \$18728%now\, \$19869%now\, \$19900%now\, \$19898%now\, \$19111%now\, \$18586%now\, \$18986_modulo6684349_id%now\, \$18468_wait662_id%now\, \$19244_v%now\, \$19612%now\, \$v4785%now\, \$19847%now\, \$19398_compare6444359_arg%now\, \$v4987%now\, \$19830%now\, \$19034_binop_int6434368_id%now\, \$18856_loop_push6494360_result%now\, \$19687_w%now\, \$19745_hd%now\, \$18894_v%now\, \$v5887%now\, \$18672%now\, \$18617%now\, \$19938%now\, \$18892_v%now\, \$19437%now\, \$18636%now\, \$18611%now\, \$19225%now\, \$19420_w06554397_arg%now\, \$18713%now\, \$18616%now\, \$18771%now\, \$v4635%now\, \$v5792%now\, \$18868_v%now\, \$v5106%now\, \$18693%now\, \$18597%now\, \$18437_loop666_result%now\, \$19426%now\, \$19763%now\, \$v5575%now\, \$v4747%now\, \$v5381%now\, \$19151_modulo6684349_result%now\, \$v5474%now\, \$18850%now\, \$18445_x%now\, \$18798_w652_arg%now\, \$18878%now\, \$v5820%now\, \$v5022%now\, \$v4968%now\, \$v4686%now\, \$19472%now\, \$v5718%now\, \$19404_b%now\, \$v4446%now\, \$19624%now\, \$18587%now\, \$v5906%now\, \$18970_r%now\, \$19545%now\, \$18534_next%now\, \$19219%now\, \$18792_wait662_id%now\, \$19265_ofs%now\, \$19618%now\, \$19411%now\, \$19468_sp%now\, \$18547%now\, \$19116_binop_int6434373_id%now\, \$19065_r%now\, \$19645%now\, \$19129_modulo6684357_result%now\, \$v5155%now\, \$v5219%now\, \$19756%now\, \$18490%now\, \$18523_aux664_arg%now\, \$v5375%now\, \$19215_argument1%now\, \$18860%now\, \$v5898%now\, \$v4643%now\, \$19174_binop_compare6454378_arg%now\, \$v5581%now\, \$v4999%now\, \$18466_loop666_result%now\, \$18469_make_block579_result%now\, \$18625_copy_root_in_ram6634345_result%now\, \$19640%now\, \$v4657%now\, \$v5501%now\, \$19323%now\, \$v5631%now\, \$19270%now\, \$19473%now\, \$19318%now\, \$19132_modulo6684349_result%now\, \$18548%now\, \$18967_modulo6684349_id%now\, \$18772%now\, \$18628%now\, \$19562%now\, \$18538%now\, \$18819_v%now\, \$19198_binop_compare6454381_arg%now\, \$19465_sp%now\, \$18526_aux664_result%now\, \$19911%now\, \$v4914%now\, \$19446_sp%now\, \$18932_r%now\, \$v4463%now\, \$19946%now\, \$19943%now\, \$v5372%now\, \$19577%now\, \$18641%now\, \$18773%now\, \$v5740%now\, \$18524_loop666_id%now\, \$18964_modulo6684356_result%now\, \$v4427%now\, \$19655%now\, \$19028_modulo6684357_arg%now\, \$v4788%now\, \$19520%now\, \$v4875%now\, \$19306_v%now\, \$v5567%now\, \$v5521%now\, \$v4644%now\, \$19343_sp%now\, \$18722%now\, \$19935%now\, \$19056_v%now\, \$18513%now\, \$18989_r%now\, \$18879_v%now\, \$v4956%now\, \$19730%now\, \$18665%now\, \$v4452%now\, \$v5783%now\, \$18710%now\, \$v5676%now\, \$19009_modulo6684357_id%now\, \$19712%now\, \$19841%now\, \$18556_forever6704344_arg%now\, \$19780_loop665_result%now\, \$19236_v%now\, \$19330_compare6444359_result%now\, \$v5600%now\, \$19330_compare6444359_arg%now\, \$18592%now\, \$19289%now\, \$19589_copy_root_in_ram6634353_arg%now\, \$v4778%now\, \$19356%now\, \$19050_modulo6684349_arg%now\, \$v5241%now\, \$18594%now\, \$v5680%now\, \$18866_v%now\, \$v5877%now\, \$19424%now\, \$v5587%now\, \$19369_b%now\, \$18481%now\, \$19050_modulo6684349_result%now\, \$19691%now\, \$18471%now\, \$19058_r%now\, \$19560_hd%now\, \$19405_compare6444359_id%now\, \$v5901%now\, \$v5435%now\, \$19353%now\, \$19059_modulo6684356_result%now\, \$18910_modulo6684349_arg%now\, \$v5706%now\, \$18486%now\, \$18501%now\, \$18532%now\, \$v4764%now\, \$19216_v%now\, \$19613_w%now\, \$18528%now\, \$19283%now\, \$v5338%now\, \$19091_binop_int6434371_result%now\, \$v4962%now\, \$19654%now\, \$v5842%now\, \$v5527%now\, \$18920_binop_int6434362_result%now\, \$19195_compare6444358_arg%now\, \$v5910%now\, \$18705_next%now\, \$19511%now\, \$v5902%now\, \$19410%now\, \$18468_wait662_arg%now\, \$v5504%now\, \$v4522%now\, \$18797_branch_if648_arg%now\, \$19696%now\, \$18955_modulo6684349_arg%now\, \$19652%now\, \$19606%now\, \$19195_compare6444358_result%now\, \$v5006%now\, \$18804%now\, \$18910_modulo6684349_result%now\, \$19502%now\, \$v5583%now\, \$18853_hd%now\, \$v5746%now\, \$v5048%now\, \$19831%now\, \$19481%now\, \$18774%now\, \$19708%now\, \$18632%now\, \$18625_copy_root_in_ram6634345_arg%now\, \$v5834%now\, \$19568%now\, \$v4723%now\, \$18519%now\, \$v4580%now\, \$19547_copy_root_in_ram6634352_arg%now\, \$19477_v%now\, \$18704%now\, \$18503%now\, \$18790_loop666_arg%now\, \$v5854%now\, \$19690%now\, \$v5786%now\, \$19498_loop665_id%now\, \$v5864%now\, \$v5886%now\, \$18923_v%now\, \$v5914%now\, \$v5798%now\, \$v5016%now\, \$19499_aux664_result%now\, \$v5554%now\, \$18675%now\, \$18463%now\, \$19469%now\, \$18700%now\, \$18744_w%now\, \$v5087%now\, \$18530%now\, \$v5423%now\, \$v5215%now\, \$18929_modulo6684349_result%now\, \$19733%now\, \$18653_hd%now\, \$19429%now\, \$18833%now\, \$v5165%now\, \$18454%now\, \$18847%now\, \$v5553%now\, \$v5075%now\, \$18692%now\, \$18719%now\, \$19940%now\, \$18712_hd%now\, \$v5417%now\, \$19125_modulo6684349_arg%now\, \$18634%now\, \$19484%now\, \$18929_modulo6684349_id%now\, \$19198_binop_compare6454381_id%now\, \$19416_w36574398_id%now\, \$18798_w652_id%now\, \$v5056%now\, \$v4439%now\, \$v5503%now\, \$19608%now\, \$v5779%now\, \$19277%now\, \$19223%now\, \$18499%now\, \$18796_make_block_n646_result%now\, \$19085_modulo6684357_id%now\, \$v5399%now\, \$v4808%now\, \$18811%now\, \$19808_forever6704342_arg%now\, \$v4508%now\, \$v5207%now\, \$v5093%now\, \$19034_binop_int6434368_result%now\, \$19627%now\, \$19881_hd%now\, \$19291_v%now\, \$18901_binop_int6434361_id%now\, \$19387_compbranch6504394_result%now\, \$19644_hd%now\, \$19347_fill6534389_id%now\, \$v5917%now\, \$19792%now\, \$19541%now\, \$v5480%now\, \$19415_sp%now\, \$19262_forever6704385_arg%now\, \$18477%now\, \$19635%now\, \$v4933%now\, \$19633%now\, \$v4566%now\, \$18917_modulo6684349_id%now\, \$18451%now\, \$19802%now\, \$19221%now\, \$19224%now\, \$v5240%now\, \$19516%now\, \$18656%now\, \$19693%now\, \$18496%now\, \$18588%now\, \$18887_v%now\, \$19360_sp%now\, \$19171_compare6444358_result%now\, \$19688_hd%now\, \$18491%now\, \$18541%now\, \$19380_compbranch6504393_arg%now\, \$19782%now\, \$v5517%now\, \$19141_modulo6684356_id%now\, \$19107_modulo6684349_id%now\, \$v4971%now\, \$v4848%now\, \$19166_binop_compare6454377_result%now\, \$19593%now\, \$18568%now\, \$v4625%now\, \$18452%now\, \$19742%now\, \$v4869%now\, \$v5590%now\, \$18468_wait662_result%now\, \$19575_hd%now\, \$19229_v%now\, \$18981_res%now\, \$v4622%now\, \$18942_v%now\, \$18543%now\, \$19513%now\, \$19555%now\, \$19692%now\, \$19370_compare6444359_result%now\, \$v4896%now\, \$v5661%now\, \$v5520%now\, \$18917_modulo6684349_result%now\, \$19116_binop_int6434373_result%now\, \$v4404%now\, \$19862%now\, \$18449%now\, \$19573%now\, \$19729%now\, \$18952_modulo6684357_id%now\, \$19252_forever6704384_arg%now\, \$19805%now\, \$18943_res%now\, \$v4564%now\, \$18926_modulo6684356_arg%now\, \$v5438%now\, \$19567%now\, \$18761%now\, \$v5350%now\, \$v5230%now\, \$v4731%now\, \$19838_copy_root_in_ram6634340_arg%now\, \$v5667%now\, \$v5535%now\, \$19008_r%now\, \$v5547%now\, \$19669%now\, \$18862%now\, \$19699%now\, \$19630%now\, \$ram_lock%now\, \$global_end_lock%now\, \$code_lock%now\)
        variable \$18463\ : value(0 to 1) := (others => '0');
        variable \$19410\, \$18469_make_block579_result\, 
                 \$19420_w06554397_arg\, \$18440_make_block579_result\, 
                 \$19344\, \$18525_loop665_arg\, \$19231\, 
                 \$18438_loop665_arg\, \$18522_loop665_arg\, \$19444\, 
                 \$19498_loop665_arg\, \$18467_loop665_arg\, 
                 \$18791_loop665_arg\, \$19780_loop665_arg\, 
                 \$19495_loop665_arg\, \$19358\, 
                 \$18793_make_block579_result\ : value(0 to 95) := (others => '0');
        variable \$19195_compare6444358_arg\, \$19330_compare6444359_arg\, 
                 \$19398_compare6444359_arg\, \$19384_compare6444359_arg\, 
                 \$19377_compare6444359_arg\, \$19370_compare6444359_arg\, 
                 \$19171_compare6444358_arg\, \$19391_compare6444359_arg\, 
                 \$19203_compare6444358_arg\, \$19405_compare6444359_arg\, 
                 \$19211_compare6444358_arg\, \$19337_compare6444359_arg\, 
                 \$19187_compare6444358_arg\, \$19179_compare6444358_arg\ : value(0 to 93) := (others => '0');
        variable \$19742\, \$19608\, \$18632\, \$18532\, \$19506\, \$19931\, 
                 \$18448_dis\, \$18766\, \$18533\, \$19462\, \$19907\, 
                 \$19818\, \$19788\, \$19542\, \$19787\, \$19554\, \$19718\, 
                 \$19463\, \$18742\, \$19505\, \$19596\, \$18566\, \$19845\, 
                 \$18709\, \$18620\, \$18578\, \$19685\, \$19464\ : value(0 to 47) := (others => '0');
        variable \$18790_loop666_arg\, \$18523_aux664_arg\, 
                 \$18798_w652_arg\, \$18466_loop666_arg\, 
                 \$19494_loop666_arg\, \$19781_aux664_arg\, 
                 \$19497_loop666_arg\, \$18524_loop666_arg\, 
                 \$18437_loop666_arg\, \$18526_aux664_arg\, 
                 \$19499_aux664_arg\, \$18856_loop_push6494360_arg\, 
                 \$19779_loop666_arg\, \$19238_w6514383_arg\, 
                 \$19496_aux664_arg\, \$18521_loop666_arg\ : value(0 to 63) := (others => '0');
        variable \$18452\, \$18451\, \$18454\, \$v5902\, \$v5910\, \$v5898\, 
                 \$v5906\, \$18453\, \$18456\, \$18455\ : value(0 to 7) := (others => '0');
        variable \$18797_branch_if648_arg\, \$18787\, \$18789\, \$18788\ : value(0 to 122) := (others => '0');
        variable \$18541\, \$19360_sp\, \$19415_sp\, \$19499_aux664_result\, 
                 \$18705_next\, \$19780_loop665_result\, \$19343_sp\, 
                 \$19446_sp\, \$18526_aux664_result\, \$19465_sp\, 
                 \$18625_copy_root_in_ram6634345_result\, \$19468_sp\, 
                 \$19265_ofs\, \$18534_next\, 
                 \$18856_loop_push6494360_result\, \$19903_next\, 
                 \$19346_sp\, \$18523_aux664_result\, \$19781_aux664_result\, 
                 \$19535_copy_root_in_ram6634354_result\, \$19514\, 
                 \$19347_fill6534389_result\, \$18467_loop665_result\, 
                 \$19518_next\, \$18571_copy_root_in_ram6634345_result\, 
                 \$18438_loop665_result\, \$18522_loop665_result\, 
                 \$18542_next\, \$19447_sp\, \$18545_next\, 
                 \$19811_copy_root_in_ram6634341_result\, \$19234_sp\, 
                 \$19409_sp\, \$19498_loop665_result\, \$19466_sp\, \$19796\, 
                 \$19789_next\, \$19507_next\, \$19496_aux664_result\, 
                 \$19412_sp\, \$19420_w06554397_result\, 
                 \$19589_copy_root_in_ram6634353_result\, \$18854_sp\, 
                 \$19467_sp\, \$18613_copy_root_in_ram6634346_result\, 
                 \$19361_fill6544390_result\, 
                 \$19601_copy_root_in_ram6634352_result\, 
                 \$18791_loop665_result\, \$19238_w6514383_result\, 
                 \$18525_loop665_result\, \$19681_next\, 
                 \$19547_copy_root_in_ram6634352_result\, 
                 \$18559_copy_root_in_ram6634347_result\, \$19800_next\, 
                 \$19495_loop665_result\, \$19515_next\, 
                 \$19838_copy_root_in_ram6634340_result\, \$19714_next\, 
                 \$19797_next\, \$18738_next\, \$19416_w36574398_result\ : value(0 to 15) := (others => '0');
        variable \$18926_modulo6684356_arg\, \$19125_modulo6684349_arg\, 
                 \$18955_modulo6684349_arg\, \$18910_modulo6684349_arg\, 
                 \$19050_modulo6684349_arg\, \$19028_modulo6684357_arg\, 
                 \$18990_modulo6684357_arg\, \$19122_modulo6684356_arg\, 
                 \$19144_modulo6684349_arg\, \$19047_modulo6684357_arg\, 
                 \$18983_modulo6684356_arg\, \$19151_modulo6684349_arg\, 
                 \$19024_modulo6684349_arg\, \$19012_modulo6684349_arg\, 
                 \$18964_modulo6684356_arg\, \$19040_modulo6684356_arg\, 
                 \$19062_modulo6684349_arg\, \$19132_modulo6684349_arg\, 
                 \$19021_modulo6684356_arg\, \$19031_modulo6684349_arg\, 
                 \$18917_modulo6684349_arg\, \$19104_modulo6684357_arg\, 
                 \$19009_modulo6684357_arg\, \$18929_modulo6684349_arg\, 
                 \$18971_modulo6684357_arg\, \$19141_modulo6684356_arg\, 
                 \$19097_modulo6684356_arg\, \$19100_modulo6684349_arg\, 
                 \$19005_modulo6684349_arg\, \$19085_modulo6684357_arg\, 
                 \$19148_modulo6684357_arg\, \$19078_modulo6684356_arg\, 
                 \$19107_modulo6684349_arg\, \$19129_modulo6684357_arg\, 
                 \$18907_modulo6684356_arg\, \$19069_modulo6684349_arg\, 
                 \$19059_modulo6684356_arg\, \$19088_modulo6684349_arg\, 
                 \$18952_modulo6684357_arg\, \$18933_modulo6684357_arg\, 
                 \$19066_modulo6684357_arg\, \$18936_modulo6684349_arg\, 
                 \$18967_modulo6684349_arg\, \$19043_modulo6684349_arg\, 
                 \$18948_modulo6684349_arg\, \$18914_modulo6684357_arg\, 
                 \$18993_modulo6684349_arg\, \$18986_modulo6684349_arg\, 
                 \$19002_modulo6684356_arg\, \$18974_modulo6684349_arg\, 
                 \$19081_modulo6684349_arg\, \$18945_modulo6684356_arg\ : value(0 to 61) := (others => '0');
        variable \$18468_wait662_arg\, \$18792_wait662_arg\, 
                 \$18439_wait662_arg\ : value(0 to 96) := (others => '0');
        variable result4399 : value(0 to 57) := (others => '0');
        variable \$v4564\, \$v4566\, \$v4567\, \$18443\, \$18462\, \$v4565\, 
                 \$v4568\, \$v4563\ : value(0 to 3) := (others => '0');
        variable \$19380_compbranch6504393_arg\, 
                 \$19373_compbranch6504392_arg\, 
                 \$19401_compbranch6504396_arg\, 
                 \$19387_compbranch6504394_arg\, 
                 \$19366_compbranch6504391_arg\, 
                 \$19326_compbranch6504387_arg\, 
                 \$19333_compbranch6504388_arg\, 
                 \$19394_compbranch6504395_arg\ : value(0 to 215) := (others => '0');
        variable \$18952_modulo6684357_id\, \$19107_modulo6684349_id\, 
                 \$19141_modulo6684356_id\, \$18917_modulo6684349_id\, 
                 \$19347_fill6534389_id\, \$18901_binop_int6434361_id\, 
                 \$19085_modulo6684357_id\, \$18798_w652_id\, 
                 \$19416_w36574398_id\, \$19198_binop_compare6454381_id\, 
                 \$18929_modulo6684349_id\, \$19498_loop665_id\, 
                 \$19405_compare6444359_id\, \$19009_modulo6684357_id\, 
                 \$18524_loop666_id\, \$18967_modulo6684349_id\, 
                 \$19116_binop_int6434373_id\, \$18792_wait662_id\, 
                 \$19034_binop_int6434368_id\, \$18468_wait662_id\, 
                 \$18986_modulo6684349_id\, \$19195_compare6444358_id\, 
                 \$19377_compare6444359_id\, \$18920_binop_int6434362_id\, 
                 \$18983_modulo6684356_id\, \$19401_compbranch6504396_id\, 
                 \$19206_binop_compare6454382_id\, \$19050_modulo6684349_id\, 
                 \$19151_modulo6684349_id\, \$19002_modulo6684356_id\, 
                 \$19053_binop_int6434369_id\, \$19529_forever6704351_id\, 
                 \$19494_loop666_id\, \$19808_forever6704342_id\, 
                 \$19373_compbranch6504392_id\, \$19122_modulo6684356_id\, 
                 \$19838_copy_root_in_ram6634340_id\, \$19780_loop665_id\, 
                 \$19174_binop_compare6454378_id\, 
                 \$19366_compbranch6504391_id\, \$18856_loop_push6494360_id\, 
                 \$19394_compbranch6504395_id\, \$19081_modulo6684349_id\, 
                 \$18955_modulo6684349_id\, \$19398_compare6444359_id\, 
                 \$19059_modulo6684356_id\, \$19420_w06554397_id\, 
                 \$19135_binop_int6434374_id\, 
                 \$19547_copy_root_in_ram6634352_id\, 
                 \$19182_binop_compare6454379_id\, \$19148_modulo6684357_id\, 
                 \$19113_forever6704372_id\, \$19072_binop_int6434370_id\, 
                 \$18439_wait662_id\, \$18556_forever6704344_id\, 
                 \$18625_copy_root_in_ram6634345_id\, 
                 \$19252_forever6704384_id\, \$19024_modulo6684349_id\, 
                 \$19781_aux664_id\, \$18914_modulo6684357_id\, 
                 \$19005_modulo6684349_id\, \$19166_binop_compare6454377_id\, 
                 \$18553_forever6704348_id\, \$19526_forever6704355_id\, 
                 \$19031_modulo6684349_id\, \$19047_modulo6684357_id\, 
                 \$18525_loop665_id\, \$19091_binop_int6434371_id\, 
                 \$19028_modulo6684357_id\, \$18795_offsetclosure_n639_id\, 
                 \$19125_modulo6684349_id\, 
                 \$18559_copy_root_in_ram6634347_id\, 
                 \$19100_modulo6684349_id\, \$18948_modulo6684349_id\, 
                 \$19361_fill6544390_id\, \$19326_compbranch6504387_id\, 
                 \$19203_compare6444358_id\, \$18437_loop666_id\, 
                 \$19097_modulo6684356_id\, \$18945_modulo6684356_id\, 
                 \$19066_modulo6684357_id\, 
                 \$19601_copy_root_in_ram6634352_id\, 
                 \$19370_compare6444359_id\, \$18522_loop665_id\, 
                 \$19171_compare6444358_id\, \$18936_modulo6684349_id\, 
                 \$19144_modulo6684349_id\, \$19190_binop_compare6454380_id\, 
                 \$18939_binop_int6434363_id\, \$18797_branch_if648_id\, 
                 \$18971_modulo6684357_id\, \$19262_forever6704385_id\, 
                 \$19330_compare6444359_id\, \$19497_loop666_id\, 
                 \$18794_apply638_id\, \$19238_w6514383_id\, 
                 \$18526_aux664_id\, \$19532_forever6704350_id\, 
                 \$19043_modulo6684349_id\, \$18990_modulo6684357_id\, 
                 \$18799_w1656_id\, \$19333_compbranch6504388_id\, 
                 \$19320_forever6704386_id\, \$18958_binop_int6434364_id\, 
                 \$18907_modulo6684356_id\, \$18790_loop666_id\, 
                 \$18964_modulo6684356_id\, \$18977_binop_int6434365_id\, 
                 \$18996_binop_int6434366_id\, \$19012_modulo6684349_id\, 
                 \$19088_modulo6684349_id\, \$19021_modulo6684356_id\, 
                 \$18993_modulo6684349_id\, \$19384_compare6444359_id\, 
                 \$19179_compare6444358_id\, \$19078_modulo6684356_id\, 
                 \$19211_compare6444358_id\, 
                 \$18571_copy_root_in_ram6634345_id\, 
                 \$18796_make_block_n646_id\, \$18521_loop666_id\, 
                 \$19387_compbranch6504394_id\, 
                 \$19535_copy_root_in_ram6634354_id\, 
                 \$19391_compare6444359_id\, \$19337_compare6444359_id\, 
                 \$18613_copy_root_in_ram6634346_id\, \$19495_loop665_id\, 
                 \$19157_forever6704375_id\, \$19062_modulo6684349_id\, 
                 \$18466_loop666_id\, \$18926_modulo6684356_id\, 
                 \$19187_compare6444358_id\, \$19163_forever6704376_id\, 
                 \$19015_binop_int6434367_id\, 
                 \$19811_copy_root_in_ram6634341_id\, 
                 \$18793_make_block579_id\, \$19129_modulo6684357_id\, 
                 \$19589_copy_root_in_ram6634353_id\, 
                 \$19040_modulo6684356_id\, \$19104_modulo6684357_id\, 
                 \$19499_aux664_id\, \$19132_modulo6684349_id\, 
                 \$19380_compbranch6504393_id\, \$18933_modulo6684357_id\, 
                 \$18974_modulo6684349_id\, \$19779_loop666_id\, 
                 \$19069_modulo6684349_id\, \$18910_modulo6684349_id\ : value(0 to 11) := (others => '0');
        variable \$19008_r\, \$18943_res\, \$18917_modulo6684349_result\, 
                 \$18981_res\, \$18929_modulo6684349_result\, 
                 \$18910_modulo6684349_result\, 
                 \$19059_modulo6684356_result\, \$19058_r\, 
                 \$19050_modulo6684349_result\, \$v5783\, \$18989_r\, 
                 \$18964_modulo6684356_result\, \$18932_r\, 
                 \$19132_modulo6684349_result\, \$19215_argument1\, 
                 \$19129_modulo6684357_result\, \$19065_r\, \$18970_r\, 
                 \$19151_modulo6684349_result\, \$19039_r\, 
                 \$19002_modulo6684356_result\, \$19340_argument2\, 
                 \$19069_modulo6684349_result\, \$19121_r\, 
                 \$19107_modulo6684349_result\, \$19095_res\, 
                 \$18983_modulo6684356_result\, \$19103_r\, \$19000_res\, 
                 \$18936_modulo6684349_result\, \$v5770\, 
                 \$19148_modulo6684357_result\, \$19433\, 
                 \$19100_modulo6684349_result\, 
                 \$19005_modulo6684349_result\, \$18951_r\, \$18963_r\, 
                 \$18914_modulo6684357_result\, 
                 \$18971_modulo6684357_result\, \$v5753\, 
                 \$18967_modulo6684349_result\, 
                 \$19021_modulo6684356_result\, \$19147_r\, \$19084_r\, 
                 \$19266\, \$18986_modulo6684349_result\, 
                 \$19078_modulo6684356_result\, 
                 \$18907_modulo6684356_result\, 
                 \$19012_modulo6684349_result\, 
                 \$19009_modulo6684357_result\, 
                 \$19047_modulo6684357_result\, 
                 \$18955_modulo6684349_result\, \$19027_r\, 
                 \$19031_modulo6684349_result\, 
                 \$19144_modulo6684349_result\, 
                 \$19125_modulo6684349_result\, \$v5799\, \$19046_r\, 
                 \$18944_r\, \$19104_modulo6684357_result\, 
                 \$19141_modulo6684356_result\, \$19120_res\, 
                 \$19040_modulo6684356_result\, \$18925_r\, \$19038_res\, 
                 \$19057_res\, \$18926_modulo6684356_result\, \$19441_arg\, 
                 \$19077_r\, \$19020_r\, \$19097_modulo6684356_result\, 
                 \$19128_r\, \$19019_res\, \$18905_res\, 
                 \$18948_modulo6684349_result\, \$18982_r\, \$19096_r\, 
                 \$18816\, \$18933_modulo6684357_result\, \$18962_res\, 
                 \$19408_argument3\, \$18913_r\, \$18906_r\, \$19139_res\, 
                 \$18952_modulo6684357_result\, 
                 \$19081_modulo6684349_result\, 
                 \$19088_modulo6684349_result\, 
                 \$19062_modulo6684349_result\, \$19076_res\, 
                 \$18974_modulo6684349_result\, \$v5760\, 
                 \$19066_modulo6684357_result\, \$19427\, 
                 \$19043_modulo6684349_result\, 
                 \$18990_modulo6684357_result\, 
                 \$19028_modulo6684357_result\, \$18924_res\, 
                 \$19122_modulo6684356_result\, \$19001_r\, \$19140_r\, 
                 \$19024_modulo6684349_result\, 
                 \$18993_modulo6684349_result\, 
                 \$19085_modulo6684357_result\, \$18945_modulo6684356_result\ : value(0 to 30) := (others => '0');
        variable \$18795_offsetclosure_n639_arg\ : value(0 to 137) := (others => '0');
        variable \$18793_make_block579_arg\ : value(0 to 103) := (others => '0');
        variable \$18469_make_block579_arg\, result4963, result4607, 
                 result4434, \$18440_make_block579_arg\ : value(0 to 127) := (others => '0');
        variable \$19630\, \$19699\, \$18862\, \$19669\, \$v5535\, \$v5667\, 
                 \$v4731\, \$v5230\, \$v5350\, \$19567\, \$v5438\, \$19805\, 
                 \$19252_forever6704384_arg\, \$19729\, \$19573\, \$19862\, 
                 \$v4404\, \$v5520\, \$v5661\, \$v4896\, 
                 \$19370_compare6444359_result\, \$19692\, \$19555\, 
                 \$19513\, \$18543\, \$v4622\, \$v5590\, \$v4869\, \$v4625\, 
                 \$18568\, \$19593\, \$v4848\, \$v4971\, \$19782\, \$18491\, 
                 \$19171_compare6444358_result\, \$18588\, \$18496\, 
                 \$19693\, \$18656\, \$19516\, \$v5240\, \$19224\, \$19221\, 
                 \$19802\, \$19633\, \$v4933\, \$19635\, \$18477\, 
                 \$19262_forever6704385_arg\, \$v5480\, \$19792\, \$v5917\, 
                 \$19627\, \$v5093\, \$v5207\, \$v4508\, 
                 \$19808_forever6704342_arg\, \$18811\, \$v4808\, \$v5399\, 
                 \$18499\, \$19223\, \$19277\, \$v5779\, \$v5503\, \$v4439\, 
                 \$v5056\, \$19484\, \$18634\, \$v5417\, \$19940\, \$18719\, 
                 \$18692\, \$v5075\, \$v5553\, \$18847\, \$v5165\, \$18833\, 
                 \$19429\, \$19733\, \$v5215\, \$v5423\, \$18530\, \$v5087\, 
                 \$18700\, \$18675\, \$v5554\, \$v5016\, \$v5798\, \$v5914\, 
                 \$v5886\, \$v5864\, \$v5786\, \$19690\, \$v5854\, \$18503\, 
                 \$v4580\, \$v4723\, \$19568\, \$v5834\, \$19708\, \$18774\, 
                 \$19481\, \$19831\, \$v5048\, \$v5746\, \$v5583\, \$19502\, 
                 \$18804\, \$v5006\, \$19195_compare6444358_result\, 
                 \$19606\, \$19652\, \$19696\, \$v4522\, \$v5504\, \$19511\, 
                 \$v5842\, \$19654\, \$v4962\, \$v5338\, \$19283\, \$18528\, 
                 \$v4764\, \$18501\, \$18486\, \$v5706\, \$v5435\, \$v5901\, 
                 \$18471\, \$19691\, \$18481\, \$19369_b\, \$19424\, 
                 \$v5877\, \$v5680\, \$18594\, \$v5241\, \$v4778\, \$19289\, 
                 \$18592\, \$v5600\, \$19330_compare6444359_result\, 
                 \$18556_forever6704344_arg\, \$19841\, \$19712\, \$v5676\, 
                 \$18710\, \$v4452\, \$18665\, \$19730\, \$v4956\, \$18513\, 
                 \$19935\, \$18722\, \$v4644\, \$v5521\, \$v4875\, \$19520\, 
                 \$v4788\, \$19655\, \$v4427\, \$v5740\, \$18773\, \$18641\, 
                 \$19577\, \$v5372\, \$19943\, \$19946\, \$v4463\, \$v4914\, 
                 \$19911\, \$18538\, \$19562\, \$18628\, \$18772\, \$18548\, 
                 \$19318\, \$19473\, \$19270\, \$19323\, \$v5501\, \$v4657\, 
                 \$19640\, \$18466_loop666_result\, \$v4999\, \$v5581\, 
                 \$v4643\, \$18860\, \$v5375\, \$18490\, \$19756\, \$v5219\, 
                 \$v5155\, \$19645\, \$18547\, \$19411\, \$19618\, \$19219\, 
                 \$19545\, \$18587\, \$19624\, \$v4446\, \$19404_b\, 
                 \$v5718\, \$19472\, \$v4686\, \$v4968\, \$v5022\, \$v5820\, 
                 \$18878\, \$18445_x\, \$v5474\, \$v5381\, \$v4747\, 
                 \$v5575\, \$19426\, \$18437_loop666_result\, \$18597\, 
                 \$18693\, \$v5106\, \$v5792\, \$v4635\, \$18771\, \$18616\, 
                 \$18713\, \$19225\, \$18611\, \$18636\, \$19938\, \$18617\, 
                 \$18672\, \$v5887\, \$19830\, \$v4987\, \$19847\, \$v4785\, 
                 \$19612\, \$18586\, \$19111\, \$19898\, \$19900\, \$19869\, 
                 \$19510\, \$v5805\, \$19604\, \$19791\, \$18743\, \$19912\, 
                 \$v4755\, \$18690\, rdy4964, \$v4411\, 
                 \$19337_compare6444359_result\, \$v5302\, \$v5229\, 
                 \$18593\, \$19632\, \$v5493\, \$v4526\, \$18686\, \$18671\, 
                 \$v5110\, \$18736\, \$19705\, \$19459\, \$18633\, \$v5593\, 
                 \$19405_compare6444359_result\, \$v5808\, \$19711\, 
                 \$19556\, \$19457\, \$19670\, \$19738\, \$18814\, \$v5408\, 
                 \$v5918\, \$19899\, \$v5500\, \$19622\, \$v5712\, \$v4737\, 
                 \$v4707\, \$v5177\, \$19695\, \$v5841\, \$19846\, \$18691\, 
                 \$18803\, \$19857\, \$v4332\, \$v5736\, \$19365\, \$v4432\, 
                 \$18585\, \$19634\, \$v5483\, \$19919\, \$19587\, \$v4600\, 
                 \$18589\, \$v4890\, \$v5531\, \$v5211\, \$v5591\, \$v4991\, 
                 \$18861\, \$v5218\, \$v4553\, \$18596\, \$v4905\, \$v5362\, 
                 \$19113_forever6704372_arg\, \$v5848\, \$18753\, \$v5510\, 
                 \$19822\, \$18678\, \$v5111\, \$v5851\, \$18658\, \$18716\, 
                 \$v5626\, \$v5341\, \$18839\, \$19461\, \$v5192\, \$v5114\, 
                 \$v5756\, \$v5572\, \$v4333\, \$v5030\, \$v5880\, \$v4670\, 
                 \$v5045\, \$v5332\, \$18871\, \$19663\, \$19160\, 
                 \$19178_res\, \$v5562\, result4572, \$v4720\, \$19258\, 
                 \$v4487\, \$v4536\, \$19757\, \$v4557\, \$18800\, \$18874\, 
                 \$19305\, \$v4459\, \$18757\, \$19552\, \$18720\, \$18609\, 
                 rdy4435, \$19278\, \$v5561\, \$19428\, \$v5695\, \$19762\, 
                 \$v5919\, \$v4774\, \$19598\, \$18621\, \$v4505\, \$v5495\, 
                 \$v4478\, \$v5782\, \$v5181\, \$19767\, \$v5459\, \$19284\, 
                 \$19494_loop666_result\, \$v5585\, \$19247\, \$19524\, 
                 \$v5444\, \$18579\, \$18493\, \$v5773\, \$18544\, \$v5602\, 
                 \$v5387\, \$19576\, \$v5890\, \$18827\, \$v5126\, \$19271\, 
                 \$v4771\, \$v4981\, \$v5894\, \$19753\, \$18607\, \$v4488\, 
                 \$v4758\, \$v5863\, \$v4884\, \$19285\, \$19747\, \$v4824\, 
                 \$v4466\, \$19945\, \$v4795\, \$v4881\, \$v5566\, \$19261\, 
                 \$18758\, \$19621\, \$19286\, \$v4857\, \$18536\, 
                 \$19497_loop666_result\, \$v5556\, 
                 \$19529_forever6704351_arg\, \$v5543\, \$18812\, \$19889\, 
                 \$v5630\, \$v5679\, \$v5051\, \$v4597\, \$19893\, \$19580\, 
                 \$19470\, \$19460\, \$v4953\, \$v5353\, \$19475\, \$19722\, 
                 \$19341\, \$v5396\, \$v4716\, \$18640\, \$v4836\, \$19605\, 
                 \$18899\, \$v4902\, \$19941\, \$v4809\, \$19768\, \$19795\, 
                 \$19749\, \$v5079\, \$18574\, \$19668\, \$v5494\, \$v5368\, 
                 \$19302\, \$v4917\, \$v5802\, \$v4827\, \$19860\, \$v5099\, 
                 \$19864\, \$v4719\, \$19921\, \$v5670\, \$v5606\, \$19876\, 
                 \$v5251\, \$v5689\, \$18714\, \$v5296\, \$19677\, \$v5039\, 
                 \$18735\, \$v4423\, \$19697\, \$19917\, \$v5709\, \$19586\, 
                 \$18701\, \$19820\, \$v4654\, \$v5084\, \$18489\, \$18550\, 
                 \$18777\, \$19719\, \$19915\, \$v4782\, \$v5222\, \$v5034\, 
                 \$v5185\, \$v5000\, \$19833\, \$19646\, \$v5867\, \$v5505\, 
                 \$19799\, \$18715\, \$18808\, \$18651\, \$18780\, \$v5724\, 
                 \$19202_res\, \$19398_compare6444359_result\, \$18748\, 
                 \$19592\, \$18786\, \$v5525\, \$v5293\, \$19927\, \$18595\, 
                 \$18674\, \$v4960\, \$v5023\, \$v5584\, \$v5356\, \$v5909\, 
                 \$19456\, \$18497\, \$18756\, \$v5411\, \$v5347\, \$v4492\, 
                 \$19316\, \$v4514\, \$18676\, \$19615\, \$19942\, \$19584\, 
                 \$19383_b\, \$v5876\, \$v5652\, \$v5491\, \$19345\, 
                 \$v5544\, \$18752\, \$19539\, \$19242\, \$19807\, \$19951\, 
                 \$v4689\, \$18515\, \$v5131\, \$19853\, \$v5605\, \$19260\, 
                 \$v5845\, \$v5814\, \$v5502\, \$18516\, \$19879\, \$v5441\, 
                 \$18886\, \$19585\, \$19451\, \$19617\, \$v5540\, \$v5314\, 
                 \$19642\, \$v5432\, \$v4813\, \$v5102\, \$v4984\, \$18781\, 
                 \$v5107\, \$v4675\, \$v5477\, \$v4496\, \$18897\, \$18702\, 
                 \$19649\, \$19414\, \$v5743\, \$v4911\, \$18654\, \$19233\, 
                 \$19755\, \$18487\, \$v4751\, \$v5560\, \$19856\, \$v5524\, 
                 \$v4746\, \$v4791\, \$v4833\, \$19500\, \$19351\, \$19665\, 
                 \$19355\, \$19293\, \$19425\, \$18724\, \$19769\, \$19700\, 
                 \$19834\, \$v5335\, \$18564\, \$v4562\, \$18498\, \$18666\, 
                 \$v4539\, \$v4605\, \$v4449\, \$18562\, \$19154\, \$18639\, 
                 \$v5141\, \$v4606\, \$19563\, \$v5359\, \$v5096\, \$v4337\, 
                 \$19566\, \$19214\, \$v4558\, \$19766\, \$18673\, \$v5260\, 
                 \$v4532\, \$v4339\, \$19892\, \$18642\, \$v5275\, \$v5254\, 
                 \$v4754\, \$19872\, \$v4972\, \$v5138\, \$v5188\, \$v5622\, 
                 \$v5405\, \$19678\, \$19110\, \$19315\, \$18508\, \$v4640\, 
                 \$v4455\, \$19832\, \$19521\, \$19594\, \$v5596\, 
                 \$19329_b\, \$19636\, \$18464_rdy\, \$19779_loop666_result\, 
                 \$v5305\, \$v4937\, \$18679\, \$18663\, \$19868\, \$18500\, 
                 \$v5664\, \$v4821\, \$19638\, \$v4540\, \$19870\, \$19519\, 
                 \$v4713\, \$v4775\, \$19743\, \$v4750\, \$v4818\, \$19660\, 
                 \$19806\, \$19561\, \$v4796\, \$19877\, \$19882\, \$v5727\, 
                 \$19772\, \$19268\, \$v4940\, \$v4700\, 
                 \$19532_forever6704350_arg\, \$19843\, \$v5492\, \$19728\, 
                 rdy4608, \$18687\, \$v4327\, \$v5066\, \$19878\, rdy4573, 
                 \$18660\, \$18669\, \$19449\, \$19731\, \$v5453\, \$v4556\, 
                 \$v4887\, \$18629\, \$19922\, \$v5072\, \$18478\, \$v5897\, 
                 \$v5563\, \$19391_compare6444359_result\, \$18898\, 
                 \$19572\, \$v5384\, \$19937\, \$v4615\, \$v5571\, \$18492\, 
                 \$19156\, \$19161\, \$v4581\, \$v5198\, \$18476\, \$19503\, 
                 \$v5696\, \$19815\, \$19310\, \$18470\, \$19639\, \$19875\, 
                 \$v5471\, \$18618\, \$18732\, \$19725\, \$v4471\, \$19512\, 
                 \$v5811\, \$v5552\, \$v5915\, \$v4335\, \$v5184\, \$18649\, 
                 \$v4683\, \$18567\, \$v4639\, \$v4802\, \$18531\, \$v4502\, 
                 \$18546\, \$19619\, \$19709\, \$19336_b\, \$v4957\, 
                 \$v4632\, \$v5233\, \$18845\, \$v4679\, \$v4839\, \$v4529\, 
                 \$v5168\, \$19543\, \$19701\, \$v5365\, \$18603\, \$19932\, 
                 \$v5134\, \$18473\, \$19259\, \$18695\, \$v4593\, \$19667\, 
                 \$v4519\, \$18622\, \$19804\, \$18790_loop666_result\, 
                 \$19211_compare6444358_result\, \$v4678\, \$v4667\, 
                 \$18813\, \$v5042\, rdy4400, \$19783\, \$v5522\, \$19774\, 
                 \$v5055\, \$v4428\, \$v5257\, \$18659\, \$v5490\, \$18869\, 
                 \$18880\, \$19944\, \$18810\, \$v4920\, \$v4978\, \$19571\, 
                 \$v5429\, \$19837\, \$18444\, \$v5574\, \$v4812\, \$v4636\, 
                 \$v4779\, \$v4546\, \$v5281\, \$v4330\, \$18891\, \$v4647\, 
                 \$v4866\, \$18806\, \$18825\, \$v5036\, \$v4996\, \$v5026\, 
                 \$18657\, \$v5059\, \$v5206\, \$18461\, \$19748\, 
                 \$19384_compare6444359_result\, \$v4338\, \$19581\, 
                 \$19597\, \$18539\, \$v5299\, \$v5536\, \$19842\, \$v5673\, 
                 \$19793\, \$18648\, \$18527\, \$19325\, \$19859\, \$19276\, 
                 \$v5658\, \$18551\, \$18495\, \$19650\, \$19939\, \$v4587\, 
                 \$18661\, \$19155\, \$18647\, \$v5769\, \$v4424\, \$19773\, 
                 \$v5482\, \$19886\, \$v5576\, \$19625\, \$v4420\, \$19487\, 
                 \$v4671\, \$18511\, \$19317\, \$18608\, \$v5311\, \$19914\, 
                 \$v5462\, \$v5390\, \$v4704\, \$18721\, \$19471\, \$19626\, 
                 \$v5550\, \$v5003\, \$19798\, \$v5447\, \$v4407\, \$18688\, 
                 \$19376_b\, \$18505\, \$v5523\, \$19304\, \$v4408\, 
                 \$v5090\, \$v5402\, \$18747\, \$18514\, \$v5169\, 
                 \$19210_res\, \$19913\, \$19801\, \$v5637\, \$v4518\, 
                 \$v4612\, \$18580\, \$18475\, \$19295\, \$v5817\, \$19540\, 
                 \$v5083\, \$18575\, \$18540\, \$18604\, \$v5468\, \$18549\, 
                 \$19901\, \$18521_loop666_result\, \$v4651\, \$19888\, 
                 \$v4619\, \$19570\, \$v5344\, \$19582\, \$v4696\, \$18782\, 
                 \$19517\, \$19557\, \$18851\, \$19871\, \$19884\, \$v4872\, 
                 \$19836\, \$19275\, \$v4571\, \$19255\, \$19538\, \$19243\, 
                 \$19544\, \$19522\, \$v5103\, 
                 \$19179_compare6444358_result\, \$v4549\, \$19920\, 
                 \$v5199\, \$v5649\, \$19891\, \$v4442\, \$v5189\, \$v4767\, 
                 \$19546\, \$v5266\, \$19249\, \$18677\, \$19883\, \$v4458\, 
                 \$v4666\, \$18472\, rdy4929, \$19734\, \$18826\, \$19785\, 
                 \$18537\, \$19771\, \$19710\, \$v4431\, \$19637\, \$19664\, 
                 \$v5570\, \$19203_compare6444358_result\, 
                 \$19377_compare6444359_result\, \$v5007\, \$v5730\, 
                 \$v4899\, \$v5147\, \$v4495\, \$v5135\, \$18863\, \$19794\, 
                 \$18749\, \$18849\, \$v4860\, \$v4799\, \$v5618\, \$v5763\, 
                 \$v5080\, \$18494\, \$v5174\, \$19821\, \$v5393\, \$v5063\, 
                 \$v5225\, \$19320_forever6704386_arg\, \$v5573\, \$v5496\, 
                 \$19873\, \$19509\, \$18770\, \$19564\, \$19923\, \$19523\, 
                 \$v5010\, \$18681\, \$v5450\, \$v5789\, \$19352\, \$v4724\, 
                 \$19849\, \$18718\, \$18750\, \$v5161\, \$v5456\, \$v5031\, 
                 \$v5545\, \$18552\, \$18601\, \$19675\, \$v4570\, \$v5511\, 
                 \$v5601\, \$19936\, \$v5329\, \$v4893\, \$v5580\, \$v4851\, 
                 \$19162\, \$18798_w652_result\, \$18799_w1656_result\, 
                 \$19826\, \$19750\, \$18734\, \$v4475\, \$19671\, \$v5893\, 
                 \$18479\, \$v5534\, \$v4975\, \$19686\, \$19610\, \$19666\, 
                 \$v4792\, \$19616\, \$v4484\, \$18465\, \$v5512\, \$v5317\, 
                 \$v4943\, \$19588\, \$19835\, \$v4923\, \$v5565\, \$v5202\, 
                 \$v5795\, \$18755\, \$19694\, \$19631\, \$18689\, 
                 \$19186_res\, \$v5269\, \$19551\, \$19303\, \$18612\, 
                 \$v5272\, \$18779\, \$19858\, \$19908\, \$v5144\, \$19724\, 
                 \$v5546\, \$18459\, \$18725\, \$19786\, \$19861\, \$19483\, 
                 \$19647\, \$19438\, \$v5170\, \$v5148\, \$18717\, \$v4462\, 
                 \$19676\, \$v5737\, \$18829\, \$v5123\, \$18831\, \$v4699\, 
                 \$v5595\, \$v5130\, \$19651\, \$v5290\, \$v5203\, \$18746\, 
                 \$18488\, \$19746\, \$v4863\, \$19565\, \$v5542\, \$19313\, 
                 \$v5426\, \$19855\, \$v5180\, \$v5516\, \$19550\, \$v5485\, 
                 \$19397_b\, \$18754\, \$18643\, \$18553_forever6704348_arg\, 
                 \$v5533\, \$19852\, \$v5237\, \$v4414\, \$v5860\, \$18684\, 
                 \$v5069\, \$18610\, \$v5027\, \$v5614\, \$v5835\, \$v5263\, 
                 \$18570\, \$v5420\, \$v4543\, \$v5247\, \$v4328\, \$19918\, 
                 \$18460\, \$19825\, \$19754\, \$18623\, \$v5465\, \$19867\, 
                 \$19157_forever6704375_arg\, \$19751\, \$18680\, \$18699\, 
                 \$v4842\, \$19726\, \$v5555\, \$v5883\, \$18591\, \$v5564\, 
                 \$19474\, \$19488\, \$v5905\, \$v5284\, \$v5278\, \$19280\, 
                 \$19558\, \$18605\, \$19578\, \$19526_forever6704355_arg\, 
                 \$19599\, \$18864\, \$v4433\, \$v5195\, \$19679\, \$v4878\, 
                 \$19359\, \$18767\, \$19698\, \$v4584\, \$19413\, \$19662\, 
                 \$18510\, \$19727\, \$19390_b\, \$v4660\, \$18733\, 
                 \$18484\, \$v4601\, \$v4995\, \$v5308\, \$v4740\, \$v5831\, 
                 \$v5164\, \$v5823\, \$19569\, \$19269\, \$v5514\, \$v4805\, 
                 \$19887\, \$v5127\, \$v4680\, \$19814\, \$19232\, \$19848\, 
                 \$v4988\, \$19854\, \$v5120\, \$19648\, \$19251\, \$18635\, 
                 \$v4908\, \$18576\, \$v4695\, \$19897\, \$18645\, \$18563\, 
                 \$v5250\, \$v4674\, \$18644\, \$v5530\, \$19885\, \$19600\, 
                 \$v5244\, \$18600\, \$18662\, \$v5481\, \$v5702\, \$v4992\, 
                 \$18447\, \$v4417\, \$v4936\, \$18485\, \$18646\, \$18664\, 
                 \$v4946\, \$v5052\, \$19623\, \$v5378\, 
                 \$19187_compare6444358_result\, \$v4552\, \$v5060\, 
                 \$v5582\, \$v5603\, \$18685\, \$v5035\, \$v4631\, \$v4845\, 
                 \$19816\, \$v4761\, \$19248\, \$v5604\, \$18670\, \$18590\, 
                 \$v4596\, \$v4728\, \$18762\, \$19314\, \$v5640\, \$v4481\, 
                 \$18723\, \$v5838\, \$19583\, \$v5828\, \$19294\, \$v5655\, 
                 \$18458\, \$18480\, \$19656\, \$v4734\, \$v4727\, \$v4491\, 
                 \$v5210\, \$18815\, \$19609\, \$19732\, \$19434\, \$v4770\, 
                 \$18502\, \$19784\, \$19611\, \$19482\, \$v5749\, \$v4569\, 
                 \$v4523\, \$19829\, \$v4926\, \$v5506\, \$18703\, \$v4628\, 
                 \$v4854\, \$v5686\, \$19916\, \$18529\, \$v4692\, \$18482\, 
                 \$v5857\, \$19486\, \$v4949\, \$19217\, \$19803\, \$19620\, 
                 \$19657\, \$v5683\, \$v5610\, \$v4952\, \$v5646\, \$19319\, 
                 \$v5515\, \$19112\, \$18805\, \$18569\, \$18837\, \$18650\, 
                 \$19504\, \$18807\, \$v5019\, \$v5776\, \$19489\, \$19819\, 
                 \$19894\, \$v4616\, \$19752\, \$v5766\, \$v5234\, \$v5586\, 
                 \$19458\, \$v5721\, \$v5212\, \$v5320\, \$v5703\, \$19419\, 
                 \$v5759\, \$18694\, \$18778\, \$19723\, \$v4472\, 
                 \$18524_loop666_result\, \$v4590\, \$v4511\, \$19890\, 
                 \$18865\, \$v5752\, \$18867\, \$19445\, \$v5117\, \$v4830\, 
                 \$v5594\, \$v5151\, \$19653\, \$18876\, \$v4443\, \$v5414\, 
                 \$19661\, \$v5733\, \$v5369\, \$v5158\, \$19641\, \$18474\, 
                 \$v5692\, \$19672\, \$19947\, \$19194_res\, \$v5592\, 
                 \$18655\, \$v5323\, \$v4515\, \$18509\, \$19525\, \$v5013\, 
                 \$18582\, \$v5226\, \$v5551\, \$v4535\, \$18630\, \$19432\, 
                 \$19827\, \$19863\, \$19170_res\, \$v4814\, \$v4710\, 
                 \$18483\, \$v4703\, \$v5152\, \$19501\, \$v5532\, \$v5076\, 
                 \$18802\, \$v4577\, \$19689\, \$19245\, \$18696\, \$v4325\, 
                 \$v4470\, \$18900\, \$v4467\, \$v5287\, \$18581\, \$v5634\, 
                 \$19292\, \$v5699\, \$v4604\, \$19163_forever6704376_arg\, 
                 \$18776\, \$19758\, \$19579\, \$18835\, \$v4650\, \$18624\, 
                 \$19250\, \$v5643\, \$18504\, \$v5484\, \$v5326\, \$v4499\, 
                 \$v4961\, \$19828\, \$v5715\, \$19874\, \$18775\, \$18801\, 
                 \$18729\, \$v5513\, \$v5486\, \$19272\, \$18751\, \$18809\, 
                 \$v5541\, \$18602\, \$v5913\, \$v4663\, \$v5526\, \$19299\, 
                 \$v4743\, \$18606\ : value(0 to 0) := (others => '0');
        variable \$18794_apply638_arg\ : value(0 to 165) := (others => '0');
        variable \$18796_make_block_n646_arg\ : value(0 to 171) := (others => '0');
        variable \$19838_copy_root_in_ram6634340_arg\, 
                 \$18468_wait662_result\, 
                 \$19547_copy_root_in_ram6634352_arg\, 
                 \$18625_copy_root_in_ram6634345_arg\, 
                 \$19589_copy_root_in_ram6634353_arg\, \$18535\, 
                 \$19416_w36574398_arg\, \$18799_w1656_arg\, 
                 \$18613_copy_root_in_ram6634346_arg\, \$19770\, 
                 \$18439_wait662_result\, \$19485\, 
                 \$18559_copy_root_in_ram6634347_arg\, 
                 \$19811_copy_root_in_ram6634341_arg\, 
                 \$19601_copy_root_in_ram6634352_arg\, 
                 \$18792_wait662_result\, \$19790\, 
                 \$19535_copy_root_in_ram6634354_arg\, 
                 \$19361_fill6544390_arg\, 
                 \$18571_copy_root_in_ram6634345_arg\, 
                 \$19347_fill6534389_arg\, \$18512\, \$19508\ : value(0 to 79) := (others => '0');
        variable \$18519\, \$19493\, \$19492\, \$18520\, \$19778\, \$19777\ : value(0 to 128) := (others => '0');
        variable \$v5547\, \$18761\, \$18449\, \$18942_v\, \$19229_v\, 
                 \$19575_hd\, \$v5517\, \$19688_hd\, \$18887_v\, \$19541\, 
                 \$19644_hd\, \$19291_v\, \$19881_hd\, \$18712_hd\, 
                 \$18653_hd\, \$18744_w\, \$19469\, \$18923_v\, \$18704\, 
                 \$19477_v\, \$18853_hd\, \$v5527\, \$19613_w\, \$19216_v\, 
                 \$19353\, \$19560_hd\, \$v5587\, \$18866_v\, \$19356\, 
                 \$19236_v\, \$18879_v\, \$19056_v\, \$v5567\, \$19306_v\, 
                 \$18819_v\, \$v5631\, \$18850\, \$19763\, \$18868_v\, 
                 \$19437\, \$18892_v\, \$18894_v\, \$19745_hd\, \$19687_w\, 
                 \$19244_v\, \$18728\, \$v5615\, \$19680\, \$18652_w\, 
                 \$18823_v\, \$v5871\, \$18836_v\, \$19629_hd\, \$18818_v\, 
                 \$v5868\, \$19037_v\, \$19237_v\, \$19574_w\, \$19476_v\, 
                 \$18840_v\, \$18885_v\, \$18883_v\, \$19193_v\, \$19744_w\, 
                 \$19933_w\, \$19607\, \$18890_v\, \$18817_v\, \$18872_v\, 
                 \$19298_v\, \$19287_v\, \$v5623\, \$18882_v\, \$18708\, 
                 \$v5627\, \$18785\, \$18870_v\, \$19228_v\, \$19823_w\, 
                 \$18741\, \$19138_v\, \$18768_w\, \$18842\, \$19297_v\, 
                 \$19865_w\, \$18844\, \$19241_v\, \$v5497\, \$18820_v\, 
                 \$19658_w\, \$18838_v\, \$19737\, \$18446_dur\, \$18737\, 
                 \$18896_v\, \$v5597\, \$19950\, \$18904_v\, \$18682_w\, 
                 \$19684\, \$19614_hd\, \$19926\, \$v5825\, \$18583_w\, 
                 \$19257_v\, \$19282_v\, \$18889_v\, \$19226\, \$19301_v\, 
                 \$18631\, \$18895_v\, \$19741\, \$19218_v\, \$19713\, 
                 \$19018_v\, \$19230_v\, \$19350_v\, \$19659_hd\, \$19844\, 
                 \$v5487\, \$19169_v\, \$19643_w\, \$18841\, \$v5872\, 
                 \$19824_hd\, \$19220\, \$18683_hd\, \$19308_v\, \$18843\, 
                 \$18824_v\, \$19256_v\, \$18877_v\, \$19119_v\, \$19227\, 
                 \$18832_v\, \$19717\, \$19288_v\, \$v5873\, 
                 \$18888_next_acc\, \$18893_v\, \$18848\, \$19324_f0\, 
                 \$18442_cy\, \$18599_hd\, \$18884_v\, \$19559_w\, \$19595\, 
                 \$18873_v\, \$19354_v\, \$19307_v\, \$19880_w\, \$19910_hd\, 
                 \$v5611\, \$19177_v\, \$18598_w\, \$19423_v\, \$19075_v\, 
                 \$18765\, \$19357_v\, \$19909_w\, \$18830_v\, \$18711_w\, 
                 \$18450\, \$19761\, \$19450_v\, \$19222\, \$19851_hd\, 
                 \$v5870\, \$18980_v\, \$19279_v\, \$18577\, \$18822_v\, 
                 \$19312_v\, \$18999_v\, \$18584_hd\, \$18834_v\, \$19817\, 
                 \$v5557\, \$19267_hd\, \$v5577\, \$18828_v\, \$19721_hd\, 
                 \$18457\, \$19296_v\, \$v5607\, \$19246_v\, \$18638_hd\, 
                 \$19720_w\, \$18852\, \$18668_hd\, \$19628_w\, \$19902\, 
                 \$v5537\, \$18565\, \$18667_w\, \$19209_v\, \$19309_v\, 
                 \$19342\, \$v5869\, \$19478_v\, \$18745_hd\, \$19364_v\, 
                 \$19185_v\, \$19930\, \$19704\, \$19274_v\, \$19201_v\, 
                 \$18961_v\, \$19850_w\, \$18846\, \$19934_hd\, \$18859\, 
                 \$18855_next_env\, \$19906\, \$19235_v\, \$18881_hd\, 
                 \$v5824\, \$19094_v\, \$19448_v\, \$18821_v\, \$18769_hd\, 
                 \$19866_hd\, \$18619\, \$18875_v\, \$v5619\, \$18637_w\, 
                 \$19553\, \$v5507\ : value(0 to 31) := (others => '0');
        variable \$19198_binop_compare6454381_arg\, 
                 \$19174_binop_compare6454378_arg\, 
                 \$18901_binop_int6434361_arg\, 
                 \$19091_binop_int6434371_arg\, 
                 \$19182_binop_compare6454379_arg\, 
                 \$19053_binop_int6434369_arg\, \$19311\, 
                 \$18958_binop_int6434364_arg\, 
                 \$18939_binop_int6434363_arg\, \$19281\, 
                 \$19116_binop_int6434373_arg\, \$19300\, 
                 \$18920_binop_int6434362_arg\, 
                 \$19206_binop_compare6454382_arg\, 
                 \$18996_binop_int6434366_arg\, 
                 \$18977_binop_int6434365_arg\, 
                 \$19015_binop_int6434367_arg\, 
                 \$19034_binop_int6434368_arg\, 
                 \$19135_binop_int6434374_arg\, 
                 \$19166_binop_compare6454377_arg\, \$19273\, \$19290\, 
                 \$19072_binop_int6434370_arg\, 
                 \$19190_binop_compare6454380_arg\ : value(0 to 153) := (others => '0');
        variable \$19116_binop_int6434373_result\, 
                 \$19166_binop_compare6454377_result\, 
                 \$19387_compbranch6504394_result\, 
                 \$19034_binop_int6434368_result\, 
                 \$18796_make_block_n646_result\, 
                 \$18920_binop_int6434362_result\, 
                 \$19091_binop_int6434371_result\, 
                 \$19380_compbranch6504393_result\, 
                 \$19394_compbranch6504395_result\, \$18794_apply638_result\, 
                 \$18901_binop_int6434361_result\, 
                 \$19174_binop_compare6454378_result\, 
                 \$18996_binop_int6434366_result\, 
                 \$19198_binop_compare6454381_result\, 
                 \$19053_binop_int6434369_result\, 
                 \$19182_binop_compare6454379_result\, 
                 \$19206_binop_compare6454382_result\, 
                 \$19015_binop_int6434367_result\, 
                 \$18977_binop_int6434365_result\, result4928, 
                 \$19366_compbranch6504391_result\, 
                 \$19333_compbranch6504388_result\, 
                 \$19135_binop_int6434374_result\, 
                 \$19373_compbranch6504392_result\, 
                 \$18795_offsetclosure_n639_result\, 
                 \$19401_compbranch6504396_result\, 
                 \$19190_binop_compare6454380_result\, 
                 \$19072_binop_int6434370_result\, 
                 \$18958_binop_int6434364_result\, 
                 \$18797_branch_if648_result\, 
                 \$18939_binop_int6434363_result\, 
                 \$19326_compbranch6504387_result\ : value(0 to 121) := (others => '0');
        variable state : t_state;
        variable state_var5924 : t_state_var5924;
        variable state_var5923 : t_state_var5923;
        variable state_var5922 : t_state_var5922;
        variable state_var5921 : t_state_var5921;
        variable state_var5920 : t_state_var5920;
        variable \$ram_lock\ : value(0 to 0);
        variable \$global_end_lock\ : value(0 to 0);
        variable \$code_lock\ : value(0 to 0);
        
    begin
      \$18606\ := \$18606%now\;
      \$19190_binop_compare6454380_arg\ := \$19190_binop_compare6454380_arg%now\;
      \$v4743\ := \$v4743%now\;
      \$19072_binop_int6434370_arg\ := \$19072_binop_int6434370_arg%now\;
      \$18910_modulo6684349_id\ := \$18910_modulo6684349_id%now\;
      \$19299\ := \$19299%now\;
      \$19069_modulo6684349_id\ := \$19069_modulo6684349_id%now\;
      \$v5526\ := \$v5526%now\;
      \$v4663\ := \$v4663%now\;
      \$v5913\ := \$v5913%now\;
      \$18602\ := \$18602%now\;
      \$v5541\ := \$v5541%now\;
      \$18809\ := \$18809%now\;
      \$18751\ := \$18751%now\;
      \$19272\ := \$19272%now\;
      \$v5486\ := \$v5486%now\;
      \$v5513\ := \$v5513%now\;
      \$18729\ := \$18729%now\;
      \$v5507\ := \$v5507%now\;
      \$18801\ := \$18801%now\;
      \$19779_loop666_id\ := \$19779_loop666_id%now\;
      \$18775\ := \$18775%now\;
      \$19874\ := \$19874%now\;
      \$v5715\ := \$v5715%now\;
      \$18974_modulo6684349_id\ := \$18974_modulo6684349_id%now\;
      \$19828\ := \$19828%now\;
      \$v4961\ := \$v4961%now\;
      \$v4499\ := \$v4499%now\;
      \$19326_compbranch6504387_result\ := \$19326_compbranch6504387_result%now\;
      \$v5326\ := \$v5326%now\;
      \$v5484\ := \$v5484%now\;
      \$18504\ := \$18504%now\;
      \$v5643\ := \$v5643%now\;
      \$18945_modulo6684356_result\ := \$18945_modulo6684356_result%now\;
      \$18933_modulo6684357_id\ := \$18933_modulo6684357_id%now\;
      \$19250\ := \$19250%now\;
      \$18624\ := \$18624%now\;
      \$v4650\ := \$v4650%now\;
      \$19553\ := \$19553%now\;
      \$18637_w\ := \$18637_w%now\;
      \$19380_compbranch6504393_id\ := \$19380_compbranch6504393_id%now\;
      \$v5619\ := \$v5619%now\;
      \$18835\ := \$18835%now\;
      \$19579\ := \$19579%now\;
      \$19758\ := \$19758%now\;
      \$19085_modulo6684357_result\ := \$19085_modulo6684357_result%now\;
      \$18776\ := \$18776%now\;
      \$18875_v\ := \$18875_v%now\;
      \$19132_modulo6684349_id\ := \$19132_modulo6684349_id%now\;
      \$18619\ := \$18619%now\;
      \$19163_forever6704376_arg\ := \$19163_forever6704376_arg%now\;
      \$v4604\ := \$v4604%now\;
      \$v5699\ := \$v5699%now\;
      \$19292\ := \$19292%now\;
      \$v5634\ := \$v5634%now\;
      \$19416_w36574398_result\ := \$19416_w36574398_result%now\;
      \$18993_modulo6684349_result\ := \$18993_modulo6684349_result%now\;
      \$18581\ := \$18581%now\;
      \$19866_hd\ := \$19866_hd%now\;
      \$v5287\ := \$v5287%now\;
      \$v4467\ := \$v4467%now\;
      \$18900\ := \$18900%now\;
      \$v4470\ := \$v4470%now\;
      \$v4325\ := \$v4325%now\;
      \$18696\ := \$18696%now\;
      \$19245\ := \$19245%now\;
      \$19024_modulo6684349_result\ := \$19024_modulo6684349_result%now\;
      \$18945_modulo6684356_arg\ := \$18945_modulo6684356_arg%now\;
      \$19689\ := \$19689%now\;
      \$v4577\ := \$v4577%now\;
      \$19140_r\ := \$19140_r%now\;
      \$18802\ := \$18802%now\;
      \$v5076\ := \$v5076%now\;
      \$19001_r\ := \$19001_r%now\;
      \$v5532\ := \$v5532%now\;
      \$19501\ := \$19501%now\;
      \$18769_hd\ := \$18769_hd%now\;
      \$v5152\ := \$v5152%now\;
      \$v4703\ := \$v4703%now\;
      \$19122_modulo6684356_result\ := \$19122_modulo6684356_result%now\;
      \$19499_aux664_id\ := \$19499_aux664_id%now\;
      \$18483\ := \$18483%now\;
      \$19290\ := \$19290%now\;
      \$19273\ := \$19273%now\;
      \$19104_modulo6684357_id\ := \$19104_modulo6684357_id%now\;
      \$v4710\ := \$v4710%now\;
      \$v4814\ := \$v4814%now\;
      \$19170_res\ := \$19170_res%now\;
      \$18924_res\ := \$18924_res%now\;
      \$19863\ := \$19863%now\;
      \$18821_v\ := \$18821_v%now\;
      \$19827\ := \$19827%now\;
      \$19432\ := \$19432%now\;
      \$19448_v\ := \$19448_v%now\;
      \$18630\ := \$18630%now\;
      \$19094_v\ := \$19094_v%now\;
      \$v4535\ := \$v4535%now\;
      \$v5551\ := \$v5551%now\;
      \$19028_modulo6684357_result\ := \$19028_modulo6684357_result%now\;
      \$18939_binop_int6434363_result\ := \$18939_binop_int6434363_result%now\;
      \$v5824\ := \$v5824%now\;
      \$18788\ := \$18788%now\;
      \$v5226\ := \$v5226%now\;
      \$18582\ := \$18582%now\;
      \$19081_modulo6684349_arg\ := \$19081_modulo6684349_arg%now\;
      \$v5013\ := \$v5013%now\;
      \$18881_hd\ := \$18881_hd%now\;
      \$19525\ := \$19525%now\;
      \$18509\ := \$18509%now\;
      \$18793_make_block579_result\ := \$18793_make_block579_result%now\;
      \$18974_modulo6684349_arg\ := \$18974_modulo6684349_arg%now\;
      \$19235_v\ := \$19235_v%now\;
      \$v4515\ := \$v4515%now\;
      \$v5323\ := \$v5323%now\;
      \$18655\ := \$18655%now\;
      \$19906\ := \$19906%now\;
      \$v5592\ := \$v5592%now\;
      \$19194_res\ := \$19194_res%now\;
      \$18990_modulo6684357_result\ := \$18990_modulo6684357_result%now\;
      \$19947\ := \$19947%now\;
      \$19672\ := \$19672%now\;
      \$v5692\ := \$v5692%now\;
      \$18474\ := \$18474%now\;
      \$19641\ := \$19641%now\;
      \$18855_next_env\ := \$18855_next_env%now\;
      \$v5158\ := \$v5158%now\;
      \$19040_modulo6684356_id\ := \$19040_modulo6684356_id%now\;
      \$v5369\ := \$v5369%now\;
      \$v5733\ := \$v5733%now\;
      \$19661\ := \$19661%now\;
      \$v5414\ := \$v5414%now\;
      \$v4443\ := \$v4443%now\;
      \$18876\ := \$18876%now\;
      \$19653\ := \$19653%now\;
      \$19508\ := \$19508%now\;
      \$19358\ := \$19358%now\;
      \$v5151\ := \$v5151%now\;
      \$v5594\ := \$v5594%now\;
      \$19043_modulo6684349_result\ := \$19043_modulo6684349_result%now\;
      \$18859\ := \$18859%now\;
      \$v4830\ := \$v4830%now\;
      \$v5117\ := \$v5117%now\;
      \$19445\ := \$19445%now\;
      \$18867\ := \$18867%now\;
      \$v5752\ := \$v5752%now\;
      \$18865\ := \$18865%now\;
      \$19890\ := \$19890%now\;
      \$v4511\ := \$v4511%now\;
      \$18455\ := \$18455%now\;
      \$18512\ := \$18512%now\;
      \$v4590\ := \$v4590%now\;
      \$19427\ := \$19427%now\;
      \$19934_hd\ := \$19934_hd%now\;
      \$18846\ := \$18846%now\;
      \$18524_loop666_result\ := \$18524_loop666_result%now\;
      \$v4472\ := \$v4472%now\;
      \$19723\ := \$19723%now\;
      \$18778\ := \$18778%now\;
      \$18694\ := \$18694%now\;
      \$v5759\ := \$v5759%now\;
      \$19066_modulo6684357_result\ := \$19066_modulo6684357_result%now\;
      \$19850_w\ := \$19850_w%now\;
      \$19419\ := \$19419%now\;
      \$18961_v\ := \$18961_v%now\;
      \$19201_v\ := \$19201_v%now\;
      \$v5703\ := \$v5703%now\;
      \$19274_v\ := \$19274_v%now\;
      \$19394_compbranch6504395_arg\ := \$19394_compbranch6504395_arg%now\;
      \$v5320\ := \$v5320%now\;
      \$19166_binop_compare6454377_arg\ := \$19166_binop_compare6454377_arg%now\;
      \$v5212\ := \$v5212%now\;
      \$19704\ := \$19704%now\;
      \$19930\ := \$19930%now\;
      \$v5721\ := \$v5721%now\;
      \$19458\ := \$19458%now\;
      \$19185_v\ := \$19185_v%now\;
      \$v5586\ := \$v5586%now\;
      \$18738_next\ := \$18738_next%now\;
      \$19364_v\ := \$19364_v%now\;
      \$v5234\ := \$v5234%now\;
      \$v5760\ := \$v5760%now\;
      \$18974_modulo6684349_result\ := \$18974_modulo6684349_result%now\;
      \$19797_next\ := \$19797_next%now\;
      \$18745_hd\ := \$18745_hd%now\;
      \$18797_branch_if648_result\ := \$18797_branch_if648_result%now\;
      \$19589_copy_root_in_ram6634353_id\ := \$19589_copy_root_in_ram6634353_id%now\;
      \$v5766\ := \$v5766%now\;
      \$19478_v\ := \$19478_v%now\;
      \$19752\ := \$19752%now\;
      \$v4616\ := \$v4616%now\;
      \$19894\ := \$19894%now\;
      \$19819\ := \$19819%now\;
      \$19489\ := \$19489%now\;
      \$v5776\ := \$v5776%now\;
      \$v5019\ := \$v5019%now\;
      \$18807\ := \$18807%now\;
      \$19504\ := \$19504%now\;
      \$18650\ := \$18650%now\;
      \$18837\ := \$18837%now\;
      \$18569\ := \$18569%now\;
      \$19129_modulo6684357_id\ := \$19129_modulo6684357_id%now\;
      \$18805\ := \$18805%now\;
      \$v5869\ := \$v5869%now\;
      \$19112\ := \$19112%now\;
      \$19135_binop_int6434374_arg\ := \$19135_binop_int6434374_arg%now\;
      \$19002_modulo6684356_arg\ := \$19002_modulo6684356_arg%now\;
      \$v5515\ := \$v5515%now\;
      \$19319\ := \$19319%now\;
      \$v5646\ := \$v5646%now\;
      \$v4952\ := \$v4952%now\;
      \$v5610\ := \$v5610%now\;
      \$v5683\ := \$v5683%now\;
      \$18958_binop_int6434364_result\ := \$18958_binop_int6434364_result%now\;
      \$19342\ := \$19342%now\;
      \$19657\ := \$19657%now\;
      \$19777\ := \$19777%now\;
      \$19620\ := \$19620%now\;
      \$18793_make_block579_id\ := \$18793_make_block579_id%now\;
      \$18521_loop666_arg\ := \$18521_loop666_arg%now\;
      \$19803\ := \$19803%now\;
      \$19217\ := \$19217%now\;
      \$v4949\ := \$v4949%now\;
      \$19486\ := \$19486%now\;
      \$v5857\ := \$v5857%now\;
      \$18482\ := \$18482%now\;
      \$v4692\ := \$v4692%now\;
      \$19309_v\ := \$19309_v%now\;
      \$18529\ := \$18529%now\;
      \$19916\ := \$19916%now\;
      \$v5686\ := \$v5686%now\;
      \$v4854\ := \$v4854%now\;
      \$v4628\ := \$v4628%now\;
      \$18703\ := \$18703%now\;
      \$v5506\ := \$v5506%now\;
      \$v4926\ := \$v4926%now\;
      \$19829\ := \$19829%now\;
      \$v4523\ := \$v4523%now\;
      \$v4569\ := \$v4569%now\;
      \$v5749\ := \$v5749%now\;
      \$19209_v\ := \$19209_v%now\;
      \$19482\ := \$19482%now\;
      \$19611\ := \$19611%now\;
      \$19811_copy_root_in_ram6634341_id\ := \$19811_copy_root_in_ram6634341_id%now\;
      \$19784\ := \$19784%now\;
      \$18502\ := \$18502%now\;
      \$v4770\ := \$v4770%now\;
      \$18667_w\ := \$18667_w%now\;
      \$19434\ := \$19434%now\;
      \$19333_compbranch6504388_arg\ := \$19333_compbranch6504388_arg%now\;
      \$19732\ := \$19732%now\;
      \$19609\ := \$19609%now\;
      \$19714_next\ := \$19714_next%now\;
      \$18815\ := \$18815%now\;
      \$v5210\ := \$v5210%now\;
      \$18565\ := \$18565%now\;
      \$v4491\ := \$v4491%now\;
      \$19076_res\ := \$19076_res%now\;
      \$v4727\ := \$v4727%now\;
      \$19015_binop_int6434367_id\ := \$19015_binop_int6434367_id%now\;
      \$18986_modulo6684349_arg\ := \$18986_modulo6684349_arg%now\;
      \$v4734\ := \$v4734%now\;
      \$19656\ := \$19656%now\;
      \$19496_aux664_arg\ := \$19496_aux664_arg%now\;
      \$18480\ := \$18480%now\;
      \$v5537\ := \$v5537%now\;
      \$18458\ := \$18458%now\;
      \$18993_modulo6684349_arg\ := \$18993_modulo6684349_arg%now\;
      \$v5655\ := \$v5655%now\;
      \$19294\ := \$19294%now\;
      \$v5828\ := \$v5828%now\;
      \$19583\ := \$19583%now\;
      \$v5838\ := \$v5838%now\;
      \$19163_forever6704376_id\ := \$19163_forever6704376_id%now\;
      \$18723\ := \$18723%now\;
      \$v4481\ := \$v4481%now\;
      \$v5640\ := \$v5640%now\;
      \$19314\ := \$19314%now\;
      \$18762\ := \$18762%now\;
      \$19034_binop_int6434368_arg\ := \$19034_binop_int6434368_arg%now\;
      \$v4728\ := \$v4728%now\;
      \$v4596\ := \$v4596%now\;
      \$19062_modulo6684349_result\ := \$19062_modulo6684349_result%now\;
      \$18914_modulo6684357_arg\ := \$18914_modulo6684357_arg%now\;
      \$18590\ := \$18590%now\;
      \$19902\ := \$19902%now\;
      \$18670\ := \$18670%now\;
      \$v5604\ := \$v5604%now\;
      \$19248\ := \$19248%now\;
      \$19088_modulo6684349_result\ := \$19088_modulo6684349_result%now\;
      \$19464\ := \$19464%now\;
      \$19072_binop_int6434370_result\ := \$19072_binop_int6434370_result%now\;
      \$v4761\ := \$v4761%now\;
      \$19816\ := \$19816%now\;
      \$19081_modulo6684349_result\ := \$19081_modulo6684349_result%now\;
      \$v4845\ := \$v4845%now\;
      \$v4631\ := \$v4631%now\;
      \$19326_compbranch6504387_arg\ := \$19326_compbranch6504387_arg%now\;
      \$v5035\ := \$v5035%now\;
      \$18685\ := \$18685%now\;
      \$v5603\ := \$v5603%now\;
      \$19628_w\ := \$19628_w%now\;
      \$v5582\ := \$v5582%now\;
      \$18948_modulo6684349_arg\ := \$18948_modulo6684349_arg%now\;
      \$v5060\ := \$v5060%now\;
      \$18668_hd\ := \$18668_hd%now\;
      \$v4552\ := \$v4552%now\;
      \$19187_compare6444358_result\ := \$19187_compare6444358_result%now\;
      \$v5378\ := \$v5378%now\;
      \$19623\ := \$19623%now\;
      \$v5052\ := \$v5052%now\;
      \$v4946\ := \$v4946%now\;
      \$18664\ := \$18664%now\;
      \$18646\ := \$18646%now\;
      \$18852\ := \$18852%now\;
      \$18485\ := \$18485%now\;
      \$19190_binop_compare6454380_result\ := \$19190_binop_compare6454380_result%now\;
      \$19043_modulo6684349_arg\ := \$19043_modulo6684349_arg%now\;
      \$v4936\ := \$v4936%now\;
      \$v4417\ := \$v4417%now\;
      \$18447\ := \$18447%now\;
      \$v4992\ := \$v4992%now\;
      \$v5702\ := \$v5702%now\;
      \$18967_modulo6684349_arg\ := \$18967_modulo6684349_arg%now\;
      \$v5481\ := \$v5481%now\;
      \$18952_modulo6684357_result\ := \$18952_modulo6684357_result%now\;
      \$18662\ := \$18662%now\;
      \$18600\ := \$18600%now\;
      \$v5244\ := \$v5244%now\;
      \$19600\ := \$19600%now\;
      \$19838_copy_root_in_ram6634340_result\ := \$19838_copy_root_in_ram6634340_result%now\;
      \$19885\ := \$19885%now\;
      \$19685\ := \$19685%now\;
      \$19187_compare6444358_id\ := \$19187_compare6444358_id%now\;
      \$18926_modulo6684356_id\ := \$18926_modulo6684356_id%now\;
      \$19720_w\ := \$19720_w%now\;
      \$v5530\ := \$v5530%now\;
      \$18644\ := \$18644%now\;
      \$18466_loop666_id\ := \$18466_loop666_id%now\;
      \$18638_hd\ := \$18638_hd%now\;
      \$v4674\ := \$v4674%now\;
      \$v5250\ := \$v5250%now\;
      \$18563\ := \$18563%now\;
      \$19062_modulo6684349_id\ := \$19062_modulo6684349_id%now\;
      \$18645\ := \$18645%now\;
      \$19897\ := \$19897%now\;
      \$19139_res\ := \$19139_res%now\;
      \$19347_fill6534389_arg\ := \$19347_fill6534389_arg%now\;
      \$19495_loop665_arg\ := \$19495_loop665_arg%now\;
      \$v4695\ := \$v4695%now\;
      \$18576\ := \$18576%now\;
      \$18578\ := \$18578%now\;
      \$18440_make_block579_arg\ := \$18440_make_block579_arg%now\;
      \$19157_forever6704375_id\ := \$19157_forever6704375_id%now\;
      \$19246_v\ := \$19246_v%now\;
      \$19495_loop665_id\ := \$19495_loop665_id%now\;
      \$19515_next\ := \$19515_next%now\;
      \$v4563\ := \$v4563%now\;
      \$v4908\ := \$v4908%now\;
      \$18635\ := \$18635%now\;
      \$19251\ := \$19251%now\;
      \$19648\ := \$19648%now\;
      \$18613_copy_root_in_ram6634346_id\ := \$18613_copy_root_in_ram6634346_id%now\;
      \$19780_loop665_arg\ := \$19780_loop665_arg%now\;
      \$18571_copy_root_in_ram6634345_arg\ := \$18571_copy_root_in_ram6634345_arg%now\;
      \$v5120\ := \$v5120%now\;
      \$19854\ := \$19854%now\;
      \$v4988\ := \$v4988%now\;
      \$v5607\ := \$v5607%now\;
      \$19848\ := \$19848%now\;
      \$19232\ := \$19232%now\;
      \$19814\ := \$19814%now\;
      \$v4680\ := \$v4680%now\;
      \$18906_r\ := \$18906_r%now\;
      \$v5127\ := \$v5127%now\;
      \$18620\ := \$18620%now\;
      \$19887\ := \$19887%now\;
      \$19296_v\ := \$19296_v%now\;
      \$18709\ := \$18709%now\;
      \$v4805\ := \$v4805%now\;
      \$v5514\ := \$v5514%now\;
      \$18913_r\ := \$18913_r%now\;
      \$18457\ := \$18457%now\;
      \$19269\ := \$19269%now\;
      \$19569\ := \$19569%now\;
      \$v5823\ := \$v5823%now\;
      \$v5164\ := \$v5164%now\;
      \$19721_hd\ := \$19721_hd%now\;
      \$v5831\ := \$v5831%now\;
      \$v4740\ := \$v4740%now\;
      \$v5308\ := \$v5308%now\;
      \$v4995\ := \$v4995%now\;
      \$v4601\ := \$v4601%now\;
      \$18484\ := \$18484%now\;
      \$18733\ := \$18733%now\;
      \$v4660\ := \$v4660%now\;
      \$19408_argument3\ := \$19408_argument3%now\;
      \$18828_v\ := \$18828_v%now\;
      \$19390_b\ := \$19390_b%now\;
      \$19727\ := \$19727%now\;
      \$18510\ := \$18510%now\;
      \$19662\ := \$19662%now\;
      \$v5577\ := \$v5577%now\;
      \$19015_binop_int6434367_arg\ := \$19015_binop_int6434367_arg%now\;
      \$19413\ := \$19413%now\;
      \$v4584\ := \$v4584%now\;
      \$19845\ := \$19845%now\;
      \$19337_compare6444359_id\ := \$19337_compare6444359_id%now\;
      \$19698\ := \$19698%now\;
      \$18566\ := \$18566%now\;
      \$18767\ := \$18767%now\;
      \$19359\ := \$19359%now\;
      \$18977_binop_int6434365_arg\ := \$18977_binop_int6434365_arg%now\;
      \$v4878\ := \$v4878%now\;
      \$19267_hd\ := \$19267_hd%now\;
      \$19679\ := \$19679%now\;
      \$v5195\ := \$v5195%now\;
      \$v4433\ := \$v4433%now\;
      \$18864\ := \$18864%now\;
      \$18996_binop_int6434366_arg\ := \$18996_binop_int6434366_arg%now\;
      \$19599\ := \$19599%now\;
      \$19526_forever6704355_arg\ := \$19526_forever6704355_arg%now\;
      \$19578\ := \$19578%now\;
      \$18605\ := \$18605%now\;
      \$19558\ := \$19558%now\;
      \$19280\ := \$19280%now\;
      \$v5278\ := \$v5278%now\;
      \$v5557\ := \$v5557%now\;
      \$19817\ := \$19817%now\;
      \$19238_w6514383_arg\ := \$19238_w6514383_arg%now\;
      \$v5284\ := \$v5284%now\;
      \$v5905\ := \$v5905%now\;
      \$19488\ := \$19488%now\;
      \$19474\ := \$19474%now\;
      \$v5564\ := \$v5564%now\;
      \$18591\ := \$18591%now\;
      \$v4568\ := \$v4568%now\;
      \$v5883\ := \$v5883%now\;
      \$v5555\ := \$v5555%now\;
      \$19726\ := \$19726%now\;
      \$v4842\ := \$v4842%now\;
      \$18834_v\ := \$18834_v%now\;
      \$19401_compbranch6504396_result\ := \$19401_compbranch6504396_result%now\;
      \$18699\ := \$18699%now\;
      \$18680\ := \$18680%now\;
      \$19751\ := \$19751%now\;
      \$19157_forever6704375_arg\ := \$19157_forever6704375_arg%now\;
      \$18584_hd\ := \$18584_hd%now\;
      \$19867\ := \$19867%now\;
      \$v5465\ := \$v5465%now\;
      \$18999_v\ := \$18999_v%now\;
      \$18623\ := \$18623%now\;
      \$19754\ := \$19754%now\;
      \$19825\ := \$19825%now\;
      \$19312_v\ := \$19312_v%now\;
      \$18936_modulo6684349_arg\ := \$18936_modulo6684349_arg%now\;
      \$18460\ := \$18460%now\;
      \$19596\ := \$19596%now\;
      \$18795_offsetclosure_n639_result\ := \$18795_offsetclosure_n639_result%now\;
      \$19918\ := \$19918%now\;
      \$v4328\ := \$v4328%now\;
      \$19373_compbranch6504392_result\ := \$19373_compbranch6504392_result%now\;
      \$v5247\ := \$v5247%now\;
      \$v4543\ := \$v4543%now\;
      \$v5420\ := \$v5420%now\;
      \$19505\ := \$19505%now\;
      \$18570\ := \$18570%now\;
      \$v5263\ := \$v5263%now\;
      \$19391_compare6444359_id\ := \$19391_compare6444359_id%now\;
      \$v5835\ := \$v5835%now\;
      \$18962_res\ := \$18962_res%now\;
      \$18822_v\ := \$18822_v%now\;
      \$v5614\ := \$v5614%now\;
      \$v5027\ := \$v5027%now\;
      \$18610\ := \$18610%now\;
      \$v5069\ := \$v5069%now\;
      \$18684\ := \$18684%now\;
      \$19535_copy_root_in_ram6634354_id\ := \$19535_copy_root_in_ram6634354_id%now\;
      \$v5860\ := \$v5860%now\;
      \$v4414\ := \$v4414%now\;
      \$v5237\ := \$v5237%now\;
      \$19066_modulo6684357_arg\ := \$19066_modulo6684357_arg%now\;
      \$19852\ := \$19852%now\;
      \$18577\ := \$18577%now\;
      \$v5533\ := \$v5533%now\;
      \$18553_forever6704348_arg\ := \$18553_forever6704348_arg%now\;
      \$19387_compbranch6504394_id\ := \$19387_compbranch6504394_id%now\;
      \$18643\ := \$18643%now\;
      \$18754\ := \$18754%now\;
      \$18933_modulo6684357_arg\ := \$18933_modulo6684357_arg%now\;
      \$19397_b\ := \$19397_b%now\;
      \$19279_v\ := \$19279_v%now\;
      \$18933_modulo6684357_result\ := \$18933_modulo6684357_result%now\;
      \$v5485\ := \$v5485%now\;
      \$19550\ := \$19550%now\;
      \$18816\ := \$18816%now\;
      \$19495_loop665_result\ := \$19495_loop665_result%now\;
      \$v5516\ := \$v5516%now\;
      \$v5180\ := \$v5180%now\;
      \$18952_modulo6684357_arg\ := \$18952_modulo6684357_arg%now\;
      \$19855\ := \$19855%now\;
      \$v5426\ := \$v5426%now\;
      \$19313\ := \$19313%now\;
      \$v5542\ := \$v5542%now\;
      \$19565\ := \$19565%now\;
      \$v4863\ := \$v4863%now\;
      \$18980_v\ := \$18980_v%now\;
      \$18521_loop666_id\ := \$18521_loop666_id%now\;
      \$v5870\ := \$v5870%now\;
      \$19800_next\ := \$19800_next%now\;
      \$19746\ := \$19746%now\;
      \$19851_hd\ := \$19851_hd%now\;
      \$18488\ := \$18488%now\;
      \$18746\ := \$18746%now\;
      \$v5203\ := \$v5203%now\;
      \$19222\ := \$19222%now\;
      \$v5290\ := \$v5290%now\;
      \$18796_make_block_n646_id\ := \$18796_make_block_n646_id%now\;
      \$19096_r\ := \$19096_r%now\;
      \$19450_v\ := \$19450_v%now\;
      \$19651\ := \$19651%now\;
      \$v5130\ := \$v5130%now\;
      \$v5595\ := \$v5595%now\;
      \$v4699\ := \$v4699%now\;
      \$18559_copy_root_in_ram6634347_result\ := \$18559_copy_root_in_ram6634347_result%now\;
      \$18831\ := \$18831%now\;
      \$v5123\ := \$v5123%now\;
      \$18829\ := \$18829%now\;
      \$19761\ := \$19761%now\;
      \$19547_copy_root_in_ram6634352_result\ := \$19547_copy_root_in_ram6634352_result%now\;
      \$v5737\ := \$v5737%now\;
      \$19676\ := \$19676%now\;
      \$18450\ := \$18450%now\;
      \$18982_r\ := \$18982_r%now\;
      \$19179_compare6444358_arg\ := \$19179_compare6444358_arg%now\;
      \$v4462\ := \$v4462%now\;
      \$18717\ := \$18717%now\;
      \$v5148\ := \$v5148%now\;
      \$18571_copy_root_in_ram6634345_id\ := \$18571_copy_root_in_ram6634345_id%now\;
      \$v5170\ := \$v5170%now\;
      \$19438\ := \$19438%now\;
      \$19647\ := \$19647%now\;
      \$19483\ := \$19483%now\;
      \$19361_fill6544390_arg\ := \$19361_fill6544390_arg%now\;
      \$19861\ := \$19861%now\;
      \$19211_compare6444358_id\ := \$19211_compare6444358_id%now\;
      \$19786\ := \$19786%now\;
      \$18725\ := \$18725%now\;
      \$18459\ := \$18459%now\;
      \$19135_binop_int6434374_result\ := \$19135_binop_int6434374_result%now\;
      \$v5546\ := \$v5546%now\;
      \$19724\ := \$19724%now\;
      \$18711_w\ := \$18711_w%now\;
      \$18948_modulo6684349_result\ := \$18948_modulo6684349_result%now\;
      \$v5144\ := \$v5144%now\;
      \$19908\ := \$19908%now\;
      \$19858\ := \$19858%now\;
      \$18779\ := \$18779%now\;
      \$v5272\ := \$v5272%now\;
      \$18612\ := \$18612%now\;
      \$19303\ := \$19303%now\;
      \$19551\ := \$19551%now\;
      \$v5269\ := \$v5269%now\;
      \$19186_res\ := \$19186_res%now\;
      \$18689\ := \$18689%now\;
      \$19631\ := \$19631%now\;
      \$18791_loop665_arg\ := \$18791_loop665_arg%now\;
      \$18905_res\ := \$18905_res%now\;
      \$19694\ := \$19694%now\;
      \$18755\ := \$18755%now\;
      \$v5795\ := \$v5795%now\;
      \$v5202\ := \$v5202%now\;
      \$v5565\ := \$v5565%now\;
      \$v4923\ := \$v4923%now\;
      \$19835\ := \$19835%now\;
      \$19588\ := \$19588%now\;
      \$v4943\ := \$v4943%now\;
      \$19078_modulo6684356_id\ := \$19078_modulo6684356_id%now\;
      \$v5317\ := \$v5317%now\;
      result4434 := \result4434%now\;
      \$v5512\ := \$v5512%now\;
      \$18465\ := \$18465%now\;
      \$v4484\ := \$v4484%now\;
      \$18830_v\ := \$18830_v%now\;
      \$19779_loop666_arg\ := \$19779_loop666_arg%now\;
      \$19616\ := \$19616%now\;
      \$v4792\ := \$v4792%now\;
      \$19088_modulo6684349_arg\ := \$19088_modulo6684349_arg%now\;
      \$19666\ := \$19666%now\;
      \$19179_compare6444358_id\ := \$19179_compare6444358_id%now\;
      \$19681_next\ := \$19681_next%now\;
      \$18742\ := \$18742%now\;
      \$18795_offsetclosure_n639_arg\ := \$18795_offsetclosure_n639_arg%now\;
      \$19384_compare6444359_id\ := \$19384_compare6444359_id%now\;
      \$18993_modulo6684349_id\ := \$18993_modulo6684349_id%now\;
      \$19610\ := \$19610%now\;
      \$18856_loop_push6494360_arg\ := \$18856_loop_push6494360_arg%now\;
      \$19909_w\ := \$19909_w%now\;
      \$19686\ := \$19686%now\;
      \$v4975\ := \$v4975%now\;
      \$19019_res\ := \$19019_res%now\;
      \$v5534\ := \$v5534%now\;
      \$18479\ := \$18479%now\;
      \$18525_loop665_result\ := \$18525_loop665_result%now\;
      \$v5893\ := \$v5893%now\;
      \$19671\ := \$19671%now\;
      \$v4475\ := \$v4475%now\;
      \$18734\ := \$18734%now\;
      \$19128_r\ := \$19128_r%now\;
      \$19750\ := \$19750%now\;
      \$19499_aux664_arg\ := \$19499_aux664_arg%now\;
      \$19826\ := \$19826%now\;
      \$18799_w1656_result\ := \$18799_w1656_result%now\;
      \$18798_w652_result\ := \$18798_w652_result%now\;
      \$18467_loop665_arg\ := \$18467_loop665_arg%now\;
      \$19021_modulo6684356_id\ := \$19021_modulo6684356_id%now\;
      \$19088_modulo6684349_id\ := \$19088_modulo6684349_id%now\;
      \$19162\ := \$19162%now\;
      \$v4851\ := \$v4851%now\;
      \$19357_v\ := \$19357_v%now\;
      \$19097_modulo6684356_result\ := \$19097_modulo6684356_result%now\;
      \$v5580\ := \$v5580%now\;
      \$19012_modulo6684349_id\ := \$19012_modulo6684349_id%now\;
      \$18765\ := \$18765%now\;
      \$v4893\ := \$v4893%now\;
      \$v5329\ := \$v5329%now\;
      \$19936\ := \$19936%now\;
      \$19020_r\ := \$19020_r%now\;
      \$19238_w6514383_result\ := \$19238_w6514383_result%now\;
      \$v5601\ := \$v5601%now\;
      \$18996_binop_int6434366_id\ := \$18996_binop_int6434366_id%now\;
      \$v5511\ := \$v5511%now\;
      \$v4570\ := \$v4570%now\;
      \$19675\ := \$19675%now\;
      \$18601\ := \$18601%now\;
      \$v4565\ := \$v4565%now\;
      \$18552\ := \$18552%now\;
      \$19077_r\ := \$19077_r%now\;
      \$v5545\ := \$v5545%now\;
      \$v5031\ := \$v5031%now\;
      \$v5456\ := \$v5456%now\;
      \$v5161\ := \$v5161%now\;
      \$19075_v\ := \$19075_v%now\;
      \$18791_loop665_result\ := \$18791_loop665_result%now\;
      \$18750\ := \$18750%now\;
      \$18718\ := \$18718%now\;
      \$19849\ := \$19849%now\;
      \$19059_modulo6684356_arg\ := \$19059_modulo6684356_arg%now\;
      \$v4724\ := \$v4724%now\;
      \$19423_v\ := \$19423_v%now\;
      \$19352\ := \$19352%now\;
      \$19601_copy_root_in_ram6634352_result\ := \$19601_copy_root_in_ram6634352_result%now\;
      \$18789\ := \$18789%now\;
      \$18977_binop_int6434365_id\ := \$18977_binop_int6434365_id%now\;
      \$v5789\ := \$v5789%now\;
      \$v5450\ := \$v5450%now\;
      \$18681\ := \$18681%now\;
      \$19206_binop_compare6454382_arg\ := \$19206_binop_compare6454382_arg%now\;
      \$v5010\ := \$v5010%now\;
      \$19523\ := \$19523%now\;
      \$18964_modulo6684356_id\ := \$18964_modulo6684356_id%now\;
      \$19923\ := \$19923%now\;
      \$19361_fill6544390_result\ := \$19361_fill6544390_result%now\;
      \$19535_copy_root_in_ram6634354_arg\ := \$19535_copy_root_in_ram6634354_arg%now\;
      \$19564\ := \$19564%now\;
      \$18770\ := \$18770%now\;
      \$19790\ := \$19790%now\;
      \$19509\ := \$19509%now\;
      \$18598_w\ := \$18598_w%now\;
      \$18462\ := \$18462%now\;
      \$19873\ := \$19873%now\;
      \$v5496\ := \$v5496%now\;
      \$v5573\ := \$v5573%now\;
      \$19177_v\ := \$19177_v%now\;
      \$19320_forever6704386_arg\ := \$19320_forever6704386_arg%now\;
      \$19069_modulo6684349_arg\ := \$19069_modulo6684349_arg%now\;
      \$v5225\ := \$v5225%now\;
      \$v5611\ := \$v5611%now\;
      \$v5063\ := \$v5063%now\;
      \$v5393\ := \$v5393%now\;
      \$19778\ := \$19778%now\;
      \$19821\ := \$19821%now\;
      \$v5174\ := \$v5174%now\;
      \$18494\ := \$18494%now\;
      \$19333_compbranch6504388_result\ := \$19333_compbranch6504388_result%now\;
      \$19441_arg\ := \$19441_arg%now\;
      \$18920_binop_int6434362_arg\ := \$18920_binop_int6434362_arg%now\;
      \$v5080\ := \$v5080%now\;
      \$18790_loop666_id\ := \$18790_loop666_id%now\;
      \$v5763\ := \$v5763%now\;
      \$v5618\ := \$v5618%now\;
      \$18613_copy_root_in_ram6634346_result\ := \$18613_copy_root_in_ram6634346_result%now\;
      \$19498_loop665_arg\ := \$19498_loop665_arg%now\;
      \$19467_sp\ := \$19467_sp%now\;
      \$v4799\ := \$v4799%now\;
      \$19187_compare6444358_arg\ := \$19187_compare6444358_arg%now\;
      \$v4860\ := \$v4860%now\;
      \$18849\ := \$18849%now\;
      \$18749\ := \$18749%now\;
      \$18907_modulo6684356_id\ := \$18907_modulo6684356_id%now\;
      \$19794\ := \$19794%now\;
      \$18863\ := \$18863%now\;
      \$19910_hd\ := \$19910_hd%now\;
      \$18958_binop_int6434364_id\ := \$18958_binop_int6434364_id%now\;
      \$v5135\ := \$v5135%now\;
      \$v4495\ := \$v4495%now\;
      \$19320_forever6704386_id\ := \$19320_forever6704386_id%now\;
      \$19300\ := \$19300%now\;
      \$19116_binop_int6434373_arg\ := \$19116_binop_int6434373_arg%now\;
      \$v5147\ := \$v5147%now\;
      \$v4899\ := \$v4899%now\;
      \$19333_compbranch6504388_id\ := \$19333_compbranch6504388_id%now\;
      \$19880_w\ := \$19880_w%now\;
      \$v5730\ := \$v5730%now\;
      \$19366_compbranch6504391_arg\ := \$19366_compbranch6504391_arg%now\;
      \$v5007\ := \$v5007%now\;
      \$19377_compare6444359_result\ := \$19377_compare6444359_result%now\;
      \$19203_compare6444358_result\ := \$19203_compare6444358_result%now\;
      \$v5570\ := \$v5570%now\;
      \$19664\ := \$19664%now\;
      \$19637\ := \$19637%now\;
      \$18926_modulo6684356_result\ := \$18926_modulo6684356_result%now\;
      \$v4431\ := \$v4431%now\;
      \$18854_sp\ := \$18854_sp%now\;
      \$19710\ := \$19710%now\;
      \$19771\ := \$19771%now\;
      \$19057_res\ := \$19057_res%now\;
      \$18907_modulo6684356_arg\ := \$18907_modulo6684356_arg%now\;
      \$18537\ := \$18537%now\;
      \$19785\ := \$19785%now\;
      \$18792_wait662_result\ := \$18792_wait662_result%now\;
      \$18826\ := \$18826%now\;
      \$19307_v\ := \$19307_v%now\;
      \$19354_v\ := \$19354_v%now\;
      \$19463\ := \$19463%now\;
      \$19734\ := \$19734%now\;
      rdy4929 := \rdy4929%now\;
      \$18799_w1656_id\ := \$18799_w1656_id%now\;
      \$19589_copy_root_in_ram6634353_result\ := \$19589_copy_root_in_ram6634353_result%now\;
      \$18472\ := \$18472%now\;
      \$v4666\ := \$v4666%now\;
      \$19129_modulo6684357_arg\ := \$19129_modulo6684357_arg%now\;
      \$v4458\ := \$v4458%now\;
      \$18873_v\ := \$18873_v%now\;
      \$19038_res\ := \$19038_res%now\;
      \$19595\ := \$19595%now\;
      \$19883\ := \$19883%now\;
      \$18677\ := \$18677%now\;
      \$19249\ := \$19249%now\;
      \$v5266\ := \$v5266%now\;
      \$19546\ := \$19546%now\;
      \$v4767\ := \$v4767%now\;
      \$v5189\ := \$v5189%now\;
      \$v4442\ := \$v4442%now\;
      \$19891\ := \$19891%now\;
      \$v5649\ := \$v5649%now\;
      \$v5199\ := \$v5199%now\;
      \$19559_w\ := \$19559_w%now\;
      \$19920\ := \$19920%now\;
      \$v4549\ := \$v4549%now\;
      \$18990_modulo6684357_id\ := \$18990_modulo6684357_id%now\;
      \$19107_modulo6684349_arg\ := \$19107_modulo6684349_arg%now\;
      \$18520\ := \$18520%now\;
      \$19420_w06554397_result\ := \$19420_w06554397_result%now\;
      \$18884_v\ := \$18884_v%now\;
      \$18925_r\ := \$18925_r%now\;
      \$19179_compare6444358_result\ := \$19179_compare6444358_result%now\;
      \$19078_modulo6684356_arg\ := \$19078_modulo6684356_arg%now\;
      \$v5103\ := \$v5103%now\;
      \$19522\ := \$19522%now\;
      \$19544\ := \$19544%now\;
      \$19243\ := \$19243%now\;
      \$19718\ := \$19718%now\;
      \$19148_modulo6684357_arg\ := \$19148_modulo6684357_arg%now\;
      \$19538\ := \$19538%now\;
      \$19255\ := \$19255%now\;
      \$v4571\ := \$v4571%now\;
      \$19275\ := \$19275%now\;
      \$19281\ := \$19281%now\;
      \$18599_hd\ := \$18599_hd%now\;
      \$19836\ := \$19836%now\;
      \$v4872\ := \$v4872%now\;
      \$19043_modulo6684349_id\ := \$19043_modulo6684349_id%now\;
      \$19884\ := \$19884%now\;
      \$19871\ := \$19871%now\;
      \$18851\ := \$18851%now\;
      \$19557\ := \$19557%now\;
      \$19517\ := \$19517%now\;
      \$19532_forever6704350_id\ := \$19532_forever6704350_id%now\;
      \$18782\ := \$18782%now\;
      \$18526_aux664_id\ := \$18526_aux664_id%now\;
      \$v4696\ := \$v4696%now\;
      \$19238_w6514383_id\ := \$19238_w6514383_id%now\;
      \$19582\ := \$19582%now\;
      \$v5344\ := \$v5344%now\;
      \$19570\ := \$19570%now\;
      \$v4619\ := \$v4619%now\;
      \$19888\ := \$19888%now\;
      \$18794_apply638_id\ := \$18794_apply638_id%now\;
      \$19497_loop666_id\ := \$19497_loop666_id%now\;
      \$v4651\ := \$v4651%now\;
      \$18521_loop666_result\ := \$18521_loop666_result%now\;
      \$19901\ := \$19901%now\;
      \$18442_cy\ := \$18442_cy%now\;
      \$19444\ := \$19444%now\;
      \$18549\ := \$18549%now\;
      \$v5468\ := \$v5468%now\;
      \$18604\ := \$18604%now\;
      \$18540\ := \$18540%now\;
      \$18575\ := \$18575%now\;
      \$19330_compare6444359_id\ := \$19330_compare6444359_id%now\;
      \$19085_modulo6684357_arg\ := \$19085_modulo6684357_arg%now\;
      \$19040_modulo6684356_result\ := \$19040_modulo6684356_result%now\;
      \$19324_f0\ := \$19324_f0%now\;
      \$v5083\ := \$v5083%now\;
      \$19540\ := \$19540%now\;
      \$v5817\ := \$v5817%now\;
      \$19554\ := \$19554%now\;
      \$19295\ := \$19295%now\;
      \$19120_res\ := \$19120_res%now\;
      \$18475\ := \$18475%now\;
      \$18580\ := \$18580%now\;
      \$v4612\ := \$v4612%now\;
      \$19005_modulo6684349_arg\ := \$19005_modulo6684349_arg%now\;
      \$v4518\ := \$v4518%now\;
      \$v5637\ := \$v5637%now\;
      \$18848\ := \$18848%now\;
      \$19801\ := \$19801%now\;
      \$18893_v\ := \$18893_v%now\;
      \$19913\ := \$19913%now\;
      \$19262_forever6704385_id\ := \$19262_forever6704385_id%now\;
      \$19210_res\ := \$19210_res%now\;
      \$v5169\ := \$v5169%now\;
      \$18514\ := \$18514%now\;
      \$18747\ := \$18747%now\;
      \$v5402\ := \$v5402%now\;
      \$v5090\ := \$v5090%now\;
      \$v4408\ := \$v4408%now\;
      \$19304\ := \$19304%now\;
      \$v5523\ := \$v5523%now\;
      \$18505\ := \$18505%now\;
      \$18888_next_acc\ := \$18888_next_acc%now\;
      \$19376_b\ := \$19376_b%now\;
      \$18688\ := \$18688%now\;
      \$19100_modulo6684349_arg\ := \$19100_modulo6684349_arg%now\;
      \$19412_sp\ := \$19412_sp%now\;
      \$v4407\ := \$v4407%now\;
      \$v5447\ := \$v5447%now\;
      \$19798\ := \$19798%now\;
      \$v5003\ := \$v5003%now\;
      \$v5873\ := \$v5873%now\;
      \$19097_modulo6684356_arg\ := \$19097_modulo6684356_arg%now\;
      \$v5550\ := \$v5550%now\;
      \$19626\ := \$19626%now\;
      \$19471\ := \$19471%now\;
      \$18721\ := \$18721%now\;
      \$18971_modulo6684357_id\ := \$18971_modulo6684357_id%now\;
      \$18797_branch_if648_id\ := \$18797_branch_if648_id%now\;
      \$v4704\ := \$v4704%now\;
      \$19288_v\ := \$19288_v%now\;
      \$v5390\ := \$v5390%now\;
      \$19366_compbranch6504391_result\ := \$19366_compbranch6504391_result%now\;
      \$v5462\ := \$v5462%now\;
      \$19914\ := \$19914%now\;
      \$v5311\ := \$v5311%now\;
      \$18608\ := \$18608%now\;
      \$19317\ := \$19317%now\;
      \$19141_modulo6684356_result\ := \$19141_modulo6684356_result%now\;
      \$18511\ := \$18511%now\;
      \$v4671\ := \$v4671%now\;
      \$19487\ := \$19487%now\;
      \$18522_loop665_arg\ := \$18522_loop665_arg%now\;
      \$v4420\ := \$v4420%now\;
      \$19625\ := \$19625%now\;
      \$v5576\ := \$v5576%now\;
      \$19886\ := \$19886%now\;
      \$v5482\ := \$v5482%now\;
      result4928 := \result4928%now\;
      \$19773\ := \$19773%now\;
      \$v4424\ := \$v4424%now\;
      \$19787\ := \$19787%now\;
      \$19104_modulo6684357_result\ := \$19104_modulo6684357_result%now\;
      \$v5769\ := \$v5769%now\;
      \$19496_aux664_result\ := \$19496_aux664_result%now\;
      \$19717\ := \$19717%now\;
      \$18647\ := \$18647%now\;
      \$19155\ := \$19155%now\;
      \$18661\ := \$18661%now\;
      \$v4587\ := \$v4587%now\;
      \$19939\ := \$19939%now\;
      \$18832_v\ := \$18832_v%now\;
      \$19227\ := \$19227%now\;
      \$19650\ := \$19650%now\;
      \$18495\ := \$18495%now\;
      \$18551\ := \$18551%now\;
      \$v5658\ := \$v5658%now\;
      \$19276\ := \$19276%now\;
      \$19859\ := \$19859%now\;
      \$19325\ := \$19325%now\;
      \$18977_binop_int6434365_result\ := \$18977_binop_int6434365_result%now\;
      \$18944_r\ := \$18944_r%now\;
      \$18527\ := \$18527%now\;
      \$19119_v\ := \$19119_v%now\;
      \$18648\ := \$18648%now\;
      \$19793\ := \$19793%now\;
      \$18877_v\ := \$18877_v%now\;
      \$18939_binop_int6434363_id\ := \$18939_binop_int6434363_id%now\;
      \$v5673\ := \$v5673%now\;
      \$19190_binop_compare6454380_id\ := \$19190_binop_compare6454380_id%now\;
      \$19842\ := \$19842%now\;
      \$19144_modulo6684349_id\ := \$19144_modulo6684349_id%now\;
      \$v5536\ := \$v5536%now\;
      \$v5299\ := \$v5299%now\;
      \$19601_copy_root_in_ram6634352_arg\ := \$19601_copy_root_in_ram6634352_arg%now\;
      \$18539\ := \$18539%now\;
      \$18936_modulo6684349_id\ := \$18936_modulo6684349_id%now\;
      \$19015_binop_int6434367_result\ := \$19015_binop_int6434367_result%now\;
      \$19171_compare6444358_id\ := \$19171_compare6444358_id%now\;
      \$19597\ := \$19597%now\;
      \$19581\ := \$19581%now\;
      \$v4338\ := \$v4338%now\;
      \$19384_compare6444359_result\ := \$19384_compare6444359_result%now\;
      \$19748\ := \$19748%now\;
      \$18522_loop665_id\ := \$18522_loop665_id%now\;
      \$18461\ := \$18461%now\;
      \$19256_v\ := \$19256_v%now\;
      \$v5206\ := \$v5206%now\;
      \$18824_v\ := \$18824_v%now\;
      \$v5059\ := \$v5059%now\;
      \$18657\ := \$18657%now\;
      \$v5026\ := \$v5026%now\;
      \$v4996\ := \$v4996%now\;
      \$v5036\ := \$v5036%now\;
      \$18825\ := \$18825%now\;
      \$18806\ := \$18806%now\;
      \$v4866\ := \$v4866%now\;
      \$v4647\ := \$v4647%now\;
      \$18891\ := \$18891%now\;
      \$18843\ := \$18843%now\;
      \$v4330\ := \$v4330%now\;
      \$19370_compare6444359_id\ := \$19370_compare6444359_id%now\;
      \$19601_copy_root_in_ram6634352_id\ := \$19601_copy_root_in_ram6634352_id%now\;
      \$v5281\ := \$v5281%now\;
      \$v4546\ := \$v4546%now\;
      \$v4779\ := \$v4779%now\;
      \$v4636\ := \$v4636%now\;
      \$v4812\ := \$v4812%now\;
      \$v5574\ := \$v5574%now\;
      \$18526_aux664_arg\ := \$18526_aux664_arg%now\;
      \$19308_v\ := \$19308_v%now\;
      \$18793_make_block579_arg\ := \$18793_make_block579_arg%now\;
      \$18437_loop666_arg\ := \$18437_loop666_arg%now\;
      \$19206_binop_compare6454382_result\ := \$19206_binop_compare6454382_result%now\;
      \$18444\ := \$18444%now\;
      \$19066_modulo6684357_id\ := \$19066_modulo6684357_id%now\;
      \$19046_r\ := \$19046_r%now\;
      \$19837\ := \$19837%now\;
      \$v5429\ := \$v5429%now\;
      \$19571\ := \$19571%now\;
      \$v4978\ := \$v4978%now\;
      \$v4920\ := \$v4920%now\;
      \$v5799\ := \$v5799%now\;
      \$18524_loop666_arg\ := \$18524_loop666_arg%now\;
      \$18810\ := \$18810%now\;
      \$19944\ := \$19944%now\;
      \$18880\ := \$18880%now\;
      \$18869\ := \$18869%now\;
      \$v5490\ := \$v5490%now\;
      \$18659\ := \$18659%now\;
      \$v5257\ := \$v5257%now\;
      \$18945_modulo6684356_id\ := \$18945_modulo6684356_id%now\;
      \$18683_hd\ := \$18683_hd%now\;
      \$v4428\ := \$v4428%now\;
      \$v5055\ := \$v5055%now\;
      \$19774\ := \$19774%now\;
      \$v5522\ := \$v5522%now\;
      \$19783\ := \$19783%now\;
      \$19125_modulo6684349_result\ := \$19125_modulo6684349_result%now\;
      \$19097_modulo6684356_id\ := \$19097_modulo6684356_id%now\;
      \$19507_next\ := \$19507_next%now\;
      rdy4400 := \rdy4400%now\;
      \$19542\ := \$19542%now\;
      \$v5042\ := \$v5042%now\;
      \$18813\ := \$18813%now\;
      \$19220\ := \$19220%now\;
      \$v4667\ := \$v4667%now\;
      \$v4678\ := \$v4678%now\;
      \$19211_compare6444358_result\ := \$19211_compare6444358_result%now\;
      \$18790_loop666_result\ := \$18790_loop666_result%now\;
      \$19804\ := \$19804%now\;
      \$18622\ := \$18622%now\;
      \$v4519\ := \$v4519%now\;
      \$19667\ := \$19667%now\;
      \$v4593\ := \$v4593%now\;
      \$19811_copy_root_in_ram6634341_arg\ := \$19811_copy_root_in_ram6634341_arg%now\;
      \$18695\ := \$18695%now\;
      \$19789_next\ := \$19789_next%now\;
      \$19259\ := \$19259%now\;
      \$18437_loop666_id\ := \$18437_loop666_id%now\;
      \$19203_compare6444358_id\ := \$19203_compare6444358_id%now\;
      \$19788\ := \$19788%now\;
      \$19141_modulo6684356_arg\ := \$19141_modulo6684356_arg%now\;
      \$18473\ := \$18473%now\;
      \$v5134\ := \$v5134%now\;
      \$19144_modulo6684349_result\ := \$19144_modulo6684349_result%now\;
      \$19932\ := \$19932%now\;
      \$18603\ := \$18603%now\;
      \$v5365\ := \$v5365%now\;
      \$19701\ := \$19701%now\;
      \$19543\ := \$19543%now\;
      \$v5168\ := \$v5168%now\;
      \$v4529\ := \$v4529%now\;
      \$v4839\ := \$v4839%now\;
      \$v4679\ := \$v4679%now\;
      \$19796\ := \$19796%now\;
      \$18845\ := \$18845%now\;
      \$v5233\ := \$v5233%now\;
      \$18438_loop665_arg\ := \$18438_loop665_arg%now\;
      \$19337_compare6444359_arg\ := \$19337_compare6444359_arg%now\;
      \$v4632\ := \$v4632%now\;
      \$v4957\ := \$v4957%now\;
      \$19336_b\ := \$19336_b%now\;
      \$19709\ := \$19709%now\;
      \$19031_modulo6684349_result\ := \$19031_modulo6684349_result%now\;
      \$19824_hd\ := \$19824_hd%now\;
      \$19619\ := \$19619%now\;
      \$18546\ := \$18546%now\;
      \$v5872\ := \$v5872%now\;
      \$19818\ := \$19818%now\;
      \$18971_modulo6684357_arg\ := \$18971_modulo6684357_arg%now\;
      \$v4502\ := \$v4502%now\;
      \$19326_compbranch6504387_id\ := \$19326_compbranch6504387_id%now\;
      \$18531\ := \$18531%now\;
      \$v4802\ := \$v4802%now\;
      \$18841\ := \$18841%now\;
      \$v4639\ := \$v4639%now\;
      \$19466_sp\ := \$19466_sp%now\;
      \$18567\ := \$18567%now\;
      \$v4683\ := \$v4683%now\;
      \$19643_w\ := \$19643_w%now\;
      \$18649\ := \$18649%now\;
      \$18929_modulo6684349_arg\ := \$18929_modulo6684349_arg%now\;
      \$v5184\ := \$v5184%now\;
      \$v4335\ := \$v4335%now\;
      \$v5915\ := \$v5915%now\;
      \$19169_v\ := \$19169_v%now\;
      \$v5487\ := \$v5487%now\;
      \$v5552\ := \$v5552%now\;
      \$19361_fill6544390_id\ := \$19361_fill6544390_id%now\;
      \$v5811\ := \$v5811%now\;
      \$19512\ := \$19512%now\;
      \$v4471\ := \$v4471%now\;
      \$19725\ := \$19725%now\;
      \$19844\ := \$19844%now\;
      \$18732\ := \$18732%now\;
      \$18618\ := \$18618%now\;
      \$19387_compbranch6504394_arg\ := \$19387_compbranch6504394_arg%now\;
      \$19027_r\ := \$19027_r%now\;
      \$v5471\ := \$v5471%now\;
      \$19659_hd\ := \$19659_hd%now\;
      \$19875\ := \$19875%now\;
      \$19639\ := \$19639%now\;
      \$18470\ := \$18470%now\;
      \$19310\ := \$19310%now\;
      \$19815\ := \$19815%now\;
      \$v5696\ := \$v5696%now\;
      \$19350_v\ := \$19350_v%now\;
      \$19503\ := \$19503%now\;
      \$19182_binop_compare6454379_result\ := \$19182_binop_compare6454379_result%now\;
      \$18955_modulo6684349_result\ := \$18955_modulo6684349_result%now\;
      \$18476\ := \$18476%now\;
      \$18443\ := \$18443%now\;
      \$19230_v\ := \$19230_v%now\;
      \$19018_v\ := \$19018_v%now\;
      \$19713\ := \$19713%now\;
      \$19218_v\ := \$19218_v%now\;
      \$19009_modulo6684357_arg\ := \$19009_modulo6684357_arg%now\;
      \$19498_loop665_result\ := \$19498_loop665_result%now\;
      \$v5198\ := \$v5198%now\;
      \$19741\ := \$19741%now\;
      \$v4581\ := \$v4581%now\;
      \$19161\ := \$19161%now\;
      \$19156\ := \$19156%now\;
      \$19104_modulo6684357_arg\ := \$19104_modulo6684357_arg%now\;
      \$18492\ := \$18492%now\;
      \$v5571\ := \$v5571%now\;
      \$v4615\ := \$v4615%now\;
      \$19937\ := \$19937%now\;
      \$18917_modulo6684349_arg\ := \$18917_modulo6684349_arg%now\;
      \$v5384\ := \$v5384%now\;
      \$18939_binop_int6434363_arg\ := \$18939_binop_int6434363_arg%now\;
      \$19572\ := \$19572%now\;
      \$18898\ := \$18898%now\;
      \$19391_compare6444359_result\ := \$19391_compare6444359_result%now\;
      \$v5563\ := \$v5563%now\;
      \$18948_modulo6684349_id\ := \$18948_modulo6684349_id%now\;
      \$v5897\ := \$v5897%now\;
      \$19100_modulo6684349_id\ := \$19100_modulo6684349_id%now\;
      \$19409_sp\ := \$19409_sp%now\;
      \$18478\ := \$18478%now\;
      \$19047_modulo6684357_result\ := \$19047_modulo6684357_result%now\;
      \$19009_modulo6684357_result\ := \$19009_modulo6684357_result%now\;
      \$v5072\ := \$v5072%now\;
      \$18895_v\ := \$18895_v%now\;
      \$18559_copy_root_in_ram6634347_id\ := \$18559_copy_root_in_ram6634347_id%now\;
      \$18559_copy_root_in_ram6634347_arg\ := \$18559_copy_root_in_ram6634347_arg%now\;
      \$19922\ := \$19922%now\;
      \$19125_modulo6684349_id\ := \$19125_modulo6684349_id%now\;
      \$18629\ := \$18629%now\;
      \$v4887\ := \$v4887%now\;
      \$v4556\ := \$v4556%now\;
      \$v5453\ := \$v5453%now\;
      \$19731\ := \$19731%now\;
      \$19449\ := \$19449%now\;
      \$18669\ := \$18669%now\;
      \$18660\ := \$18660%now\;
      rdy4573 := \rdy4573%now\;
      \$18795_offsetclosure_n639_id\ := \$18795_offsetclosure_n639_id%now\;
      \$19401_compbranch6504396_arg\ := \$19401_compbranch6504396_arg%now\;
      \$19878\ := \$19878%now\;
      \$v5066\ := \$v5066%now\;
      \$18631\ := \$18631%now\;
      \$v4327\ := \$v4327%now\;
      \$19234_sp\ := \$19234_sp%now\;
      \$18687\ := \$18687%now\;
      \$19811_copy_root_in_ram6634341_result\ := \$19811_copy_root_in_ram6634341_result%now\;
      rdy4608 := \rdy4608%now\;
      \$19728\ := \$19728%now\;
      \$v5492\ := \$v5492%now\;
      \$19843\ := \$19843%now\;
      \$19532_forever6704350_arg\ := \$19532_forever6704350_arg%now\;
      \$19028_modulo6684357_id\ := \$19028_modulo6684357_id%now\;
      \$18958_binop_int6434364_arg\ := \$18958_binop_int6434364_arg%now\;
      \$v4700\ := \$v4700%now\;
      \$19301_v\ := \$19301_v%now\;
      \$v4940\ := \$v4940%now\;
      \$19012_modulo6684349_result\ := \$19012_modulo6684349_result%now\;
      \$19268\ := \$19268%now\;
      \$19772\ := \$19772%now\;
      \$19226\ := \$19226%now\;
      \$v5727\ := \$v5727%now\;
      \$18889_v\ := \$18889_v%now\;
      \$19882\ := \$19882%now\;
      \$19877\ := \$19877%now\;
      \$19091_binop_int6434371_id\ := \$19091_binop_int6434371_id%now\;
      \$v4796\ := \$v4796%now\;
      \$18907_modulo6684356_result\ := \$18907_modulo6684356_result%now\;
      \$19561\ := \$19561%now\;
      \$19282_v\ := \$19282_v%now\;
      \$19806\ := \$19806%now\;
      \$19257_v\ := \$19257_v%now\;
      \$19660\ := \$19660%now\;
      \$18583_w\ := \$18583_w%now\;
      \$v4818\ := \$v4818%now\;
      \$v4750\ := \$v4750%now\;
      \$19492\ := \$19492%now\;
      \$18525_loop665_id\ := \$18525_loop665_id%now\;
      \$19311\ := \$19311%now\;
      \$19743\ := \$19743%now\;
      \$v4775\ := \$v4775%now\;
      \$v4713\ := \$v4713%now\;
      \$19519\ := \$19519%now\;
      \$19870\ := \$19870%now\;
      \$v4540\ := \$v4540%now\;
      \$19638\ := \$19638%now\;
      \$v4821\ := \$v4821%now\;
      \$v5664\ := \$v5664%now\;
      \$19211_compare6444358_arg\ := \$19211_compare6444358_arg%now\;
      \$18500\ := \$18500%now\;
      \$18545_next\ := \$18545_next%now\;
      \$19078_modulo6684356_result\ := \$19078_modulo6684356_result%now\;
      \$19868\ := \$19868%now\;
      \$19047_modulo6684357_id\ := \$19047_modulo6684357_id%now\;
      \$18663\ := \$18663%now\;
      \$18679\ := \$18679%now\;
      \$19053_binop_int6434369_result\ := \$19053_binop_int6434369_result%now\;
      \$v4937\ := \$v4937%now\;
      \$v5305\ := \$v5305%now\;
      \$18986_modulo6684349_result\ := \$18986_modulo6684349_result%now\;
      \$19266\ := \$19266%now\;
      \$19447_sp\ := \$19447_sp%now\;
      \$19084_r\ := \$19084_r%now\;
      \$19779_loop666_result\ := \$19779_loop666_result%now\;
      \$v5825\ := \$v5825%now\;
      \$18464_rdy\ := \$18464_rdy%now\;
      \$19636\ := \$19636%now\;
      \$19329_b\ := \$19329_b%now\;
      \$v5596\ := \$v5596%now\;
      \$19031_modulo6684349_id\ := \$19031_modulo6684349_id%now\;
      \$19526_forever6704355_id\ := \$19526_forever6704355_id%now\;
      \$19926\ := \$19926%now\;
      \$19614_hd\ := \$19614_hd%now\;
      \$19594\ := \$19594%now\;
      \$18542_next\ := \$18542_next%now\;
      \$18553_forever6704348_id\ := \$18553_forever6704348_id%now\;
      \$19521\ := \$19521%now\;
      \$19832\ := \$19832%now\;
      \$v4455\ := \$v4455%now\;
      \$v4640\ := \$v4640%now\;
      \$19053_binop_int6434369_arg\ := \$19053_binop_int6434369_arg%now\;
      \$18508\ := \$18508%now\;
      \$19684\ := \$19684%now\;
      \$19315\ := \$19315%now\;
      \$19166_binop_compare6454377_id\ := \$19166_binop_compare6454377_id%now\;
      \$19110\ := \$19110%now\;
      \$19678\ := \$19678%now\;
      \$v5405\ := \$v5405%now\;
      \$v5622\ := \$v5622%now\;
      \$v5188\ := \$v5188%now\;
      \$v5138\ := \$v5138%now\;
      \$19198_binop_compare6454381_result\ := \$19198_binop_compare6454381_result%now\;
      \$v4972\ := \$v4972%now\;
      \$19872\ := \$19872%now\;
      \$19031_modulo6684349_arg\ := \$19031_modulo6684349_arg%now\;
      \$19405_compare6444359_arg\ := \$19405_compare6444359_arg%now\;
      \$v4754\ := \$v4754%now\;
      \$v5254\ := \$v5254%now\;
      \$v5275\ := \$v5275%now\;
      \$18642\ := \$18642%now\;
      \$19892\ := \$19892%now\;
      \$v4339\ := \$v4339%now\;
      \$v4532\ := \$v4532%now\;
      \$v5260\ := \$v5260%now\;
      \$19021_modulo6684356_arg\ := \$19021_modulo6684356_arg%now\;
      \$18996_binop_int6434366_result\ := \$18996_binop_int6434366_result%now\;
      \$19005_modulo6684349_id\ := \$19005_modulo6684349_id%now\;
      \$18522_loop665_result\ := \$18522_loop665_result%now\;
      \$18682_w\ := \$18682_w%now\;
      \$18914_modulo6684357_id\ := \$18914_modulo6684357_id%now\;
      \$18673\ := \$18673%now\;
      \$19766\ := \$19766%now\;
      \$v4558\ := \$v4558%now\;
      \$19214\ := \$19214%now\;
      \$19566\ := \$19566%now\;
      \$v4337\ := \$v4337%now\;
      \$v5096\ := \$v5096%now\;
      \$v5359\ := \$v5359%now\;
      \$19174_binop_compare6454378_result\ := \$19174_binop_compare6454378_result%now\;
      \$19563\ := \$19563%now\;
      \$v4606\ := \$v4606%now\;
      \$v5141\ := \$v5141%now\;
      \$18639\ := \$18639%now\;
      \$19154\ := \$19154%now\;
      \$18562\ := \$18562%now\;
      \$v4449\ := \$v4449%now\;
      \$v4605\ := \$v4605%now\;
      \$v4539\ := \$v4539%now\;
      \$18666\ := \$18666%now\;
      \$19781_aux664_id\ := \$19781_aux664_id%now\;
      \$18904_v\ := \$18904_v%now\;
      \$18498\ := \$18498%now\;
      \$v4562\ := \$v4562%now\;
      \$19497_loop666_arg\ := \$19497_loop666_arg%now\;
      \$18564\ := \$18564%now\;
      \$v5335\ := \$v5335%now\;
      \$19834\ := \$19834%now\;
      \$19700\ := \$19700%now\;
      \$19769\ := \$19769%now\;
      \$19907\ := \$19907%now\;
      \$18724\ := \$18724%now\;
      \$19425\ := \$19425%now\;
      \$19293\ := \$19293%now\;
      \$19147_r\ := \$19147_r%now\;
      \$19950\ := \$19950%now\;
      \$19355\ := \$19355%now\;
      \$19024_modulo6684349_id\ := \$19024_modulo6684349_id%now\;
      \$19665\ := \$19665%now\;
      \$19351\ := \$19351%now\;
      \$19500\ := \$19500%now\;
      \$v4833\ := \$v4833%now\;
      \$v4791\ := \$v4791%now\;
      \$v4746\ := \$v4746%now\;
      \$v5524\ := \$v5524%now\;
      \$19856\ := \$19856%now\;
      \$18456\ := \$18456%now\;
      \$19021_modulo6684356_result\ := \$19021_modulo6684356_result%now\;
      \$v5560\ := \$v5560%now\;
      \$v4751\ := \$v4751%now\;
      \$18487\ := \$18487%now\;
      \$19755\ := \$19755%now\;
      \$19233\ := \$19233%now\;
      \$18654\ := \$18654%now\;
      \$v4911\ := \$v4911%now\;
      \$v5743\ := \$v5743%now\;
      \$19414\ := \$19414%now\;
      \$19649\ := \$19649%now\;
      \$18702\ := \$18702%now\;
      \$18897\ := \$18897%now\;
      \$v4496\ := \$v4496%now\;
      \$18967_modulo6684349_result\ := \$18967_modulo6684349_result%now\;
      \$v5477\ := \$v5477%now\;
      \$v4675\ := \$v4675%now\;
      \$v5107\ := \$v5107%now\;
      \$19485\ := \$19485%now\;
      \$v5597\ := \$v5597%now\;
      \$19132_modulo6684349_arg\ := \$19132_modulo6684349_arg%now\;
      \$18781\ := \$18781%now\;
      \$19252_forever6704384_id\ := \$19252_forever6704384_id%now\;
      \$v4984\ := \$v4984%now\;
      \$v5753\ := \$v5753%now\;
      \$18896_v\ := \$18896_v%now\;
      \$18737\ := \$18737%now\;
      \$18439_wait662_result\ := \$18439_wait662_result%now\;
      \$v5102\ := \$v5102%now\;
      \$v4813\ := \$v4813%now\;
      \$v5432\ := \$v5432%now\;
      \$19642\ := \$19642%now\;
      \$18446_dur\ := \$18446_dur%now\;
      \$18625_copy_root_in_ram6634345_id\ := \$18625_copy_root_in_ram6634345_id%now\;
      \$v5314\ := \$v5314%now\;
      \$v5540\ := \$v5540%now\;
      \$19617\ := \$19617%now\;
      \$19451\ := \$19451%now\;
      \$18556_forever6704344_id\ := \$18556_forever6704344_id%now\;
      \$19585\ := \$19585%now\;
      \$18886\ := \$18886%now\;
      \$18439_wait662_id\ := \$18439_wait662_id%now\;
      \$v5441\ := \$v5441%now\;
      \$19737\ := \$19737%now\;
      \$19879\ := \$19879%now\;
      \$19072_binop_int6434370_id\ := \$19072_binop_int6434370_id%now\;
      \$19462\ := \$19462%now\;
      \$18516\ := \$18516%now\;
      \$18838_v\ := \$18838_v%now\;
      \$v5502\ := \$v5502%now\;
      \$v5814\ := \$v5814%now\;
      \$v5845\ := \$v5845%now\;
      \$18438_loop665_result\ := \$18438_loop665_result%now\;
      \$19658_w\ := \$19658_w%now\;
      \$19182_binop_compare6454379_arg\ := \$19182_binop_compare6454379_arg%now\;
      \$18901_binop_int6434361_result\ := \$18901_binop_int6434361_result%now\;
      \$18453\ := \$18453%now\;
      \$19260\ := \$19260%now\;
      \$v5605\ := \$v5605%now\;
      \$18971_modulo6684357_result\ := \$18971_modulo6684357_result%now\;
      \$19853\ := \$19853%now\;
      \$v5131\ := \$v5131%now\;
      \$18820_v\ := \$18820_v%now\;
      \$18571_copy_root_in_ram6634345_result\ := \$18571_copy_root_in_ram6634345_result%now\;
      \$18515\ := \$18515%now\;
      \$v4689\ := \$v4689%now\;
      \$18914_modulo6684357_result\ := \$18914_modulo6684357_result%now\;
      \$v5497\ := \$v5497%now\;
      \$19951\ := \$19951%now\;
      \$19807\ := \$19807%now\;
      \$19241_v\ := \$19241_v%now\;
      \$19242\ := \$19242%now\;
      \$19539\ := \$19539%now\;
      \$18752\ := \$18752%now\;
      \$v5544\ := \$v5544%now\;
      result4607 := \result4607%now\;
      \$19091_binop_int6434371_arg\ := \$19091_binop_int6434371_arg%now\;
      \$19345\ := \$19345%now\;
      \$v5491\ := \$v5491%now\;
      \$18844\ := \$18844%now\;
      \$18963_r\ := \$18963_r%now\;
      \$v5652\ := \$v5652%now\;
      \$v5876\ := \$v5876%now\;
      \$19113_forever6704372_id\ := \$19113_forever6704372_id%now\;
      \$19383_b\ := \$19383_b%now\;
      \$19584\ := \$19584%now\;
      \$19942\ := \$19942%now\;
      \$19615\ := \$19615%now\;
      \$18676\ := \$18676%now\;
      \$v4514\ := \$v4514%now\;
      \$19316\ := \$19316%now\;
      \$19148_modulo6684357_id\ := \$19148_modulo6684357_id%now\;
      \$v4492\ := \$v4492%now\;
      \$v5347\ := \$v5347%now\;
      \$v5411\ := \$v5411%now\;
      \$18756\ := \$18756%now\;
      \$19865_w\ := \$19865_w%now\;
      \$18533\ := \$18533%now\;
      \$19297_v\ := \$19297_v%now\;
      \$18497\ := \$18497%now\;
      \$19062_modulo6684349_arg\ := \$19062_modulo6684349_arg%now\;
      \$19456\ := \$19456%now\;
      \$v5909\ := \$v5909%now\;
      \$v5356\ := \$v5356%now\;
      \$v5584\ := \$v5584%now\;
      \$v5023\ := \$v5023%now\;
      \$18766\ := \$18766%now\;
      \$19770\ := \$19770%now\;
      \$v4960\ := \$v4960%now\;
      \$18674\ := \$18674%now\;
      \$18595\ := \$18595%now\;
      \$19927\ := \$19927%now\;
      \$v5293\ := \$v5293%now\;
      \$v5525\ := \$v5525%now\;
      \$18786\ := \$18786%now\;
      \$19592\ := \$19592%now\;
      \$18748\ := \$18748%now\;
      \$18448_dis\ := \$18448_dis%now\;
      \$19398_compare6444359_result\ := \$19398_compare6444359_result%now\;
      \$19202_res\ := \$19202_res%now\;
      \$18951_r\ := \$18951_r%now\;
      \$19040_modulo6684356_arg\ := \$19040_modulo6684356_arg%now\;
      \$v5724\ := \$v5724%now\;
      \$18780\ := \$18780%now\;
      \$18651\ := \$18651%now\;
      \$19518_next\ := \$19518_next%now\;
      \$19005_modulo6684349_result\ := \$19005_modulo6684349_result%now\;
      \$18808\ := \$18808%now\;
      \$18715\ := \$18715%now\;
      \$19799\ := \$19799%now\;
      \$v5505\ := \$v5505%now\;
      \$v5867\ := \$v5867%now\;
      \$19646\ := \$19646%now\;
      \$19833\ := \$19833%now\;
      \$19182_binop_compare6454379_id\ := \$19182_binop_compare6454379_id%now\;
      \$v5000\ := \$v5000%now\;
      \$v5185\ := \$v5185%now\;
      \$v5034\ := \$v5034%now\;
      \$18467_loop665_result\ := \$18467_loop665_result%now\;
      \$v5222\ := \$v5222%now\;
      \$v4782\ := \$v4782%now\;
      \$19547_copy_root_in_ram6634352_id\ := \$19547_copy_root_in_ram6634352_id%now\;
      \$19915\ := \$19915%now\;
      \$19719\ := \$19719%now\;
      \$18777\ := \$18777%now\;
      \$18550\ := \$18550%now\;
      \$18842\ := \$18842%now\;
      \$18489\ := \$18489%now\;
      \$18439_wait662_arg\ := \$18439_wait662_arg%now\;
      \$19100_modulo6684349_result\ := \$19100_modulo6684349_result%now\;
      \$19135_binop_int6434374_id\ := \$19135_binop_int6434374_id%now\;
      \$18796_make_block_n646_arg\ := \$18796_make_block_n646_arg%now\;
      \$v5084\ := \$v5084%now\;
      \$v4654\ := \$v4654%now\;
      \$19820\ := \$19820%now\;
      \$18901_binop_int6434361_arg\ := \$18901_binop_int6434361_arg%now\;
      \$18701\ := \$18701%now\;
      \$18768_w\ := \$18768_w%now\;
      \$19586\ := \$19586%now\;
      \$v5709\ := \$v5709%now\;
      \$18613_copy_root_in_ram6634346_arg\ := \$18613_copy_root_in_ram6634346_arg%now\;
      \$19917\ := \$19917%now\;
      \$19138_v\ := \$19138_v%now\;
      \$19697\ := \$19697%now\;
      \$v4423\ := \$v4423%now\;
      result4963 := \result4963%now\;
      \$18794_apply638_arg\ := \$18794_apply638_arg%now\;
      \$18792_wait662_arg\ := \$18792_wait662_arg%now\;
      \$18741\ := \$18741%now\;
      \$18735\ := \$18735%now\;
      \$v5039\ := \$v5039%now\;
      \$19677\ := \$19677%now\;
      \$v5296\ := \$v5296%now\;
      \$18714\ := \$18714%now\;
      \$19231\ := \$19231%now\;
      \$v5689\ := \$v5689%now\;
      \$v5251\ := \$v5251%now\;
      \$19876\ := \$19876%now\;
      \$v5606\ := \$v5606%now\;
      \$v5670\ := \$v5670%now\;
      \$18794_apply638_result\ := \$18794_apply638_result%now\;
      \$19921\ := \$19921%now\;
      \$19420_w06554397_id\ := \$19420_w06554397_id%now\;
      \$v4719\ := \$v4719%now\;
      \$19059_modulo6684356_id\ := \$19059_modulo6684356_id%now\;
      \$19864\ := \$19864%now\;
      \$19347_fill6534389_result\ := \$19347_fill6534389_result%now\;
      \$v5099\ := \$v5099%now\;
      \$19860\ := \$19860%now\;
      \$19781_aux664_arg\ := \$19781_aux664_arg%now\;
      \$v4827\ := \$v4827%now\;
      \$18964_modulo6684356_arg\ := \$18964_modulo6684356_arg%now\;
      \$v5802\ := \$v5802%now\;
      \$v4917\ := \$v4917%now\;
      \$19302\ := \$19302%now\;
      \$v5368\ := \$v5368%now\;
      \$19823_w\ := \$19823_w%now\;
      \$v5494\ := \$v5494%now\;
      \$19668\ := \$19668%now\;
      \$19398_compare6444359_id\ := \$19398_compare6444359_id%now\;
      \$18574\ := \$18574%now\;
      \$19228_v\ := \$19228_v%now\;
      \$v5079\ := \$v5079%now\;
      \$19749\ := \$19749%now\;
      \$19795\ := \$19795%now\;
      \$19203_compare6444358_arg\ := \$19203_compare6444358_arg%now\;
      \$19768\ := \$19768%now\;
      \$v4809\ := \$v4809%now\;
      \$19941\ := \$19941%now\;
      \$v4902\ := \$v4902%now\;
      \$18899\ := \$18899%now\;
      \$19605\ := \$19605%now\;
      \$19514\ := \$19514%now\;
      \$v4836\ := \$v4836%now\;
      \$18640\ := \$18640%now\;
      \$v4716\ := \$v4716%now\;
      \$v5396\ := \$v5396%now\;
      \$19341\ := \$19341%now\;
      \$18870_v\ := \$18870_v%now\;
      \$19722\ := \$19722%now\;
      \$19475\ := \$19475%now\;
      \$v5353\ := \$v5353%now\;
      \$v4953\ := \$v4953%now\;
      \$19460\ := \$19460%now\;
      \$19470\ := \$19470%now\;
      \$19580\ := \$19580%now\;
      \$19893\ := \$19893%now\;
      \$v4597\ := \$v4597%now\;
      \$v5051\ := \$v5051%now\;
      \$v5679\ := \$v5679%now\;
      \$v5630\ := \$v5630%now\;
      \$19889\ := \$19889%now\;
      \$18812\ := \$18812%now\;
      \$v5543\ := \$v5543%now\;
      \$18955_modulo6684349_id\ := \$18955_modulo6684349_id%now\;
      \$19529_forever6704351_arg\ := \$19529_forever6704351_arg%now\;
      \$v5556\ := \$v5556%now\;
      \$19497_loop666_result\ := \$19497_loop666_result%now\;
      \$18536\ := \$18536%now\;
      \$19433\ := \$19433%now\;
      \$v4857\ := \$v4857%now\;
      \$19286\ := \$19286%now\;
      \$19621\ := \$19621%now\;
      \$18758\ := \$18758%now\;
      \$19261\ := \$19261%now\;
      \$v5566\ := \$v5566%now\;
      \$v4881\ := \$v4881%now\;
      \$19148_modulo6684357_result\ := \$19148_modulo6684357_result%now\;
      \$v4795\ := \$v4795%now\;
      \$19945\ := \$19945%now\;
      \$v4466\ := \$v4466%now\;
      \$v4824\ := \$v4824%now\;
      \$19747\ := \$19747%now\;
      \$19081_modulo6684349_id\ := \$19081_modulo6684349_id%now\;
      \$19285\ := \$19285%now\;
      \$v4884\ := \$v4884%now\;
      \$v5863\ := \$v5863%now\;
      \$19394_compbranch6504395_result\ := \$19394_compbranch6504395_result%now\;
      \$19535_copy_root_in_ram6634354_result\ := \$19535_copy_root_in_ram6634354_result%now\;
      \$v4758\ := \$v4758%now\;
      \$v4488\ := \$v4488%now\;
      \$19012_modulo6684349_arg\ := \$19012_modulo6684349_arg%now\;
      \$18607\ := \$18607%now\;
      \$19753\ := \$19753%now\;
      \$18785\ := \$18785%now\;
      \$19394_compbranch6504395_id\ := \$19394_compbranch6504395_id%now\;
      \$v5894\ := \$v5894%now\;
      \$18799_w1656_arg\ := \$18799_w1656_arg%now\;
      \$18856_loop_push6494360_id\ := \$18856_loop_push6494360_id%now\;
      \$v4981\ := \$v4981%now\;
      \$19391_compare6444359_arg\ := \$19391_compare6444359_arg%now\;
      \$19366_compbranch6504391_id\ := \$19366_compbranch6504391_id%now\;
      \$v4771\ := \$v4771%now\;
      \$19781_aux664_result\ := \$19781_aux664_result%now\;
      \$19174_binop_compare6454378_id\ := \$19174_binop_compare6454378_id%now\;
      \$19416_w36574398_arg\ := \$19416_w36574398_arg%now\;
      \$v5627\ := \$v5627%now\;
      \$19271\ := \$19271%now\;
      \$v5126\ := \$v5126%now\;
      \$18708\ := \$18708%now\;
      \$19780_loop665_id\ := \$19780_loop665_id%now\;
      \$18827\ := \$18827%now\;
      \$v5890\ := \$v5890%now\;
      \$18882_v\ := \$18882_v%now\;
      \$18525_loop665_arg\ := \$18525_loop665_arg%now\;
      \$v5623\ := \$v5623%now\;
      \$19344\ := \$19344%now\;
      \$19576\ := \$19576%now\;
      \$19171_compare6444358_arg\ := \$19171_compare6444358_arg%now\;
      \$19838_copy_root_in_ram6634340_id\ := \$19838_copy_root_in_ram6634340_id%now\;
      \$v5387\ := \$v5387%now\;
      \$19373_compbranch6504392_arg\ := \$19373_compbranch6504392_arg%now\;
      \$v5602\ := \$v5602%now\;
      \$18544\ := \$18544%now\;
      \$v5773\ := \$v5773%now\;
      \$18493\ := \$18493%now\;
      \$18579\ := \$18579%now\;
      \$v5444\ := \$v5444%now\;
      \$19524\ := \$19524%now\;
      \$19247\ := \$19247%now\;
      \$19122_modulo6684356_id\ := \$19122_modulo6684356_id%now\;
      \$v5585\ := \$v5585%now\;
      \$19494_loop666_result\ := \$19494_loop666_result%now\;
      \$19284\ := \$19284%now\;
      \$19373_compbranch6504392_id\ := \$19373_compbranch6504392_id%now\;
      \$19287_v\ := \$19287_v%now\;
      \$19808_forever6704342_id\ := \$19808_forever6704342_id%now\;
      \$v5459\ := \$v5459%now\;
      \$19767\ := \$19767%now\;
      \$v5181\ := \$v5181%now\;
      \$19494_loop666_id\ := \$19494_loop666_id%now\;
      \$19529_forever6704351_id\ := \$19529_forever6704351_id%now\;
      \$v5782\ := \$v5782%now\;
      \$19053_binop_int6434369_id\ := \$19053_binop_int6434369_id%now\;
      \$v4478\ := \$v4478%now\;
      \$v5495\ := \$v5495%now\;
      \$v4505\ := \$v4505%now\;
      \$18621\ := \$18621%now\;
      \$19598\ := \$19598%now\;
      \$v4774\ := \$v4774%now\;
      \$18523_aux664_result\ := \$18523_aux664_result%now\;
      \$v5919\ := \$v5919%now\;
      \$19298_v\ := \$19298_v%now\;
      \$18872_v\ := \$18872_v%now\;
      \$18817_v\ := \$18817_v%now\;
      \$19762\ := \$19762%now\;
      \$19002_modulo6684356_id\ := \$19002_modulo6684356_id%now\;
      \$v5695\ := \$v5695%now\;
      \$v5770\ := \$v5770%now\;
      \$19024_modulo6684349_arg\ := \$19024_modulo6684349_arg%now\;
      \$18936_modulo6684349_result\ := \$18936_modulo6684349_result%now\;
      \$19428\ := \$19428%now\;
      \$18890_v\ := \$18890_v%now\;
      \$v5561\ := \$v5561%now\;
      \$18535\ := \$18535%now\;
      \$19151_modulo6684349_arg\ := \$19151_modulo6684349_arg%now\;
      result4399 := \result4399%now\;
      \$19278\ := \$19278%now\;
      rdy4435 := \rdy4435%now\;
      \$19000_res\ := \$19000_res%now\;
      \$18609\ := \$18609%now\;
      \$18720\ := \$18720%now\;
      \$19552\ := \$19552%now\;
      \$18757\ := \$18757%now\;
      \$v4459\ := \$v4459%now\;
      \$19305\ := \$19305%now\;
      \$18874\ := \$18874%now\;
      \$18800\ := \$18800%now\;
      \$19607\ := \$19607%now\;
      \$v4557\ := \$v4557%now\;
      \$19757\ := \$19757%now\;
      \$v4536\ := \$v4536%now\;
      \$19933_w\ := \$19933_w%now\;
      \$v4487\ := \$v4487%now\;
      \$19258\ := \$19258%now\;
      \$v4720\ := \$v4720%now\;
      \$19151_modulo6684349_id\ := \$19151_modulo6684349_id%now\;
      \$19744_w\ := \$19744_w%now\;
      result4572 := \result4572%now\;
      \$19103_r\ := \$19103_r%now\;
      \$v5562\ := \$v5562%now\;
      \$19178_res\ := \$19178_res%now\;
      \$19160\ := \$19160%now\;
      \$19663\ := \$19663%now\;
      \$18871\ := \$18871%now\;
      \$v5332\ := \$v5332%now\;
      \$v5045\ := \$v5045%now\;
      \$19193_v\ := \$19193_v%now\;
      \$v4670\ := \$v4670%now\;
      \$v5880\ := \$v5880%now\;
      \$v5030\ := \$v5030%now\;
      \$18883_v\ := \$18883_v%now\;
      \$v4333\ := \$v4333%now\;
      \$v5572\ := \$v5572%now\;
      \$18983_modulo6684356_result\ := \$18983_modulo6684356_result%now\;
      \$19493\ := \$19493%now\;
      \$19095_res\ := \$19095_res%now\;
      \$v5756\ := \$v5756%now\;
      \$18983_modulo6684356_arg\ := \$18983_modulo6684356_arg%now\;
      \$v5114\ := \$v5114%now\;
      \$v5192\ := \$v5192%now\;
      \$19461\ := \$19461%now\;
      \$19107_modulo6684349_result\ := \$19107_modulo6684349_result%now\;
      \$18839\ := \$18839%now\;
      \$v5341\ := \$v5341%now\;
      \$v5626\ := \$v5626%now\;
      \$19050_modulo6684349_id\ := \$19050_modulo6684349_id%now\;
      \$18787\ := \$18787%now\;
      \$18716\ := \$18716%now\;
      \$19121_r\ := \$19121_r%now\;
      \$19206_binop_compare6454382_id\ := \$19206_binop_compare6454382_id%now\;
      \$18885_v\ := \$18885_v%now\;
      \$18658\ := \$18658%now\;
      \$v5851\ := \$v5851%now\;
      \$19069_modulo6684349_result\ := \$19069_modulo6684349_result%now\;
      \$v5111\ := \$v5111%now\;
      \$18678\ := \$18678%now\;
      \$19822\ := \$19822%now\;
      \$v5510\ := \$v5510%now\;
      \$18753\ := \$18753%now\;
      \$v5848\ := \$v5848%now\;
      \$19113_forever6704372_arg\ := \$19113_forever6704372_arg%now\;
      \$18840_v\ := \$18840_v%now\;
      \$v5362\ := \$v5362%now\;
      \$v4905\ := \$v4905%now\;
      \$18596\ := \$18596%now\;
      \$v4553\ := \$v4553%now\;
      \$v5218\ := \$v5218%now\;
      \$18440_make_block579_result\ := \$18440_make_block579_result%now\;
      \$19401_compbranch6504396_id\ := \$19401_compbranch6504396_id%now\;
      \$19380_compbranch6504393_result\ := \$19380_compbranch6504393_result%now\;
      \$19047_modulo6684357_arg\ := \$19047_modulo6684357_arg%now\;
      \$18861\ := \$18861%now\;
      \$19931\ := \$19931%now\;
      \$19340_argument2\ := \$19340_argument2%now\;
      \$v4991\ := \$v4991%now\;
      \$18983_modulo6684356_id\ := \$18983_modulo6684356_id%now\;
      \$v5591\ := \$v5591%now\;
      \$v5211\ := \$v5211%now\;
      \$18920_binop_int6434362_id\ := \$18920_binop_int6434362_id%now\;
      \$v5531\ := \$v5531%now\;
      \$19002_modulo6684356_result\ := \$19002_modulo6684356_result%now\;
      \$v4890\ := \$v4890%now\;
      \$18589\ := \$18589%now\;
      \$19144_modulo6684349_arg\ := \$19144_modulo6684349_arg%now\;
      \$v4600\ := \$v4600%now\;
      \$19476_v\ := \$19476_v%now\;
      \$19587\ := \$19587%now\;
      \$19919\ := \$19919%now\;
      \$19574_w\ := \$19574_w%now\;
      \$19237_v\ := \$19237_v%now\;
      \$19037_v\ := \$19037_v%now\;
      \$v5483\ := \$v5483%now\;
      \$19634\ := \$19634%now\;
      \$18585\ := \$18585%now\;
      \$v4432\ := \$v4432%now\;
      \$19365\ := \$19365%now\;
      \$v5736\ := \$v5736%now\;
      \$v4332\ := \$v4332%now\;
      \$19857\ := \$19857%now\;
      \$v5868\ := \$v5868%now\;
      \$18803\ := \$18803%now\;
      \$19346_sp\ := \$19346_sp%now\;
      \$18691\ := \$18691%now\;
      \$19846\ := \$19846%now\;
      \$v5841\ := \$v5841%now\;
      \$19695\ := \$19695%now\;
      \$19494_loop666_arg\ := \$19494_loop666_arg%now\;
      \$v5177\ := \$v5177%now\;
      \$v4707\ := \$v4707%now\;
      \$19122_modulo6684356_arg\ := \$19122_modulo6684356_arg%now\;
      \$v4737\ := \$v4737%now\;
      \$v5712\ := \$v5712%now\;
      \$19370_compare6444359_arg\ := \$19370_compare6444359_arg%now\;
      \$19622\ := \$19622%now\;
      \$v4567\ := \$v4567%now\;
      \$v5500\ := \$v5500%now\;
      \$19899\ := \$19899%now\;
      \$v5918\ := \$v5918%now\;
      \$v5408\ := \$v5408%now\;
      \$19039_r\ := \$19039_r%now\;
      \$18814\ := \$18814%now\;
      \$19738\ := \$19738%now\;
      \$19670\ := \$19670%now\;
      \$19457\ := \$19457%now\;
      \$19377_compare6444359_id\ := \$19377_compare6444359_id%now\;
      \$19556\ := \$19556%now\;
      \$19711\ := \$19711%now\;
      \$v5808\ := \$v5808%now\;
      \$19377_compare6444359_arg\ := \$19377_compare6444359_arg%now\;
      \$19405_compare6444359_result\ := \$19405_compare6444359_result%now\;
      \$v5593\ := \$v5593%now\;
      \$19903_next\ := \$19903_next%now\;
      \$18818_v\ := \$18818_v%now\;
      \$18633\ := \$18633%now\;
      \$18466_loop666_arg\ := \$18466_loop666_arg%now\;
      \$19459\ := \$19459%now\;
      \$19705\ := \$19705%now\;
      \$19629_hd\ := \$19629_hd%now\;
      \$18836_v\ := \$18836_v%now\;
      \$19384_compare6444359_arg\ := \$19384_compare6444359_arg%now\;
      \$18736\ := \$18736%now\;
      \$v5110\ := \$v5110%now\;
      \$18671\ := \$18671%now\;
      \$18686\ := \$18686%now\;
      \$v4526\ := \$v4526%now\;
      \$18990_modulo6684357_arg\ := \$18990_modulo6684357_arg%now\;
      \$v5493\ := \$v5493%now\;
      \$19632\ := \$19632%now\;
      \$v5871\ := \$v5871%now\;
      \$18823_v\ := \$18823_v%now\;
      \$18593\ := \$18593%now\;
      \$v5229\ := \$v5229%now\;
      \$v5302\ := \$v5302%now\;
      \$18652_w\ := \$18652_w%now\;
      \$19506\ := \$19506%now\;
      \$19337_compare6444359_result\ := \$19337_compare6444359_result%now\;
      \$v4411\ := \$v4411%now\;
      \$19680\ := \$19680%now\;
      rdy4964 := \rdy4964%now\;
      \$18690\ := \$18690%now\;
      \$v4755\ := \$v4755%now\;
      \$v5615\ := \$v5615%now\;
      \$19195_compare6444358_id\ := \$19195_compare6444358_id%now\;
      \$19912\ := \$19912%now\;
      \$18469_make_block579_arg\ := \$18469_make_block579_arg%now\;
      \$18743\ := \$18743%now\;
      \$19791\ := \$19791%now\;
      \$19604\ := \$19604%now\;
      \$v5805\ := \$v5805%now\;
      \$19510\ := \$19510%now\;
      \$18728\ := \$18728%now\;
      \$19869\ := \$19869%now\;
      \$19900\ := \$19900%now\;
      \$19898\ := \$19898%now\;
      \$19111\ := \$19111%now\;
      \$18586\ := \$18586%now\;
      \$18986_modulo6684349_id\ := \$18986_modulo6684349_id%now\;
      \$18468_wait662_id\ := \$18468_wait662_id%now\;
      \$19244_v\ := \$19244_v%now\;
      \$19612\ := \$19612%now\;
      \$v4785\ := \$v4785%now\;
      \$19847\ := \$19847%now\;
      \$19398_compare6444359_arg\ := \$19398_compare6444359_arg%now\;
      \$v4987\ := \$v4987%now\;
      \$19830\ := \$19830%now\;
      \$19034_binop_int6434368_id\ := \$19034_binop_int6434368_id%now\;
      \$18856_loop_push6494360_result\ := \$18856_loop_push6494360_result%now\;
      \$19687_w\ := \$19687_w%now\;
      \$19745_hd\ := \$19745_hd%now\;
      \$18894_v\ := \$18894_v%now\;
      \$v5887\ := \$v5887%now\;
      \$18672\ := \$18672%now\;
      \$18617\ := \$18617%now\;
      \$19938\ := \$19938%now\;
      \$18892_v\ := \$18892_v%now\;
      \$19437\ := \$19437%now\;
      \$18636\ := \$18636%now\;
      \$18611\ := \$18611%now\;
      \$19225\ := \$19225%now\;
      \$19420_w06554397_arg\ := \$19420_w06554397_arg%now\;
      \$18713\ := \$18713%now\;
      \$18616\ := \$18616%now\;
      \$18771\ := \$18771%now\;
      \$v4635\ := \$v4635%now\;
      \$v5792\ := \$v5792%now\;
      \$18868_v\ := \$18868_v%now\;
      \$v5106\ := \$v5106%now\;
      \$18693\ := \$18693%now\;
      \$18597\ := \$18597%now\;
      \$18437_loop666_result\ := \$18437_loop666_result%now\;
      \$19426\ := \$19426%now\;
      \$19763\ := \$19763%now\;
      \$v5575\ := \$v5575%now\;
      \$v4747\ := \$v4747%now\;
      \$v5381\ := \$v5381%now\;
      \$19151_modulo6684349_result\ := \$19151_modulo6684349_result%now\;
      \$v5474\ := \$v5474%now\;
      \$18850\ := \$18850%now\;
      \$18445_x\ := \$18445_x%now\;
      \$18798_w652_arg\ := \$18798_w652_arg%now\;
      \$18878\ := \$18878%now\;
      \$v5820\ := \$v5820%now\;
      \$v5022\ := \$v5022%now\;
      \$v4968\ := \$v4968%now\;
      \$v4686\ := \$v4686%now\;
      \$19472\ := \$19472%now\;
      \$v5718\ := \$v5718%now\;
      \$19404_b\ := \$19404_b%now\;
      \$v4446\ := \$v4446%now\;
      \$19624\ := \$19624%now\;
      \$18587\ := \$18587%now\;
      \$v5906\ := \$v5906%now\;
      \$18970_r\ := \$18970_r%now\;
      \$19545\ := \$19545%now\;
      \$18534_next\ := \$18534_next%now\;
      \$19219\ := \$19219%now\;
      \$18792_wait662_id\ := \$18792_wait662_id%now\;
      \$19265_ofs\ := \$19265_ofs%now\;
      \$19618\ := \$19618%now\;
      \$19411\ := \$19411%now\;
      \$19468_sp\ := \$19468_sp%now\;
      \$18547\ := \$18547%now\;
      \$19116_binop_int6434373_id\ := \$19116_binop_int6434373_id%now\;
      \$19065_r\ := \$19065_r%now\;
      \$19645\ := \$19645%now\;
      \$19129_modulo6684357_result\ := \$19129_modulo6684357_result%now\;
      \$v5155\ := \$v5155%now\;
      \$v5219\ := \$v5219%now\;
      \$19756\ := \$19756%now\;
      \$18490\ := \$18490%now\;
      \$18523_aux664_arg\ := \$18523_aux664_arg%now\;
      \$v5375\ := \$v5375%now\;
      \$19215_argument1\ := \$19215_argument1%now\;
      \$18860\ := \$18860%now\;
      \$v5898\ := \$v5898%now\;
      \$v4643\ := \$v4643%now\;
      \$19174_binop_compare6454378_arg\ := \$19174_binop_compare6454378_arg%now\;
      \$v5581\ := \$v5581%now\;
      \$v4999\ := \$v4999%now\;
      \$18466_loop666_result\ := \$18466_loop666_result%now\;
      \$18469_make_block579_result\ := \$18469_make_block579_result%now\;
      \$18625_copy_root_in_ram6634345_result\ := \$18625_copy_root_in_ram6634345_result%now\;
      \$19640\ := \$19640%now\;
      \$v4657\ := \$v4657%now\;
      \$v5501\ := \$v5501%now\;
      \$19323\ := \$19323%now\;
      \$v5631\ := \$v5631%now\;
      \$19270\ := \$19270%now\;
      \$19473\ := \$19473%now\;
      \$19318\ := \$19318%now\;
      \$19132_modulo6684349_result\ := \$19132_modulo6684349_result%now\;
      \$18548\ := \$18548%now\;
      \$18967_modulo6684349_id\ := \$18967_modulo6684349_id%now\;
      \$18772\ := \$18772%now\;
      \$18628\ := \$18628%now\;
      \$19562\ := \$19562%now\;
      \$18538\ := \$18538%now\;
      \$18819_v\ := \$18819_v%now\;
      \$19198_binop_compare6454381_arg\ := \$19198_binop_compare6454381_arg%now\;
      \$19465_sp\ := \$19465_sp%now\;
      \$18526_aux664_result\ := \$18526_aux664_result%now\;
      \$19911\ := \$19911%now\;
      \$v4914\ := \$v4914%now\;
      \$19446_sp\ := \$19446_sp%now\;
      \$18932_r\ := \$18932_r%now\;
      \$v4463\ := \$v4463%now\;
      \$19946\ := \$19946%now\;
      \$19943\ := \$19943%now\;
      \$v5372\ := \$v5372%now\;
      \$19577\ := \$19577%now\;
      \$18641\ := \$18641%now\;
      \$18773\ := \$18773%now\;
      \$v5740\ := \$v5740%now\;
      \$18524_loop666_id\ := \$18524_loop666_id%now\;
      \$18964_modulo6684356_result\ := \$18964_modulo6684356_result%now\;
      \$v4427\ := \$v4427%now\;
      \$19655\ := \$19655%now\;
      \$19028_modulo6684357_arg\ := \$19028_modulo6684357_arg%now\;
      \$v4788\ := \$v4788%now\;
      \$19520\ := \$19520%now\;
      \$v4875\ := \$v4875%now\;
      \$19306_v\ := \$19306_v%now\;
      \$v5567\ := \$v5567%now\;
      \$v5521\ := \$v5521%now\;
      \$v4644\ := \$v4644%now\;
      \$19343_sp\ := \$19343_sp%now\;
      \$18722\ := \$18722%now\;
      \$19935\ := \$19935%now\;
      \$19056_v\ := \$19056_v%now\;
      \$18513\ := \$18513%now\;
      \$18989_r\ := \$18989_r%now\;
      \$18879_v\ := \$18879_v%now\;
      \$v4956\ := \$v4956%now\;
      \$19730\ := \$19730%now\;
      \$18665\ := \$18665%now\;
      \$v4452\ := \$v4452%now\;
      \$v5783\ := \$v5783%now\;
      \$18710\ := \$18710%now\;
      \$v5676\ := \$v5676%now\;
      \$19009_modulo6684357_id\ := \$19009_modulo6684357_id%now\;
      \$19712\ := \$19712%now\;
      \$19841\ := \$19841%now\;
      \$18556_forever6704344_arg\ := \$18556_forever6704344_arg%now\;
      \$19780_loop665_result\ := \$19780_loop665_result%now\;
      \$19236_v\ := \$19236_v%now\;
      \$19330_compare6444359_result\ := \$19330_compare6444359_result%now\;
      \$v5600\ := \$v5600%now\;
      \$19330_compare6444359_arg\ := \$19330_compare6444359_arg%now\;
      \$18592\ := \$18592%now\;
      \$19289\ := \$19289%now\;
      \$19589_copy_root_in_ram6634353_arg\ := \$19589_copy_root_in_ram6634353_arg%now\;
      \$v4778\ := \$v4778%now\;
      \$19356\ := \$19356%now\;
      \$19050_modulo6684349_arg\ := \$19050_modulo6684349_arg%now\;
      \$v5241\ := \$v5241%now\;
      \$18594\ := \$18594%now\;
      \$v5680\ := \$v5680%now\;
      \$18866_v\ := \$18866_v%now\;
      \$v5877\ := \$v5877%now\;
      \$19424\ := \$19424%now\;
      \$v5587\ := \$v5587%now\;
      \$19369_b\ := \$19369_b%now\;
      \$18481\ := \$18481%now\;
      \$19050_modulo6684349_result\ := \$19050_modulo6684349_result%now\;
      \$19691\ := \$19691%now\;
      \$18471\ := \$18471%now\;
      \$19058_r\ := \$19058_r%now\;
      \$19560_hd\ := \$19560_hd%now\;
      \$19405_compare6444359_id\ := \$19405_compare6444359_id%now\;
      \$v5901\ := \$v5901%now\;
      \$v5435\ := \$v5435%now\;
      \$19353\ := \$19353%now\;
      \$19059_modulo6684356_result\ := \$19059_modulo6684356_result%now\;
      \$18910_modulo6684349_arg\ := \$18910_modulo6684349_arg%now\;
      \$v5706\ := \$v5706%now\;
      \$18486\ := \$18486%now\;
      \$18501\ := \$18501%now\;
      \$18532\ := \$18532%now\;
      \$v4764\ := \$v4764%now\;
      \$19216_v\ := \$19216_v%now\;
      \$19613_w\ := \$19613_w%now\;
      \$18528\ := \$18528%now\;
      \$19283\ := \$19283%now\;
      \$v5338\ := \$v5338%now\;
      \$19091_binop_int6434371_result\ := \$19091_binop_int6434371_result%now\;
      \$v4962\ := \$v4962%now\;
      \$19654\ := \$19654%now\;
      \$v5842\ := \$v5842%now\;
      \$v5527\ := \$v5527%now\;
      \$18920_binop_int6434362_result\ := \$18920_binop_int6434362_result%now\;
      \$19195_compare6444358_arg\ := \$19195_compare6444358_arg%now\;
      \$v5910\ := \$v5910%now\;
      \$18705_next\ := \$18705_next%now\;
      \$19511\ := \$19511%now\;
      \$v5902\ := \$v5902%now\;
      \$19410\ := \$19410%now\;
      \$18468_wait662_arg\ := \$18468_wait662_arg%now\;
      \$v5504\ := \$v5504%now\;
      \$v4522\ := \$v4522%now\;
      \$18797_branch_if648_arg\ := \$18797_branch_if648_arg%now\;
      \$19696\ := \$19696%now\;
      \$18955_modulo6684349_arg\ := \$18955_modulo6684349_arg%now\;
      \$19652\ := \$19652%now\;
      \$19606\ := \$19606%now\;
      \$19195_compare6444358_result\ := \$19195_compare6444358_result%now\;
      \$v5006\ := \$v5006%now\;
      \$18804\ := \$18804%now\;
      \$18910_modulo6684349_result\ := \$18910_modulo6684349_result%now\;
      \$19502\ := \$19502%now\;
      \$v5583\ := \$v5583%now\;
      \$18853_hd\ := \$18853_hd%now\;
      \$v5746\ := \$v5746%now\;
      \$v5048\ := \$v5048%now\;
      \$19831\ := \$19831%now\;
      \$19481\ := \$19481%now\;
      \$18774\ := \$18774%now\;
      \$19708\ := \$19708%now\;
      \$18632\ := \$18632%now\;
      \$18625_copy_root_in_ram6634345_arg\ := \$18625_copy_root_in_ram6634345_arg%now\;
      \$v5834\ := \$v5834%now\;
      \$19568\ := \$19568%now\;
      \$v4723\ := \$v4723%now\;
      \$18519\ := \$18519%now\;
      \$v4580\ := \$v4580%now\;
      \$19547_copy_root_in_ram6634352_arg\ := \$19547_copy_root_in_ram6634352_arg%now\;
      \$19477_v\ := \$19477_v%now\;
      \$18704\ := \$18704%now\;
      \$18503\ := \$18503%now\;
      \$18790_loop666_arg\ := \$18790_loop666_arg%now\;
      \$v5854\ := \$v5854%now\;
      \$19690\ := \$19690%now\;
      \$v5786\ := \$v5786%now\;
      \$19498_loop665_id\ := \$19498_loop665_id%now\;
      \$v5864\ := \$v5864%now\;
      \$v5886\ := \$v5886%now\;
      \$18923_v\ := \$18923_v%now\;
      \$v5914\ := \$v5914%now\;
      \$v5798\ := \$v5798%now\;
      \$v5016\ := \$v5016%now\;
      \$19499_aux664_result\ := \$19499_aux664_result%now\;
      \$v5554\ := \$v5554%now\;
      \$18675\ := \$18675%now\;
      \$18463\ := \$18463%now\;
      \$19469\ := \$19469%now\;
      \$18700\ := \$18700%now\;
      \$18744_w\ := \$18744_w%now\;
      \$v5087\ := \$v5087%now\;
      \$18530\ := \$18530%now\;
      \$v5423\ := \$v5423%now\;
      \$v5215\ := \$v5215%now\;
      \$18929_modulo6684349_result\ := \$18929_modulo6684349_result%now\;
      \$19733\ := \$19733%now\;
      \$18653_hd\ := \$18653_hd%now\;
      \$19429\ := \$19429%now\;
      \$18833\ := \$18833%now\;
      \$v5165\ := \$v5165%now\;
      \$18454\ := \$18454%now\;
      \$18847\ := \$18847%now\;
      \$v5553\ := \$v5553%now\;
      \$v5075\ := \$v5075%now\;
      \$18692\ := \$18692%now\;
      \$18719\ := \$18719%now\;
      \$19940\ := \$19940%now\;
      \$18712_hd\ := \$18712_hd%now\;
      \$v5417\ := \$v5417%now\;
      \$19125_modulo6684349_arg\ := \$19125_modulo6684349_arg%now\;
      \$18634\ := \$18634%now\;
      \$19484\ := \$19484%now\;
      \$18929_modulo6684349_id\ := \$18929_modulo6684349_id%now\;
      \$19198_binop_compare6454381_id\ := \$19198_binop_compare6454381_id%now\;
      \$19416_w36574398_id\ := \$19416_w36574398_id%now\;
      \$18798_w652_id\ := \$18798_w652_id%now\;
      \$v5056\ := \$v5056%now\;
      \$v4439\ := \$v4439%now\;
      \$v5503\ := \$v5503%now\;
      \$19608\ := \$19608%now\;
      \$v5779\ := \$v5779%now\;
      \$19277\ := \$19277%now\;
      \$19223\ := \$19223%now\;
      \$18499\ := \$18499%now\;
      \$18796_make_block_n646_result\ := \$18796_make_block_n646_result%now\;
      \$19085_modulo6684357_id\ := \$19085_modulo6684357_id%now\;
      \$v5399\ := \$v5399%now\;
      \$v4808\ := \$v4808%now\;
      \$18811\ := \$18811%now\;
      \$19808_forever6704342_arg\ := \$19808_forever6704342_arg%now\;
      \$v4508\ := \$v4508%now\;
      \$v5207\ := \$v5207%now\;
      \$v5093\ := \$v5093%now\;
      \$19034_binop_int6434368_result\ := \$19034_binop_int6434368_result%now\;
      \$19627\ := \$19627%now\;
      \$19881_hd\ := \$19881_hd%now\;
      \$19291_v\ := \$19291_v%now\;
      \$18901_binop_int6434361_id\ := \$18901_binop_int6434361_id%now\;
      \$19387_compbranch6504394_result\ := \$19387_compbranch6504394_result%now\;
      \$19644_hd\ := \$19644_hd%now\;
      \$19347_fill6534389_id\ := \$19347_fill6534389_id%now\;
      \$v5917\ := \$v5917%now\;
      \$19792\ := \$19792%now\;
      \$19541\ := \$19541%now\;
      \$v5480\ := \$v5480%now\;
      \$19415_sp\ := \$19415_sp%now\;
      \$19262_forever6704385_arg\ := \$19262_forever6704385_arg%now\;
      \$18477\ := \$18477%now\;
      \$19635\ := \$19635%now\;
      \$v4933\ := \$v4933%now\;
      \$19633\ := \$19633%now\;
      \$v4566\ := \$v4566%now\;
      \$18917_modulo6684349_id\ := \$18917_modulo6684349_id%now\;
      \$18451\ := \$18451%now\;
      \$19802\ := \$19802%now\;
      \$19221\ := \$19221%now\;
      \$19224\ := \$19224%now\;
      \$v5240\ := \$v5240%now\;
      \$19516\ := \$19516%now\;
      \$18656\ := \$18656%now\;
      \$19693\ := \$19693%now\;
      \$18496\ := \$18496%now\;
      \$18588\ := \$18588%now\;
      \$18887_v\ := \$18887_v%now\;
      \$19360_sp\ := \$19360_sp%now\;
      \$19171_compare6444358_result\ := \$19171_compare6444358_result%now\;
      \$19688_hd\ := \$19688_hd%now\;
      \$18491\ := \$18491%now\;
      \$18541\ := \$18541%now\;
      \$19380_compbranch6504393_arg\ := \$19380_compbranch6504393_arg%now\;
      \$19782\ := \$19782%now\;
      \$v5517\ := \$v5517%now\;
      \$19141_modulo6684356_id\ := \$19141_modulo6684356_id%now\;
      \$19107_modulo6684349_id\ := \$19107_modulo6684349_id%now\;
      \$v4971\ := \$v4971%now\;
      \$v4848\ := \$v4848%now\;
      \$19166_binop_compare6454377_result\ := \$19166_binop_compare6454377_result%now\;
      \$19593\ := \$19593%now\;
      \$18568\ := \$18568%now\;
      \$v4625\ := \$v4625%now\;
      \$18452\ := \$18452%now\;
      \$19742\ := \$19742%now\;
      \$v4869\ := \$v4869%now\;
      \$v5590\ := \$v5590%now\;
      \$18468_wait662_result\ := \$18468_wait662_result%now\;
      \$19575_hd\ := \$19575_hd%now\;
      \$19229_v\ := \$19229_v%now\;
      \$18981_res\ := \$18981_res%now\;
      \$v4622\ := \$v4622%now\;
      \$18942_v\ := \$18942_v%now\;
      \$18543\ := \$18543%now\;
      \$19513\ := \$19513%now\;
      \$19555\ := \$19555%now\;
      \$19692\ := \$19692%now\;
      \$19370_compare6444359_result\ := \$19370_compare6444359_result%now\;
      \$v4896\ := \$v4896%now\;
      \$v5661\ := \$v5661%now\;
      \$v5520\ := \$v5520%now\;
      \$18917_modulo6684349_result\ := \$18917_modulo6684349_result%now\;
      \$19116_binop_int6434373_result\ := \$19116_binop_int6434373_result%now\;
      \$v4404\ := \$v4404%now\;
      \$19862\ := \$19862%now\;
      \$18449\ := \$18449%now\;
      \$19573\ := \$19573%now\;
      \$19729\ := \$19729%now\;
      \$18952_modulo6684357_id\ := \$18952_modulo6684357_id%now\;
      \$19252_forever6704384_arg\ := \$19252_forever6704384_arg%now\;
      \$19805\ := \$19805%now\;
      \$18943_res\ := \$18943_res%now\;
      \$v4564\ := \$v4564%now\;
      \$18926_modulo6684356_arg\ := \$18926_modulo6684356_arg%now\;
      \$v5438\ := \$v5438%now\;
      \$19567\ := \$19567%now\;
      \$18761\ := \$18761%now\;
      \$v5350\ := \$v5350%now\;
      \$v5230\ := \$v5230%now\;
      \$v4731\ := \$v4731%now\;
      \$19838_copy_root_in_ram6634340_arg\ := \$19838_copy_root_in_ram6634340_arg%now\;
      \$v5667\ := \$v5667%now\;
      \$v5535\ := \$v5535%now\;
      \$19008_r\ := \$19008_r%now\;
      \$v5547\ := \$v5547%now\;
      \$19669\ := \$19669%now\;
      \$18862\ := \$18862%now\;
      \$19699\ := \$19699%now\;
      \$19630\ := \$19630%now\;
      \$ram_lock\ := \$ram_lock%now\;
      \$global_end_lock\ := \$global_end_lock%now\;
      \$code_lock\ := \$code_lock%now\;
      state := \state%now\;
      state_var5924 := \state_var5924%now\;
      state_var5923 := \state_var5923%now\;
      state_var5922 := \state_var5922%now\;
      state_var5921 := \state_var5921%now\;
      state_var5920 := \state_var5920%now\;
      case state is
      when \$18437_LOOP666\ =>
        \$v4408\ := work.Int.ge(\$18437_loop666_arg\(0 to 15), work.Int.add(
                                                               \$18437_loop666_arg\(48 to 63), X"000" & X"1"));
        if \$v4408\(0) = '1' then
          \$18437_loop666_result\ := eclat_unit;
          \$19945\ := \$18437_loop666_result\;
          \$v4417\ := \$ram_lock\;
          if \$v4417\(0) = '1' then
            state := Q_WAIT4416;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$19930\(0 to 30),16)));
            \$ram_write\ <= eclat_resize(\$18438_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
            state := PAUSE_SET4415;
          end if;
        else
          \$v4407\ := \$ram_lock\;
          if \$v4407\(0) = '1' then
            state := Q_WAIT4406;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$18437_loop666_arg\(32 to 47), \$18437_loop666_arg\(0 to 15))));
            state := PAUSE_GET4405;
          end if;
        end if;
      when \$18438_LOOP665\ =>
        \$v4432\ := work.Int.ge(\$18438_loop665_arg\(0 to 15), work.Int.add(
                                                               \$18438_loop665_arg\(80 to 95), X"000" & X"1"));
        if \$v4432\(0) = '1' then
          \$18438_loop665_result\ := \$18438_loop665_arg\(16 to 31);
          state := \$18438_LOOP665\;
        else
          \$v4431\ := \$ram_lock\;
          if \$v4431\(0) = '1' then
            state := Q_WAIT4430;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$18438_loop665_arg\(64 to 79), \$18438_loop665_arg\(0 to 15))));
            state := PAUSE_GET4429;
          end if;
        end if;
      when \$18439_WAIT662\ =>
        if \$v4325\(0) = '1' then
          
        else
          \$v4325\ := eclat_true;
          \$19778\ := \$18439_wait662_arg\(1 to 32) & \$18439_wait662_arg\(33 to 64) & X"0" & X"fa0" & X"0" & X"fa0" & X"0" & X"fa0" & 
          work.Int.add(X"0" & X"fa0", X"1770") & eclat_false;
        end if;
        case state_var5924 is
        when \$19779_LOOP666\ =>
          \$v4443\ := work.Int.ge(\$19779_loop666_arg\(0 to 15), work.Int.add(
                                                                 \$19779_loop666_arg\(48 to 63), X"000" & X"1"));
          if \$v4443\(0) = '1' then
            \$19779_loop666_result\ := eclat_unit;
            case \$19779_loop666_id\ is
            when "000000000010" =>
              \$19921\ := \$19779_loop666_result\;
              \$v4452\ := \$ram_lock\;
              if \$v4452\(0) = '1' then
                state_var5924 := Q_WAIT4451;
              else
                acquire(\$ram_lock\);
                \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$19906\(0 to 30),16)));
                \$ram_write\ <= eclat_resize(\$19780_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                state_var5924 := PAUSE_SET4450;
              end if;
            when "000000000110" =>
              \$19835\ := \$19779_loop666_result\;
              \$v4481\ := \$ram_lock\;
              if \$v4481\(0) = '1' then
                state_var5924 := Q_WAIT4480;
              else
                acquire(\$ram_lock\);
                \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$19817\(0 to 30),16)));
                \$ram_write\ <= eclat_resize(\$19811_copy_root_in_ram6634341_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                state_var5924 := PAUSE_SET4479;
              end if;
            when "000000001000" =>
              \$19862\ := \$19779_loop666_result\;
              \$v4508\ := \$ram_lock\;
              if \$v4508\(0) = '1' then
                state_var5924 := Q_WAIT4507;
              else
                acquire(\$ram_lock\);
                \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$19844\(0 to 30),16)));
                \$ram_write\ <= eclat_resize(\$19838_copy_root_in_ram6634340_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                state_var5924 := PAUSE_SET4506;
              end if;
            when "000000001010" =>
              \$19877\ := \$19779_loop666_result\;
              \$v4529\ := \$ram_lock\;
              if \$v4529\(0) = '1' then
                state_var5924 := Q_WAIT4528;
              else
                acquire(\$ram_lock\);
                \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18439_wait662_arg\(33 to 63),16)));
                \$ram_write\ <= eclat_resize(\$19787\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                state_var5924 := PAUSE_SET4527;
              end if;
            when "000000001011" =>
              \$19892\ := \$19779_loop666_result\;
              \$v4546\ := \$ram_lock\;
              if \$v4546\(0) = '1' then
                state_var5924 := Q_WAIT4545;
              else
                acquire(\$ram_lock\);
                \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18439_wait662_arg\(1 to 31),16)));
                \$ram_write\ <= eclat_resize(\$19778\(112 to 127),31) & eclat_false; \$ram_write_request\ <= '1';
                state_var5924 := PAUSE_SET4544;
              end if;
            when others =>
              
            end case;
          else
            \$v4442\ := \$ram_lock\;
            if \$v4442\(0) = '1' then
              state_var5924 := Q_WAIT4441;
            else
              acquire(\$ram_lock\);
              \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$19779_loop666_arg\(32 to 47), \$19779_loop666_arg\(0 to 15))));
              state_var5924 := PAUSE_GET4440;
            end if;
          end if;
        when \$19780_LOOP665\ =>
          \$v4467\ := work.Int.ge(\$19780_loop665_arg\(0 to 15), work.Int.add(
                                                                 \$19780_loop665_arg\(80 to 95), X"000" & X"1"));
          if \$v4467\(0) = '1' then
            \$19780_loop665_result\ := \$19780_loop665_arg\(16 to 31);
            \$19903_next\ := \$19780_loop665_result\;
            \$19781_aux664_arg\ := work.Int.add(\$19781_aux664_arg\(0 to 15), 
                                                work.Int.add(eclat_resize(
                                                             work.Int.lsr(
                                                             eclat_resize(eclat_resize(\$19902\(0 to 30),16),31), X"0000000" & X"2"),16), X"000" & X"1")) & \$19903_next\ & \$19781_aux664_arg\(32 to 47) & \$19781_aux664_arg\(48 to 63);
            state_var5924 := \$19781_AUX664\;
          else
            \$v4466\ := \$ram_lock\;
            if \$v4466\(0) = '1' then
              state_var5924 := Q_WAIT4465;
            else
              acquire(\$ram_lock\);
              \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$19780_loop665_arg\(64 to 79), \$19780_loop665_arg\(0 to 15))));
              state_var5924 := PAUSE_GET4464;
            end if;
          end if;
        when \$19781_AUX664\ =>
          \$19897\ := work.Print.print_string(clk,of_string("     scan="));
          \$19898\ := work.Int.print(clk,\$19781_aux664_arg\(0 to 15));
          \$19899\ := work.Print.print_string(clk,of_string(" | next="));
          \$19900\ := work.Int.print(clk,\$19781_aux664_arg\(16 to 31));
          \$19901\ := work.Print.print_newline(clk,eclat_unit);
          \$v4471\ := work.Int.ge(\$19781_aux664_arg\(0 to 15), \$19781_aux664_arg\(16 to 31));
          if \$v4471\(0) = '1' then
            \$19781_aux664_result\ := \$19781_aux664_arg\(16 to 31);
            \$19800_next\ := \$19781_aux664_result\;
            \$19801\ := work.Print.print_string(clk,of_string("memory copied in to_space : "));
            \$19802\ := work.Int.print(clk,work.Int.sub(\$19800_next\, \$19778\(112 to 127)));
            \$19803\ := work.Print.print_string(clk,of_string(" words"));
            \$19804\ := work.Print.print_newline(clk,eclat_unit);
            \$v4472\ := work.Int.gt(work.Int.sub(\$19800_next\, \$19778\(112 to 127)), X"1770");
            if \$v4472\(0) = '1' then
              \$19805\ := work.Print.print_string(clk,of_string("fatal error: "));
              \$19806\ := work.Print.print_string(clk,of_string("Out of memory"));
              \$19807\ := work.Print.print_newline(clk,eclat_unit);
              \$19808_forever6704342_id\ := "000000000100";
              \$19808_forever6704342_arg\ := eclat_unit;
              state_var5924 := \$19808_FOREVER6704342\;
            else
              \$19790\ := \$19787\(0 to 31) & \$19788\(0 to 31) & \$19800_next\;
              \$19791\ := work.Print.print_newline(clk,eclat_unit);
              \$19792\ := work.Print.print_newline(clk,eclat_unit);
              \$19793\ := work.Print.print_string(clk,of_string("[================= GC END ======================]"));
              \$19794\ := work.Print.print_newline(clk,eclat_unit);
              \$19795\ := work.Print.print_newline(clk,eclat_unit);
              result4434 := \$19790\(0 to 31) & \$19790\(32 to 63) & \$19790\(64 to 79) & 
              work.Int.add(\$19790\(64 to 79), \$18439_wait662_arg\(81 to 96)) & \$19778\(112 to 127) & \$19778\(96 to 111);
              rdy4435 := eclat_true;
              state_var5924 := IDLE4436;
            end if;
          else
            \$v4470\ := \$ram_lock\;
            if \$v4470\(0) = '1' then
              state_var5924 := Q_WAIT4469;
            else
              acquire(\$ram_lock\);
              \$ram_ptr\ <= to_integer(unsigned(\$19781_aux664_arg\(0 to 15)));
              state_var5924 := PAUSE_GET4468;
            end if;
          end if;
        when \$19808_FOREVER6704342\ =>
          \$19808_forever6704342_arg\ := eclat_unit;
          state_var5924 := \$19808_FOREVER6704342\;
        when \$19811_COPY_ROOT_IN_RAM6634341\ =>
          \$v4496\ := work.Int.ge(\$19811_copy_root_in_ram6634341_arg\(0 to 15), \$19811_copy_root_in_ram6634341_arg\(16 to 31));
          if \$v4496\(0) = '1' then
            \$19811_copy_root_in_ram6634341_result\ := \$19811_copy_root_in_ram6634341_arg\(32 to 47);
            \$19797_next\ := \$19811_copy_root_in_ram6634341_result\;
            \$19798\ := work.Print.print_string(clk,of_string("======================================="));
            \$19799\ := work.Print.print_newline(clk,eclat_unit);
            \$19781_aux664_id\ := "000000000101";
            \$19781_aux664_arg\ := \$19778\(112 to 127) & \$19797_next\ & \$19778\(96 to 111) & \$19778\(112 to 127);
            state_var5924 := \$19781_AUX664\;
          else
            \$19814\ := work.Print.print_string(clk,of_string("racine:"));
            \$19815\ := work.Int.print(clk,\$19811_copy_root_in_ram6634341_arg\(0 to 15));
            \$19816\ := work.Print.print_newline(clk,eclat_unit);
            \$v4495\ := \$ram_lock\;
            if \$v4495\(0) = '1' then
              state_var5924 := Q_WAIT4494;
            else
              acquire(\$ram_lock\);
              \$ram_ptr\ <= to_integer(unsigned(\$19811_copy_root_in_ram6634341_arg\(0 to 15)));
              state_var5924 := PAUSE_GET4493;
            end if;
          end if;
        when \$19838_COPY_ROOT_IN_RAM6634340\ =>
          \$v4523\ := work.Int.ge(\$19838_copy_root_in_ram6634340_arg\(0 to 15), \$19838_copy_root_in_ram6634340_arg\(16 to 31));
          if \$v4523\(0) = '1' then
            \$19838_copy_root_in_ram6634340_result\ := \$19838_copy_root_in_ram6634340_arg\(32 to 47);
            \$19789_next\ := \$19838_copy_root_in_ram6634340_result\;
            \$v4499\ := \$global_end_lock\;
            if \$v4499\(0) = '1' then
              state_var5924 := Q_WAIT4498;
            else
              acquire(\$global_end_lock\);
              \$global_end_ptr\ <= 0;
              state_var5924 := PAUSE_GET4497;
            end if;
          else
            \$19841\ := work.Print.print_string(clk,of_string("racine:"));
            \$19842\ := work.Int.print(clk,\$19838_copy_root_in_ram6634340_arg\(0 to 15));
            \$19843\ := work.Print.print_newline(clk,eclat_unit);
            \$v4522\ := \$ram_lock\;
            if \$v4522\(0) = '1' then
              state_var5924 := Q_WAIT4521;
            else
              acquire(\$ram_lock\);
              \$ram_ptr\ <= to_integer(unsigned(\$19838_copy_root_in_ram6634340_arg\(0 to 15)));
              state_var5924 := PAUSE_GET4520;
            end if;
          end if;
        when PAUSE_GET4440 =>
          \$19926\ := \$ram_value\;
          release(\$ram_lock\);
          \$v4439\ := \$ram_lock\;
          if \$v4439\(0) = '1' then
            state_var5924 := Q_WAIT4438;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(\$19779_loop666_arg\(16 to 31), \$19779_loop666_arg\(0 to 15))));
            \$ram_write\ <= \$19926\; \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4437;
          end if;
        when PAUSE_GET4456 =>
          \$19910_hd\ := \$ram_value\;
          release(\$ram_lock\);
          \$19911\ := work.Print.print_string(clk,of_string("bloc "));
          \$19912\ := work.Int.print(clk,eclat_resize(\$19906\(0 to 30),16));
          \$19913\ := work.Print.print_string(clk,of_string(" of size "));
          \$19914\ := work.Int.print(clk,work.Int.add(eclat_resize(work.Int.lsr(
                                                                   \$19910_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
          \$19915\ := work.Print.print_string(clk,of_string(" from "));
          \$19916\ := work.Int.print(clk,eclat_resize(\$19906\(0 to 30),16));
          \$19917\ := work.Print.print_string(clk,of_string(" to "));
          \$19918\ := work.Int.print(clk,\$19780_loop665_arg\(16 to 31));
          \$19919\ := work.Print.print_newline(clk,eclat_unit);
          \$v4455\ := \$ram_lock\;
          if \$v4455\(0) = '1' then
            state_var5924 := Q_WAIT4454;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(\$19780_loop665_arg\(16 to 31)));
            \$ram_write\ <= \$19910_hd\; \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4453;
          end if;
        when PAUSE_GET4460 =>
          \$19909_w\ := \$ram_value\;
          release(\$ram_lock\);
          \$v4459\ := eclat_if(work.Bool.lnot(""&\$19909_w\(31)) & eclat_if(
                                                                   work.Int.le(
                                                                   \$19780_loop665_arg\(48 to 63), eclat_resize(\$19909_w\(0 to 30),16)) & 
                                                                   work.Int.lt(
                                                                   eclat_resize(\$19909_w\(0 to 30),16), 
                                                                   work.Int.add(
                                                                   \$19780_loop665_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false);
          if \$v4459\(0) = '1' then
            \$19907\ := \$19909_w\ & \$19780_loop665_arg\(16 to 31);
            \$v4446\ := \$ram_lock\;
            if \$v4446\(0) = '1' then
              state_var5924 := Q_WAIT4445;
            else
              acquire(\$ram_lock\);
              \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(\$19780_loop665_arg\(64 to 79), \$19780_loop665_arg\(0 to 15))));
              \$ram_write\ <= \$19907\(0 to 31); \$ram_write_request\ <= '1';
              state_var5924 := PAUSE_SET4444;
            end if;
          else
            \$v4458\ := \$ram_lock\;
            if \$v4458\(0) = '1' then
              state_var5924 := Q_WAIT4457;
            else
              acquire(\$ram_lock\);
              \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$19906\(0 to 30),16)));
              state_var5924 := PAUSE_GET4456;
            end if;
          end if;
        when PAUSE_GET4464 =>
          \$19906\ := \$ram_value\;
          release(\$ram_lock\);
          \$v4463\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$19906\(31)) & 
                                     eclat_if(work.Int.le(\$19780_loop665_arg\(32 to 47), eclat_resize(\$19906\(0 to 30),16)) & 
                                     work.Int.lt(eclat_resize(\$19906\(0 to 30),16), 
                                                 work.Int.add(\$19780_loop665_arg\(32 to 47), X"1770")) & eclat_false) & eclat_false));
          if \$v4463\(0) = '1' then
            \$19907\ := \$19906\ & \$19780_loop665_arg\(16 to 31);
            \$v4446\ := \$ram_lock\;
            if \$v4446\(0) = '1' then
              state_var5924 := Q_WAIT4445;
            else
              acquire(\$ram_lock\);
              \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(\$19780_loop665_arg\(64 to 79), \$19780_loop665_arg\(0 to 15))));
              \$ram_write\ <= \$19907\(0 to 31); \$ram_write_request\ <= '1';
              state_var5924 := PAUSE_SET4444;
            end if;
          else
            \$v4462\ := \$ram_lock\;
            if \$v4462\(0) = '1' then
              state_var5924 := Q_WAIT4461;
            else
              acquire(\$ram_lock\);
              \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19906\(0 to 30),16), X"000" & X"1")));
              state_var5924 := PAUSE_GET4460;
            end if;
          end if;
        when PAUSE_GET4468 =>
          \$19902\ := \$ram_value\;
          release(\$ram_lock\);
          \$19780_loop665_id\ := "000000000011";
          \$19780_loop665_arg\ := X"000" & X"1" & \$19781_aux664_arg\(16 to 31) & \$19781_aux664_arg\(32 to 47) & \$19781_aux664_arg\(48 to 63) & \$19781_aux664_arg\(0 to 15) & eclat_resize(
          work.Int.lsr(eclat_resize(eclat_resize(\$19902\(0 to 30),16),31), X"0000000" & X"2"),16);
          state_var5924 := \$19780_LOOP665\;
        when PAUSE_GET4485 =>
          \$19824_hd\ := \$ram_value\;
          release(\$ram_lock\);
          \$19825\ := work.Print.print_string(clk,of_string("bloc "));
          \$19826\ := work.Int.print(clk,eclat_resize(\$19817\(0 to 30),16));
          \$19827\ := work.Print.print_string(clk,of_string(" of size "));
          \$19828\ := work.Int.print(clk,work.Int.add(eclat_resize(work.Int.lsr(
                                                                   \$19824_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
          \$19829\ := work.Print.print_string(clk,of_string(" from "));
          \$19830\ := work.Int.print(clk,eclat_resize(\$19817\(0 to 30),16));
          \$19831\ := work.Print.print_string(clk,of_string(" to "));
          \$19832\ := work.Int.print(clk,\$19811_copy_root_in_ram6634341_arg\(32 to 47));
          \$19833\ := work.Print.print_newline(clk,eclat_unit);
          \$v4484\ := \$ram_lock\;
          if \$v4484\(0) = '1' then
            state_var5924 := Q_WAIT4483;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(\$19811_copy_root_in_ram6634341_arg\(32 to 47)));
            \$ram_write\ <= \$19824_hd\; \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4482;
          end if;
        when PAUSE_GET4489 =>
          \$19823_w\ := \$ram_value\;
          release(\$ram_lock\);
          \$v4488\ := eclat_if(work.Bool.lnot(""&\$19823_w\(31)) & eclat_if(
                                                                   work.Int.le(
                                                                   \$19811_copy_root_in_ram6634341_arg\(64 to 79), eclat_resize(\$19823_w\(0 to 30),16)) & 
                                                                   work.Int.lt(
                                                                   eclat_resize(\$19823_w\(0 to 30),16), 
                                                                   work.Int.add(
                                                                   \$19811_copy_root_in_ram6634341_arg\(64 to 79), X"1770")) & eclat_false) & eclat_false);
          if \$v4488\(0) = '1' then
            \$19818\ := \$19823_w\ & \$19811_copy_root_in_ram6634341_arg\(32 to 47);
            \$v4475\ := \$ram_lock\;
            if \$v4475\(0) = '1' then
              state_var5924 := Q_WAIT4474;
            else
              acquire(\$ram_lock\);
              \$ram_ptr_write\ <= to_integer(unsigned(\$19811_copy_root_in_ram6634341_arg\(0 to 15)));
              \$ram_write\ <= \$19818\(0 to 31); \$ram_write_request\ <= '1';
              state_var5924 := PAUSE_SET4473;
            end if;
          else
            \$v4487\ := \$ram_lock\;
            if \$v4487\(0) = '1' then
              state_var5924 := Q_WAIT4486;
            else
              acquire(\$ram_lock\);
              \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$19817\(0 to 30),16)));
              state_var5924 := PAUSE_GET4485;
            end if;
          end if;
        when PAUSE_GET4493 =>
          \$19817\ := \$ram_value\;
          release(\$ram_lock\);
          \$v4492\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$19817\(31)) & 
                                     eclat_if(work.Int.le(\$19811_copy_root_in_ram6634341_arg\(48 to 63), eclat_resize(\$19817\(0 to 30),16)) & 
                                     work.Int.lt(eclat_resize(\$19817\(0 to 30),16), 
                                                 work.Int.add(\$19811_copy_root_in_ram6634341_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false));
          if \$v4492\(0) = '1' then
            \$19818\ := \$19817\ & \$19811_copy_root_in_ram6634341_arg\(32 to 47);
            \$v4475\ := \$ram_lock\;
            if \$v4475\(0) = '1' then
              state_var5924 := Q_WAIT4474;
            else
              acquire(\$ram_lock\);
              \$ram_ptr_write\ <= to_integer(unsigned(\$19811_copy_root_in_ram6634341_arg\(0 to 15)));
              \$ram_write\ <= \$19818\(0 to 31); \$ram_write_request\ <= '1';
              state_var5924 := PAUSE_SET4473;
            end if;
          else
            \$v4491\ := \$ram_lock\;
            if \$v4491\(0) = '1' then
              state_var5924 := Q_WAIT4490;
            else
              acquire(\$ram_lock\);
              \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19817\(0 to 30),16), X"000" & X"1")));
              state_var5924 := PAUSE_GET4489;
            end if;
          end if;
        when PAUSE_GET4497 =>
          \$19796\ := \$global_end_value\;
          release(\$global_end_lock\);
          \$19811_copy_root_in_ram6634341_id\ := "000000000111";
          \$19811_copy_root_in_ram6634341_arg\ := X"3e80" & \$19796\ & \$19789_next\ & \$19778\(96 to 111) & \$19778\(112 to 127);
          state_var5924 := \$19811_COPY_ROOT_IN_RAM6634341\;
        when PAUSE_GET4512 =>
          \$19851_hd\ := \$ram_value\;
          release(\$ram_lock\);
          \$19852\ := work.Print.print_string(clk,of_string("bloc "));
          \$19853\ := work.Int.print(clk,eclat_resize(\$19844\(0 to 30),16));
          \$19854\ := work.Print.print_string(clk,of_string(" of size "));
          \$19855\ := work.Int.print(clk,work.Int.add(eclat_resize(work.Int.lsr(
                                                                   \$19851_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
          \$19856\ := work.Print.print_string(clk,of_string(" from "));
          \$19857\ := work.Int.print(clk,eclat_resize(\$19844\(0 to 30),16));
          \$19858\ := work.Print.print_string(clk,of_string(" to "));
          \$19859\ := work.Int.print(clk,\$19838_copy_root_in_ram6634340_arg\(32 to 47));
          \$19860\ := work.Print.print_newline(clk,eclat_unit);
          \$v4511\ := \$ram_lock\;
          if \$v4511\(0) = '1' then
            state_var5924 := Q_WAIT4510;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(\$19838_copy_root_in_ram6634340_arg\(32 to 47)));
            \$ram_write\ <= \$19851_hd\; \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4509;
          end if;
        when PAUSE_GET4516 =>
          \$19850_w\ := \$ram_value\;
          release(\$ram_lock\);
          \$v4515\ := eclat_if(work.Bool.lnot(""&\$19850_w\(31)) & eclat_if(
                                                                   work.Int.le(
                                                                   \$19838_copy_root_in_ram6634340_arg\(64 to 79), eclat_resize(\$19850_w\(0 to 30),16)) & 
                                                                   work.Int.lt(
                                                                   eclat_resize(\$19850_w\(0 to 30),16), 
                                                                   work.Int.add(
                                                                   \$19838_copy_root_in_ram6634340_arg\(64 to 79), X"1770")) & eclat_false) & eclat_false);
          if \$v4515\(0) = '1' then
            \$19845\ := \$19850_w\ & \$19838_copy_root_in_ram6634340_arg\(32 to 47);
            \$v4502\ := \$ram_lock\;
            if \$v4502\(0) = '1' then
              state_var5924 := Q_WAIT4501;
            else
              acquire(\$ram_lock\);
              \$ram_ptr_write\ <= to_integer(unsigned(\$19838_copy_root_in_ram6634340_arg\(0 to 15)));
              \$ram_write\ <= \$19845\(0 to 31); \$ram_write_request\ <= '1';
              state_var5924 := PAUSE_SET4500;
            end if;
          else
            \$v4514\ := \$ram_lock\;
            if \$v4514\(0) = '1' then
              state_var5924 := Q_WAIT4513;
            else
              acquire(\$ram_lock\);
              \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$19844\(0 to 30),16)));
              state_var5924 := PAUSE_GET4512;
            end if;
          end if;
        when PAUSE_GET4520 =>
          \$19844\ := \$ram_value\;
          release(\$ram_lock\);
          \$v4519\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$19844\(31)) & 
                                     eclat_if(work.Int.le(\$19838_copy_root_in_ram6634340_arg\(48 to 63), eclat_resize(\$19844\(0 to 30),16)) & 
                                     work.Int.lt(eclat_resize(\$19844\(0 to 30),16), 
                                                 work.Int.add(\$19838_copy_root_in_ram6634340_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false));
          if \$v4519\(0) = '1' then
            \$19845\ := \$19844\ & \$19838_copy_root_in_ram6634340_arg\(32 to 47);
            \$v4502\ := \$ram_lock\;
            if \$v4502\(0) = '1' then
              state_var5924 := Q_WAIT4501;
            else
              acquire(\$ram_lock\);
              \$ram_ptr_write\ <= to_integer(unsigned(\$19838_copy_root_in_ram6634340_arg\(0 to 15)));
              \$ram_write\ <= \$19845\(0 to 31); \$ram_write_request\ <= '1';
              state_var5924 := PAUSE_SET4500;
            end if;
          else
            \$v4518\ := \$ram_lock\;
            if \$v4518\(0) = '1' then
              state_var5924 := Q_WAIT4517;
            else
              acquire(\$ram_lock\);
              \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19844\(0 to 30),16), X"000" & X"1")));
              state_var5924 := PAUSE_GET4516;
            end if;
          end if;
        when PAUSE_GET4533 =>
          \$19866_hd\ := \$ram_value\;
          release(\$ram_lock\);
          \$19867\ := work.Print.print_string(clk,of_string("bloc "));
          \$19868\ := work.Int.print(clk,eclat_resize(\$18439_wait662_arg\(33 to 63),16));
          \$19869\ := work.Print.print_string(clk,of_string(" of size "));
          \$19870\ := work.Int.print(clk,work.Int.add(eclat_resize(work.Int.lsr(
                                                                   \$19866_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
          \$19871\ := work.Print.print_string(clk,of_string(" from "));
          \$19872\ := work.Int.print(clk,eclat_resize(\$18439_wait662_arg\(33 to 63),16));
          \$19873\ := work.Print.print_string(clk,of_string(" to "));
          \$19874\ := work.Int.print(clk,\$19787\(32 to 47));
          \$19875\ := work.Print.print_newline(clk,eclat_unit);
          \$v4532\ := \$ram_lock\;
          if \$v4532\(0) = '1' then
            state_var5924 := Q_WAIT4531;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(\$19787\(32 to 47)));
            \$ram_write\ <= \$19866_hd\; \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4530;
          end if;
        when PAUSE_GET4537 =>
          \$19865_w\ := \$ram_value\;
          release(\$ram_lock\);
          \$v4536\ := eclat_if(work.Bool.lnot(""&\$19865_w\(31)) & eclat_if(
                                                                   work.Int.le(
                                                                   \$19778\(112 to 127), eclat_resize(\$19865_w\(0 to 30),16)) & 
                                                                   work.Int.lt(
                                                                   eclat_resize(\$19865_w\(0 to 30),16), 
                                                                   work.Int.add(
                                                                   \$19778\(112 to 127), X"1770")) & eclat_false) & eclat_false);
          if \$v4536\(0) = '1' then
            \$19788\ := \$19865_w\ & \$19787\(32 to 47);
            \$19838_copy_root_in_ram6634340_id\ := "000000001001";
            \$19838_copy_root_in_ram6634340_arg\ := X"0" & X"3e8" & \$18439_wait662_arg\(65 to 80) & \$19788\(32 to 47) & \$19778\(96 to 111) & \$19778\(112 to 127);
            state_var5924 := \$19838_COPY_ROOT_IN_RAM6634340\;
          else
            \$v4535\ := \$ram_lock\;
            if \$v4535\(0) = '1' then
              state_var5924 := Q_WAIT4534;
            else
              acquire(\$ram_lock\);
              \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18439_wait662_arg\(33 to 63),16)));
              state_var5924 := PAUSE_GET4533;
            end if;
          end if;
        when PAUSE_GET4550 =>
          \$19881_hd\ := \$ram_value\;
          release(\$ram_lock\);
          \$19882\ := work.Print.print_string(clk,of_string("bloc "));
          \$19883\ := work.Int.print(clk,eclat_resize(\$18439_wait662_arg\(1 to 31),16));
          \$19884\ := work.Print.print_string(clk,of_string(" of size "));
          \$19885\ := work.Int.print(clk,work.Int.add(eclat_resize(work.Int.lsr(
                                                                   \$19881_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
          \$19886\ := work.Print.print_string(clk,of_string(" from "));
          \$19887\ := work.Int.print(clk,eclat_resize(\$18439_wait662_arg\(1 to 31),16));
          \$19888\ := work.Print.print_string(clk,of_string(" to "));
          \$19889\ := work.Int.print(clk,\$19778\(112 to 127));
          \$19890\ := work.Print.print_newline(clk,eclat_unit);
          \$v4549\ := \$ram_lock\;
          if \$v4549\(0) = '1' then
            state_var5924 := Q_WAIT4548;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(\$19778\(112 to 127)));
            \$ram_write\ <= \$19881_hd\; \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4547;
          end if;
        when PAUSE_GET4554 =>
          \$19880_w\ := \$ram_value\;
          release(\$ram_lock\);
          \$v4553\ := eclat_if(work.Bool.lnot(""&\$19880_w\(31)) & eclat_if(
                                                                   work.Int.le(
                                                                   \$19778\(112 to 127), eclat_resize(\$19880_w\(0 to 30),16)) & 
                                                                   work.Int.lt(
                                                                   eclat_resize(\$19880_w\(0 to 30),16), 
                                                                   work.Int.add(
                                                                   \$19778\(112 to 127), X"1770")) & eclat_false) & eclat_false);
          if \$v4553\(0) = '1' then
            \$19787\ := \$19880_w\ & \$19778\(112 to 127);
            \$v4540\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$18439_wait662_arg\(64)) & 
                                       eclat_if(work.Int.le(\$19778\(96 to 111), eclat_resize(\$18439_wait662_arg\(33 to 63),16)) & 
                                       work.Int.lt(eclat_resize(\$18439_wait662_arg\(33 to 63),16), 
                                                   work.Int.add(\$19778\(96 to 111), X"1770")) & eclat_false) & eclat_false));
            if \$v4540\(0) = '1' then
              \$19788\ := \$18439_wait662_arg\(33 to 64) & \$19787\(32 to 47);
              \$19838_copy_root_in_ram6634340_id\ := "000000001001";
              \$19838_copy_root_in_ram6634340_arg\ := X"0" & X"3e8" & \$18439_wait662_arg\(65 to 80) & \$19788\(32 to 47) & \$19778\(96 to 111) & \$19778\(112 to 127);
              state_var5924 := \$19838_COPY_ROOT_IN_RAM6634340\;
            else
              \$v4539\ := \$ram_lock\;
              if \$v4539\(0) = '1' then
                state_var5924 := Q_WAIT4538;
              else
                acquire(\$ram_lock\);
                \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18439_wait662_arg\(33 to 63),16), X"000" & X"1")));
                state_var5924 := PAUSE_GET4537;
              end if;
            end if;
          else
            \$v4552\ := \$ram_lock\;
            if \$v4552\(0) = '1' then
              state_var5924 := Q_WAIT4551;
            else
              acquire(\$ram_lock\);
              \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18439_wait662_arg\(1 to 31),16)));
              state_var5924 := PAUSE_GET4550;
            end if;
          end if;
        when PAUSE_SET4437 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$19927\ := eclat_unit;
          \$19779_loop666_arg\ := work.Int.add(\$19779_loop666_arg\(0 to 15), X"000" & X"1") & \$19779_loop666_arg\(16 to 31) & \$19779_loop666_arg\(32 to 47) & \$19779_loop666_arg\(48 to 63);
          state_var5924 := \$19779_LOOP666\;
        when PAUSE_SET4444 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$19908\ := eclat_unit;
          \$19780_loop665_arg\ := work.Int.add(\$19780_loop665_arg\(0 to 15), X"000" & X"1") & \$19907\(32 to 47) & \$19780_loop665_arg\(32 to 47) & \$19780_loop665_arg\(48 to 63) & \$19780_loop665_arg\(64 to 79) & \$19780_loop665_arg\(80 to 95);
          state_var5924 := \$19780_LOOP665\;
        when PAUSE_SET4447 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$19923\ := eclat_unit;
          \$19907\ := eclat_resize(\$19780_loop665_arg\(16 to 31),31) & eclat_false & 
          work.Int.add(\$19780_loop665_arg\(16 to 31), work.Int.add(eclat_resize(
                                                                    work.Int.lsr(
                                                                    \$19910_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
          \$v4446\ := \$ram_lock\;
          if \$v4446\(0) = '1' then
            state_var5924 := Q_WAIT4445;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(\$19780_loop665_arg\(64 to 79), \$19780_loop665_arg\(0 to 15))));
            \$ram_write\ <= \$19907\(0 to 31); \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4444;
          end if;
        when PAUSE_SET4450 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$19922\ := eclat_unit;
          \$v4449\ := \$ram_lock\;
          if \$v4449\(0) = '1' then
            state_var5924 := Q_WAIT4448;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19906\(0 to 30),16), X"000" & X"1")));
            \$ram_write\ <= eclat_resize(\$19780_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4447;
          end if;
        when PAUSE_SET4453 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$19920\ := eclat_unit;
          \$19779_loop666_id\ := "000000000010";
          \$19779_loop666_arg\ := X"000" & X"1" & \$19780_loop665_arg\(16 to 31) & eclat_resize(\$19906\(0 to 30),16) & eclat_resize(
          work.Int.lsr(\$19910_hd\(0 to 30), X"0000000" & X"2"),16);
          state_var5924 := \$19779_LOOP666\;
        when PAUSE_SET4473 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$19819\ := eclat_unit;
          \$19820\ := work.Print.print_string(clk,of_string(" next="));
          \$19821\ := work.Int.print(clk,\$19818\(32 to 47));
          \$19822\ := work.Print.print_newline(clk,eclat_unit);
          \$19811_copy_root_in_ram6634341_arg\ := work.Int.add(\$19811_copy_root_in_ram6634341_arg\(0 to 15), X"000" & X"1") & \$19811_copy_root_in_ram6634341_arg\(16 to 31) & \$19818\(32 to 47) & \$19811_copy_root_in_ram6634341_arg\(48 to 63) & \$19811_copy_root_in_ram6634341_arg\(64 to 79);
          state_var5924 := \$19811_COPY_ROOT_IN_RAM6634341\;
        when PAUSE_SET4476 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$19837\ := eclat_unit;
          \$19818\ := eclat_resize(\$19811_copy_root_in_ram6634341_arg\(32 to 47),31) & eclat_false & 
          work.Int.add(\$19811_copy_root_in_ram6634341_arg\(32 to 47), 
                       work.Int.add(eclat_resize(work.Int.lsr(\$19824_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
          \$v4475\ := \$ram_lock\;
          if \$v4475\(0) = '1' then
            state_var5924 := Q_WAIT4474;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(\$19811_copy_root_in_ram6634341_arg\(0 to 15)));
            \$ram_write\ <= \$19818\(0 to 31); \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4473;
          end if;
        when PAUSE_SET4479 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$19836\ := eclat_unit;
          \$v4478\ := \$ram_lock\;
          if \$v4478\(0) = '1' then
            state_var5924 := Q_WAIT4477;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19817\(0 to 30),16), X"000" & X"1")));
            \$ram_write\ <= eclat_resize(\$19811_copy_root_in_ram6634341_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4476;
          end if;
        when PAUSE_SET4482 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$19834\ := eclat_unit;
          \$19779_loop666_id\ := "000000000110";
          \$19779_loop666_arg\ := X"000" & X"1" & \$19811_copy_root_in_ram6634341_arg\(32 to 47) & eclat_resize(\$19817\(0 to 30),16) & eclat_resize(
          work.Int.lsr(\$19824_hd\(0 to 30), X"0000000" & X"2"),16);
          state_var5924 := \$19779_LOOP666\;
        when PAUSE_SET4500 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$19846\ := eclat_unit;
          \$19847\ := work.Print.print_string(clk,of_string(" next="));
          \$19848\ := work.Int.print(clk,\$19845\(32 to 47));
          \$19849\ := work.Print.print_newline(clk,eclat_unit);
          \$19838_copy_root_in_ram6634340_arg\ := work.Int.add(\$19838_copy_root_in_ram6634340_arg\(0 to 15), X"000" & X"1") & \$19838_copy_root_in_ram6634340_arg\(16 to 31) & \$19845\(32 to 47) & \$19838_copy_root_in_ram6634340_arg\(48 to 63) & \$19838_copy_root_in_ram6634340_arg\(64 to 79);
          state_var5924 := \$19838_COPY_ROOT_IN_RAM6634340\;
        when PAUSE_SET4503 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$19864\ := eclat_unit;
          \$19845\ := eclat_resize(\$19838_copy_root_in_ram6634340_arg\(32 to 47),31) & eclat_false & 
          work.Int.add(\$19838_copy_root_in_ram6634340_arg\(32 to 47), 
                       work.Int.add(eclat_resize(work.Int.lsr(\$19851_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
          \$v4502\ := \$ram_lock\;
          if \$v4502\(0) = '1' then
            state_var5924 := Q_WAIT4501;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(\$19838_copy_root_in_ram6634340_arg\(0 to 15)));
            \$ram_write\ <= \$19845\(0 to 31); \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4500;
          end if;
        when PAUSE_SET4506 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$19863\ := eclat_unit;
          \$v4505\ := \$ram_lock\;
          if \$v4505\(0) = '1' then
            state_var5924 := Q_WAIT4504;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19844\(0 to 30),16), X"000" & X"1")));
            \$ram_write\ <= eclat_resize(\$19838_copy_root_in_ram6634340_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4503;
          end if;
        when PAUSE_SET4509 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$19861\ := eclat_unit;
          \$19779_loop666_id\ := "000000001000";
          \$19779_loop666_arg\ := X"000" & X"1" & \$19838_copy_root_in_ram6634340_arg\(32 to 47) & eclat_resize(\$19844\(0 to 30),16) & eclat_resize(
          work.Int.lsr(\$19851_hd\(0 to 30), X"0000000" & X"2"),16);
          state_var5924 := \$19779_LOOP666\;
        when PAUSE_SET4524 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$19879\ := eclat_unit;
          \$19788\ := eclat_resize(\$19787\(32 to 47),31) & eclat_false & 
          work.Int.add(\$19787\(32 to 47), work.Int.add(eclat_resize(
                                                        work.Int.lsr(
                                                        \$19866_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
          \$19838_copy_root_in_ram6634340_id\ := "000000001001";
          \$19838_copy_root_in_ram6634340_arg\ := X"0" & X"3e8" & \$18439_wait662_arg\(65 to 80) & \$19788\(32 to 47) & \$19778\(96 to 111) & \$19778\(112 to 127);
          state_var5924 := \$19838_COPY_ROOT_IN_RAM6634340\;
        when PAUSE_SET4527 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$19878\ := eclat_unit;
          \$v4526\ := \$ram_lock\;
          if \$v4526\(0) = '1' then
            state_var5924 := Q_WAIT4525;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18439_wait662_arg\(33 to 63),16), X"000" & X"1")));
            \$ram_write\ <= eclat_resize(\$19787\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4524;
          end if;
        when PAUSE_SET4530 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$19876\ := eclat_unit;
          \$19779_loop666_id\ := "000000001010";
          \$19779_loop666_arg\ := X"000" & X"1" & \$19787\(32 to 47) & eclat_resize(\$18439_wait662_arg\(33 to 63),16) & eclat_resize(
          work.Int.lsr(\$19866_hd\(0 to 30), X"0000000" & X"2"),16);
          state_var5924 := \$19779_LOOP666\;
        when PAUSE_SET4541 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$19894\ := eclat_unit;
          \$19787\ := eclat_resize(\$19778\(112 to 127),31) & eclat_false & 
          work.Int.add(\$19778\(112 to 127), work.Int.add(eclat_resize(
                                                          work.Int.lsr(
                                                          \$19881_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
          \$v4540\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$18439_wait662_arg\(64)) & 
                                     eclat_if(work.Int.le(\$19778\(96 to 111), eclat_resize(\$18439_wait662_arg\(33 to 63),16)) & 
                                     work.Int.lt(eclat_resize(\$18439_wait662_arg\(33 to 63),16), 
                                                 work.Int.add(\$19778\(96 to 111), X"1770")) & eclat_false) & eclat_false));
          if \$v4540\(0) = '1' then
            \$19788\ := \$18439_wait662_arg\(33 to 64) & \$19787\(32 to 47);
            \$19838_copy_root_in_ram6634340_id\ := "000000001001";
            \$19838_copy_root_in_ram6634340_arg\ := X"0" & X"3e8" & \$18439_wait662_arg\(65 to 80) & \$19788\(32 to 47) & \$19778\(96 to 111) & \$19778\(112 to 127);
            state_var5924 := \$19838_COPY_ROOT_IN_RAM6634340\;
          else
            \$v4539\ := \$ram_lock\;
            if \$v4539\(0) = '1' then
              state_var5924 := Q_WAIT4538;
            else
              acquire(\$ram_lock\);
              \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18439_wait662_arg\(33 to 63),16), X"000" & X"1")));
              state_var5924 := PAUSE_GET4537;
            end if;
          end if;
        when PAUSE_SET4544 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$19893\ := eclat_unit;
          \$v4543\ := \$ram_lock\;
          if \$v4543\(0) = '1' then
            state_var5924 := Q_WAIT4542;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18439_wait662_arg\(1 to 31),16), X"000" & X"1")));
            \$ram_write\ <= eclat_resize(\$19778\(112 to 127),31) & eclat_false; \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4541;
          end if;
        when PAUSE_SET4547 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$19891\ := eclat_unit;
          \$19779_loop666_id\ := "000000001011";
          \$19779_loop666_arg\ := X"000" & X"1" & \$19778\(112 to 127) & eclat_resize(\$18439_wait662_arg\(1 to 31),16) & eclat_resize(
          work.Int.lsr(\$19881_hd\(0 to 30), X"0000000" & X"2"),16);
          state_var5924 := \$19779_LOOP666\;
        when Q_WAIT4438 =>
          \$v4439\ := \$ram_lock\;
          if \$v4439\(0) = '1' then
            state_var5924 := Q_WAIT4438;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(\$19779_loop666_arg\(16 to 31), \$19779_loop666_arg\(0 to 15))));
            \$ram_write\ <= \$19926\; \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4437;
          end if;
        when Q_WAIT4441 =>
          \$v4442\ := \$ram_lock\;
          if \$v4442\(0) = '1' then
            state_var5924 := Q_WAIT4441;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$19779_loop666_arg\(32 to 47), \$19779_loop666_arg\(0 to 15))));
            state_var5924 := PAUSE_GET4440;
          end if;
        when Q_WAIT4445 =>
          \$v4446\ := \$ram_lock\;
          if \$v4446\(0) = '1' then
            state_var5924 := Q_WAIT4445;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(\$19780_loop665_arg\(64 to 79), \$19780_loop665_arg\(0 to 15))));
            \$ram_write\ <= \$19907\(0 to 31); \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4444;
          end if;
        when Q_WAIT4448 =>
          \$v4449\ := \$ram_lock\;
          if \$v4449\(0) = '1' then
            state_var5924 := Q_WAIT4448;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19906\(0 to 30),16), X"000" & X"1")));
            \$ram_write\ <= eclat_resize(\$19780_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4447;
          end if;
        when Q_WAIT4451 =>
          \$v4452\ := \$ram_lock\;
          if \$v4452\(0) = '1' then
            state_var5924 := Q_WAIT4451;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$19906\(0 to 30),16)));
            \$ram_write\ <= eclat_resize(\$19780_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4450;
          end if;
        when Q_WAIT4454 =>
          \$v4455\ := \$ram_lock\;
          if \$v4455\(0) = '1' then
            state_var5924 := Q_WAIT4454;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(\$19780_loop665_arg\(16 to 31)));
            \$ram_write\ <= \$19910_hd\; \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4453;
          end if;
        when Q_WAIT4457 =>
          \$v4458\ := \$ram_lock\;
          if \$v4458\(0) = '1' then
            state_var5924 := Q_WAIT4457;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$19906\(0 to 30),16)));
            state_var5924 := PAUSE_GET4456;
          end if;
        when Q_WAIT4461 =>
          \$v4462\ := \$ram_lock\;
          if \$v4462\(0) = '1' then
            state_var5924 := Q_WAIT4461;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19906\(0 to 30),16), X"000" & X"1")));
            state_var5924 := PAUSE_GET4460;
          end if;
        when Q_WAIT4465 =>
          \$v4466\ := \$ram_lock\;
          if \$v4466\(0) = '1' then
            state_var5924 := Q_WAIT4465;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$19780_loop665_arg\(64 to 79), \$19780_loop665_arg\(0 to 15))));
            state_var5924 := PAUSE_GET4464;
          end if;
        when Q_WAIT4469 =>
          \$v4470\ := \$ram_lock\;
          if \$v4470\(0) = '1' then
            state_var5924 := Q_WAIT4469;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(\$19781_aux664_arg\(0 to 15)));
            state_var5924 := PAUSE_GET4468;
          end if;
        when Q_WAIT4474 =>
          \$v4475\ := \$ram_lock\;
          if \$v4475\(0) = '1' then
            state_var5924 := Q_WAIT4474;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(\$19811_copy_root_in_ram6634341_arg\(0 to 15)));
            \$ram_write\ <= \$19818\(0 to 31); \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4473;
          end if;
        when Q_WAIT4477 =>
          \$v4478\ := \$ram_lock\;
          if \$v4478\(0) = '1' then
            state_var5924 := Q_WAIT4477;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19817\(0 to 30),16), X"000" & X"1")));
            \$ram_write\ <= eclat_resize(\$19811_copy_root_in_ram6634341_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4476;
          end if;
        when Q_WAIT4480 =>
          \$v4481\ := \$ram_lock\;
          if \$v4481\(0) = '1' then
            state_var5924 := Q_WAIT4480;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$19817\(0 to 30),16)));
            \$ram_write\ <= eclat_resize(\$19811_copy_root_in_ram6634341_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4479;
          end if;
        when Q_WAIT4483 =>
          \$v4484\ := \$ram_lock\;
          if \$v4484\(0) = '1' then
            state_var5924 := Q_WAIT4483;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(\$19811_copy_root_in_ram6634341_arg\(32 to 47)));
            \$ram_write\ <= \$19824_hd\; \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4482;
          end if;
        when Q_WAIT4486 =>
          \$v4487\ := \$ram_lock\;
          if \$v4487\(0) = '1' then
            state_var5924 := Q_WAIT4486;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$19817\(0 to 30),16)));
            state_var5924 := PAUSE_GET4485;
          end if;
        when Q_WAIT4490 =>
          \$v4491\ := \$ram_lock\;
          if \$v4491\(0) = '1' then
            state_var5924 := Q_WAIT4490;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19817\(0 to 30),16), X"000" & X"1")));
            state_var5924 := PAUSE_GET4489;
          end if;
        when Q_WAIT4494 =>
          \$v4495\ := \$ram_lock\;
          if \$v4495\(0) = '1' then
            state_var5924 := Q_WAIT4494;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(\$19811_copy_root_in_ram6634341_arg\(0 to 15)));
            state_var5924 := PAUSE_GET4493;
          end if;
        when Q_WAIT4498 =>
          \$v4499\ := \$global_end_lock\;
          if \$v4499\(0) = '1' then
            state_var5924 := Q_WAIT4498;
          else
            acquire(\$global_end_lock\);
            \$global_end_ptr\ <= 0;
            state_var5924 := PAUSE_GET4497;
          end if;
        when Q_WAIT4501 =>
          \$v4502\ := \$ram_lock\;
          if \$v4502\(0) = '1' then
            state_var5924 := Q_WAIT4501;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(\$19838_copy_root_in_ram6634340_arg\(0 to 15)));
            \$ram_write\ <= \$19845\(0 to 31); \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4500;
          end if;
        when Q_WAIT4504 =>
          \$v4505\ := \$ram_lock\;
          if \$v4505\(0) = '1' then
            state_var5924 := Q_WAIT4504;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19844\(0 to 30),16), X"000" & X"1")));
            \$ram_write\ <= eclat_resize(\$19838_copy_root_in_ram6634340_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4503;
          end if;
        when Q_WAIT4507 =>
          \$v4508\ := \$ram_lock\;
          if \$v4508\(0) = '1' then
            state_var5924 := Q_WAIT4507;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$19844\(0 to 30),16)));
            \$ram_write\ <= eclat_resize(\$19838_copy_root_in_ram6634340_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4506;
          end if;
        when Q_WAIT4510 =>
          \$v4511\ := \$ram_lock\;
          if \$v4511\(0) = '1' then
            state_var5924 := Q_WAIT4510;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(\$19838_copy_root_in_ram6634340_arg\(32 to 47)));
            \$ram_write\ <= \$19851_hd\; \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4509;
          end if;
        when Q_WAIT4513 =>
          \$v4514\ := \$ram_lock\;
          if \$v4514\(0) = '1' then
            state_var5924 := Q_WAIT4513;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$19844\(0 to 30),16)));
            state_var5924 := PAUSE_GET4512;
          end if;
        when Q_WAIT4517 =>
          \$v4518\ := \$ram_lock\;
          if \$v4518\(0) = '1' then
            state_var5924 := Q_WAIT4517;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19844\(0 to 30),16), X"000" & X"1")));
            state_var5924 := PAUSE_GET4516;
          end if;
        when Q_WAIT4521 =>
          \$v4522\ := \$ram_lock\;
          if \$v4522\(0) = '1' then
            state_var5924 := Q_WAIT4521;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(\$19838_copy_root_in_ram6634340_arg\(0 to 15)));
            state_var5924 := PAUSE_GET4520;
          end if;
        when Q_WAIT4525 =>
          \$v4526\ := \$ram_lock\;
          if \$v4526\(0) = '1' then
            state_var5924 := Q_WAIT4525;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18439_wait662_arg\(33 to 63),16), X"000" & X"1")));
            \$ram_write\ <= eclat_resize(\$19787\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4524;
          end if;
        when Q_WAIT4528 =>
          \$v4529\ := \$ram_lock\;
          if \$v4529\(0) = '1' then
            state_var5924 := Q_WAIT4528;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18439_wait662_arg\(33 to 63),16)));
            \$ram_write\ <= eclat_resize(\$19787\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4527;
          end if;
        when Q_WAIT4531 =>
          \$v4532\ := \$ram_lock\;
          if \$v4532\(0) = '1' then
            state_var5924 := Q_WAIT4531;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(\$19787\(32 to 47)));
            \$ram_write\ <= \$19866_hd\; \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4530;
          end if;
        when Q_WAIT4534 =>
          \$v4535\ := \$ram_lock\;
          if \$v4535\(0) = '1' then
            state_var5924 := Q_WAIT4534;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18439_wait662_arg\(33 to 63),16)));
            state_var5924 := PAUSE_GET4533;
          end if;
        when Q_WAIT4538 =>
          \$v4539\ := \$ram_lock\;
          if \$v4539\(0) = '1' then
            state_var5924 := Q_WAIT4538;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18439_wait662_arg\(33 to 63),16), X"000" & X"1")));
            state_var5924 := PAUSE_GET4537;
          end if;
        when Q_WAIT4542 =>
          \$v4543\ := \$ram_lock\;
          if \$v4543\(0) = '1' then
            state_var5924 := Q_WAIT4542;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18439_wait662_arg\(1 to 31),16), X"000" & X"1")));
            \$ram_write\ <= eclat_resize(\$19778\(112 to 127),31) & eclat_false; \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4541;
          end if;
        when Q_WAIT4545 =>
          \$v4546\ := \$ram_lock\;
          if \$v4546\(0) = '1' then
            state_var5924 := Q_WAIT4545;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18439_wait662_arg\(1 to 31),16)));
            \$ram_write\ <= eclat_resize(\$19778\(112 to 127),31) & eclat_false; \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4544;
          end if;
        when Q_WAIT4548 =>
          \$v4549\ := \$ram_lock\;
          if \$v4549\(0) = '1' then
            state_var5924 := Q_WAIT4548;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(\$19778\(112 to 127)));
            \$ram_write\ <= \$19881_hd\; \$ram_write_request\ <= '1';
            state_var5924 := PAUSE_SET4547;
          end if;
        when Q_WAIT4551 =>
          \$v4552\ := \$ram_lock\;
          if \$v4552\(0) = '1' then
            state_var5924 := Q_WAIT4551;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18439_wait662_arg\(1 to 31),16)));
            state_var5924 := PAUSE_GET4550;
          end if;
        when Q_WAIT4555 =>
          \$v4556\ := \$ram_lock\;
          if \$v4556\(0) = '1' then
            state_var5924 := Q_WAIT4555;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18439_wait662_arg\(1 to 31),16), X"000" & X"1")));
            state_var5924 := PAUSE_GET4554;
          end if;
        when IDLE4436 =>
          rdy4435 := eclat_false;
          \$v4558\ := work.Int.gt(work.Int.add(\$19778\(80 to 95), \$18439_wait662_arg\(81 to 96)), 
                                  work.Int.add(\$19778\(96 to 111), X"1770"));
          if \$v4558\(0) = '1' then
            \$19782\ := work.Print.print_newline(clk,eclat_unit);
            \$19783\ := work.Print.print_newline(clk,eclat_unit);
            \$19784\ := work.Print.print_string(clk,of_string("[================= GC START ======================]"));
            \$19785\ := work.Print.print_newline(clk,eclat_unit);
            \$19786\ := work.Print.print_newline(clk,eclat_unit);
            \$v4557\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$18439_wait662_arg\(32)) & 
                                       eclat_if(work.Int.le(\$19778\(96 to 111), eclat_resize(\$18439_wait662_arg\(1 to 31),16)) & 
                                       work.Int.lt(eclat_resize(\$18439_wait662_arg\(1 to 31),16), 
                                                   work.Int.add(\$19778\(96 to 111), X"1770")) & eclat_false) & eclat_false));
            if \$v4557\(0) = '1' then
              \$19787\ := \$18439_wait662_arg\(1 to 32) & \$19778\(112 to 127);
              \$v4540\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$18439_wait662_arg\(64)) & 
                                         eclat_if(work.Int.le(\$19778\(96 to 111), eclat_resize(\$18439_wait662_arg\(33 to 63),16)) & 
                                         work.Int.lt(eclat_resize(\$18439_wait662_arg\(33 to 63),16), 
                                                     work.Int.add(\$19778\(96 to 111), X"1770")) & eclat_false) & eclat_false));
              if \$v4540\(0) = '1' then
                \$19788\ := \$18439_wait662_arg\(33 to 64) & \$19787\(32 to 47);
                \$19838_copy_root_in_ram6634340_id\ := "000000001001";
                \$19838_copy_root_in_ram6634340_arg\ := X"0" & X"3e8" & \$18439_wait662_arg\(65 to 80) & \$19788\(32 to 47) & \$19778\(96 to 111) & \$19778\(112 to 127);
                state_var5924 := \$19838_COPY_ROOT_IN_RAM6634340\;
              else
                \$v4539\ := \$ram_lock\;
                if \$v4539\(0) = '1' then
                  state_var5924 := Q_WAIT4538;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18439_wait662_arg\(33 to 63),16), X"000" & X"1")));
                  state_var5924 := PAUSE_GET4537;
                end if;
              end if;
            else
              \$v4556\ := \$ram_lock\;
              if \$v4556\(0) = '1' then
                state_var5924 := Q_WAIT4555;
              else
                acquire(\$ram_lock\);
                \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18439_wait662_arg\(1 to 31),16), X"000" & X"1")));
                state_var5924 := PAUSE_GET4554;
              end if;
            end if;
          else
            result4434 := \$18439_wait662_arg\(1 to 32) & \$18439_wait662_arg\(33 to 64) & \$19778\(80 to 95) & 
            work.Int.add(\$19778\(80 to 95), \$18439_wait662_arg\(81 to 96)) & \$19778\(96 to 111) & \$19778\(112 to 127);
            rdy4435 := eclat_true;
            state_var5924 := IDLE4436;
          end if;
        end case;
        
        if rdy4435(0) = '1' then
          
        else
          result4434 := \$19778\(0 to 31) & \$19778\(32 to 63) & \$19778\(64 to 79) & \$19778\(80 to 95) & \$19778\(96 to 111) & \$19778\(112 to 127);
        end if;
        \$19778\ := result4434 & rdy4435;
        \$19777\ := \$19778\;
        \$v4433\ := ""&\$19777\(128);
        if \$v4433\(0) = '1' then
          \$18439_wait662_result\ := \$19777\(0 to 31) & \$19777\(32 to 63) & \$19777\(64 to 79);
          \$19770\ := \$18439_wait662_result\;
          \$19771\ := work.Print.print_string(clk,of_string("size:"));
          \$19772\ := work.Int.print(clk,eclat_if(work.Int.eq(\$18440_make_block579_arg\(112 to 127), X"000" & X"0") & X"000" & X"1" & \$18440_make_block579_arg\(112 to 127)));
          \$19773\ := work.Print.print_newline(clk,eclat_unit);
          \$v4562\ := \$ram_lock\;
          if \$v4562\(0) = '1' then
            state := Q_WAIT4561;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(\$19770\(64 to 79)));
            \$ram_write\ <= work.Int.lor(work.Int.lsl(eclat_resize(\$18440_make_block579_arg\(80 to 111),31), X"000000" & X"18"), 
                                         work.Int.lsl(eclat_resize(eclat_if(
                                                                   work.Int.eq(
                                                                   \$18440_make_block579_arg\(112 to 127), X"000" & X"0") & X"000" & X"1" & \$18440_make_block579_arg\(112 to 127)),31), X"0000000" & X"2")) & eclat_true; \$ram_write_request\ <= '1';
            state := PAUSE_SET4560;
          end if;
        else
          \$18439_wait662_arg\ := eclat_unit & \$18439_wait662_arg\(1 to 32) & \$18439_wait662_arg\(33 to 64) & \$18439_wait662_arg\(65 to 80) & \$18439_wait662_arg\(81 to 96);
          state := \$18439_WAIT662\;
        end if;
      when \$18440_MAKE_BLOCK579\ =>
        \$19766\ := work.Print.print_string(clk,of_string("GC-ALLOC:(size="));
        \$19767\ := work.Int.print(clk,work.Int.add(eclat_if(work.Int.eq(
                                                             \$18440_make_block579_arg\(112 to 127), X"000" & X"0") & X"000" & X"1" & \$18440_make_block579_arg\(112 to 127)), X"000" & X"1"));
        \$19768\ := work.Print.print_string(clk,of_string(")"));
        \$19769\ := work.Print.print_newline(clk,eclat_unit);
        \$18439_wait662_id\ := "000000001100";
        \$18439_wait662_arg\ := eclat_unit & \$18440_make_block579_arg\(16 to 47) & \$18440_make_block579_arg\(48 to 79) & \$18440_make_block579_arg\(0 to 15) & 
        work.Int.add(eclat_if(work.Int.eq(\$18440_make_block579_arg\(112 to 127), X"000" & X"0") & X"000" & X"1" & \$18440_make_block579_arg\(112 to 127)), X"000" & X"1");
        state := \$18439_WAIT662\;
      when PAUSE_GET4405 =>
        \$19950\ := \$ram_value\;
        release(\$ram_lock\);
        \$v4404\ := \$ram_lock\;
        if \$v4404\(0) = '1' then
          state := Q_WAIT4403;
        else
          acquire(\$ram_lock\);
          \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(\$18437_loop666_arg\(16 to 31), \$18437_loop666_arg\(0 to 15))));
          \$ram_write\ <= \$19950\; \$ram_write_request\ <= '1';
          state := PAUSE_SET4402;
        end if;
      when PAUSE_GET4421 =>
        \$19934_hd\ := \$ram_value\;
        release(\$ram_lock\);
        \$19935\ := work.Print.print_string(clk,of_string("bloc "));
        \$19936\ := work.Int.print(clk,eclat_resize(\$19930\(0 to 30),16));
        \$19937\ := work.Print.print_string(clk,of_string(" of size "));
        \$19938\ := work.Int.print(clk,work.Int.add(eclat_resize(work.Int.lsr(
                                                                 \$19934_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
        \$19939\ := work.Print.print_string(clk,of_string(" from "));
        \$19940\ := work.Int.print(clk,eclat_resize(\$19930\(0 to 30),16));
        \$19941\ := work.Print.print_string(clk,of_string(" to "));
        \$19942\ := work.Int.print(clk,\$18438_loop665_arg\(16 to 31));
        \$19943\ := work.Print.print_newline(clk,eclat_unit);
        \$v4420\ := \$ram_lock\;
        if \$v4420\(0) = '1' then
          state := Q_WAIT4419;
        else
          acquire(\$ram_lock\);
          \$ram_ptr_write\ <= to_integer(unsigned(\$18438_loop665_arg\(16 to 31)));
          \$ram_write\ <= \$19934_hd\; \$ram_write_request\ <= '1';
          state := PAUSE_SET4418;
        end if;
      when PAUSE_GET4425 =>
        \$19933_w\ := \$ram_value\;
        release(\$ram_lock\);
        \$v4424\ := eclat_if(work.Bool.lnot(""&\$19933_w\(31)) & eclat_if(
                                                                 work.Int.le(
                                                                 \$18438_loop665_arg\(48 to 63), eclat_resize(\$19933_w\(0 to 30),16)) & 
                                                                 work.Int.lt(
                                                                 eclat_resize(\$19933_w\(0 to 30),16), 
                                                                 work.Int.add(
                                                                 \$18438_loop665_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false);
        if \$v4424\(0) = '1' then
          \$19931\ := \$19933_w\ & \$18438_loop665_arg\(16 to 31);
          \$v4411\ := \$ram_lock\;
          if \$v4411\(0) = '1' then
            state := Q_WAIT4410;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(\$18438_loop665_arg\(64 to 79), \$18438_loop665_arg\(0 to 15))));
            \$ram_write\ <= \$19931\(0 to 31); \$ram_write_request\ <= '1';
            state := PAUSE_SET4409;
          end if;
        else
          \$v4423\ := \$ram_lock\;
          if \$v4423\(0) = '1' then
            state := Q_WAIT4422;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$19930\(0 to 30),16)));
            state := PAUSE_GET4421;
          end if;
        end if;
      when PAUSE_GET4429 =>
        \$19930\ := \$ram_value\;
        release(\$ram_lock\);
        \$v4428\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$19930\(31)) & 
                                   eclat_if(work.Int.le(\$18438_loop665_arg\(32 to 47), eclat_resize(\$19930\(0 to 30),16)) & 
                                   work.Int.lt(eclat_resize(\$19930\(0 to 30),16), 
                                               work.Int.add(\$18438_loop665_arg\(32 to 47), X"1770")) & eclat_false) & eclat_false));
        if \$v4428\(0) = '1' then
          \$19931\ := \$19930\ & \$18438_loop665_arg\(16 to 31);
          \$v4411\ := \$ram_lock\;
          if \$v4411\(0) = '1' then
            state := Q_WAIT4410;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(\$18438_loop665_arg\(64 to 79), \$18438_loop665_arg\(0 to 15))));
            \$ram_write\ <= \$19931\(0 to 31); \$ram_write_request\ <= '1';
            state := PAUSE_SET4409;
          end if;
        else
          \$v4427\ := \$ram_lock\;
          if \$v4427\(0) = '1' then
            state := Q_WAIT4426;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19930\(0 to 30),16), X"000" & X"1")));
            state := PAUSE_GET4425;
          end if;
        end if;
      when PAUSE_SET4402 =>
        \$ram_write_request\ <= '0';
        release(\$ram_lock\);
        \$19951\ := eclat_unit;
        \$18437_loop666_arg\ := work.Int.add(\$18437_loop666_arg\(0 to 15), X"000" & X"1") & \$18437_loop666_arg\(16 to 31) & \$18437_loop666_arg\(32 to 47) & \$18437_loop666_arg\(48 to 63);
        state := \$18437_LOOP666\;
      when PAUSE_SET4409 =>
        \$ram_write_request\ <= '0';
        release(\$ram_lock\);
        \$19932\ := eclat_unit;
        \$18438_loop665_arg\ := work.Int.add(\$18438_loop665_arg\(0 to 15), X"000" & X"1") & \$19931\(32 to 47) & \$18438_loop665_arg\(32 to 47) & \$18438_loop665_arg\(48 to 63) & \$18438_loop665_arg\(64 to 79) & \$18438_loop665_arg\(80 to 95);
        state := \$18438_LOOP665\;
      when PAUSE_SET4412 =>
        \$ram_write_request\ <= '0';
        release(\$ram_lock\);
        \$19947\ := eclat_unit;
        \$19931\ := eclat_resize(\$18438_loop665_arg\(16 to 31),31) & eclat_false & 
        work.Int.add(\$18438_loop665_arg\(16 to 31), work.Int.add(eclat_resize(
                                                                  work.Int.lsr(
                                                                  \$19934_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
        \$v4411\ := \$ram_lock\;
        if \$v4411\(0) = '1' then
          state := Q_WAIT4410;
        else
          acquire(\$ram_lock\);
          \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(\$18438_loop665_arg\(64 to 79), \$18438_loop665_arg\(0 to 15))));
          \$ram_write\ <= \$19931\(0 to 31); \$ram_write_request\ <= '1';
          state := PAUSE_SET4409;
        end if;
      when PAUSE_SET4415 =>
        \$ram_write_request\ <= '0';
        release(\$ram_lock\);
        \$19946\ := eclat_unit;
        \$v4414\ := \$ram_lock\;
        if \$v4414\(0) = '1' then
          state := Q_WAIT4413;
        else
          acquire(\$ram_lock\);
          \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19930\(0 to 30),16), X"000" & X"1")));
          \$ram_write\ <= eclat_resize(\$18438_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
          state := PAUSE_SET4412;
        end if;
      when PAUSE_SET4418 =>
        \$ram_write_request\ <= '0';
        release(\$ram_lock\);
        \$19944\ := eclat_unit;
        \$18437_loop666_id\ := "000000000001";
        \$18437_loop666_arg\ := X"000" & X"1" & \$18438_loop665_arg\(16 to 31) & eclat_resize(\$19930\(0 to 30),16) & eclat_resize(
        work.Int.lsr(\$19934_hd\(0 to 30), X"0000000" & X"2"),16);
        state := \$18437_LOOP666\;
      when PAUSE_SET4560 =>
        \$ram_write_request\ <= '0';
        release(\$ram_lock\);
        \$19774\ := eclat_unit;
        \$18440_make_block579_result\ := \$19770\(0 to 31) & \$19770\(32 to 63) & eclat_resize(\$19770\(64 to 79),31) & eclat_false;
        state := \$18440_MAKE_BLOCK579\;
      when Q_WAIT4403 =>
        \$v4404\ := \$ram_lock\;
        if \$v4404\(0) = '1' then
          state := Q_WAIT4403;
        else
          acquire(\$ram_lock\);
          \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(\$18437_loop666_arg\(16 to 31), \$18437_loop666_arg\(0 to 15))));
          \$ram_write\ <= \$19950\; \$ram_write_request\ <= '1';
          state := PAUSE_SET4402;
        end if;
      when Q_WAIT4406 =>
        \$v4407\ := \$ram_lock\;
        if \$v4407\(0) = '1' then
          state := Q_WAIT4406;
        else
          acquire(\$ram_lock\);
          \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$18437_loop666_arg\(32 to 47), \$18437_loop666_arg\(0 to 15))));
          state := PAUSE_GET4405;
        end if;
      when Q_WAIT4410 =>
        \$v4411\ := \$ram_lock\;
        if \$v4411\(0) = '1' then
          state := Q_WAIT4410;
        else
          acquire(\$ram_lock\);
          \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(\$18438_loop665_arg\(64 to 79), \$18438_loop665_arg\(0 to 15))));
          \$ram_write\ <= \$19931\(0 to 31); \$ram_write_request\ <= '1';
          state := PAUSE_SET4409;
        end if;
      when Q_WAIT4413 =>
        \$v4414\ := \$ram_lock\;
        if \$v4414\(0) = '1' then
          state := Q_WAIT4413;
        else
          acquire(\$ram_lock\);
          \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19930\(0 to 30),16), X"000" & X"1")));
          \$ram_write\ <= eclat_resize(\$18438_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
          state := PAUSE_SET4412;
        end if;
      when Q_WAIT4416 =>
        \$v4417\ := \$ram_lock\;
        if \$v4417\(0) = '1' then
          state := Q_WAIT4416;
        else
          acquire(\$ram_lock\);
          \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$19930\(0 to 30),16)));
          \$ram_write\ <= eclat_resize(\$18438_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
          state := PAUSE_SET4415;
        end if;
      when Q_WAIT4419 =>
        \$v4420\ := \$ram_lock\;
        if \$v4420\(0) = '1' then
          state := Q_WAIT4419;
        else
          acquire(\$ram_lock\);
          \$ram_ptr_write\ <= to_integer(unsigned(\$18438_loop665_arg\(16 to 31)));
          \$ram_write\ <= \$19934_hd\; \$ram_write_request\ <= '1';
          state := PAUSE_SET4418;
        end if;
      when Q_WAIT4422 =>
        \$v4423\ := \$ram_lock\;
        if \$v4423\(0) = '1' then
          state := Q_WAIT4422;
        else
          acquire(\$ram_lock\);
          \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$19930\(0 to 30),16)));
          state := PAUSE_GET4421;
        end if;
      when Q_WAIT4426 =>
        \$v4427\ := \$ram_lock\;
        if \$v4427\(0) = '1' then
          state := Q_WAIT4426;
        else
          acquire(\$ram_lock\);
          \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19930\(0 to 30),16), X"000" & X"1")));
          state := PAUSE_GET4425;
        end if;
      when Q_WAIT4430 =>
        \$v4431\ := \$ram_lock\;
        if \$v4431\(0) = '1' then
          state := Q_WAIT4430;
        else
          acquire(\$ram_lock\);
          \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$18438_loop665_arg\(64 to 79), \$18438_loop665_arg\(0 to 15))));
          state := PAUSE_GET4429;
        end if;
      when Q_WAIT4561 =>
        \$v4562\ := \$ram_lock\;
        if \$v4562\(0) = '1' then
          state := Q_WAIT4561;
        else
          acquire(\$ram_lock\);
          \$ram_ptr_write\ <= to_integer(unsigned(\$19770\(64 to 79)));
          \$ram_write\ <= work.Int.lor(work.Int.lsl(eclat_resize(\$18440_make_block579_arg\(80 to 111),31), X"000000" & X"18"), 
                                       work.Int.lsl(eclat_resize(eclat_if(
                                                                 work.Int.eq(
                                                                 \$18440_make_block579_arg\(112 to 127), X"000" & X"0") & X"000" & X"1" & \$18440_make_block579_arg\(112 to 127)),31), X"0000000" & X"2")) & eclat_true; \$ram_write_request\ <= '1';
          state := PAUSE_SET4560;
        end if;
      when IDLE4401 =>
        rdy4400 := eclat_false;
        \$v5919\ := work.Bool.lnot(""&argument(10));
        if \$v5919\(0) = '1' then
          result4399 := ""&argument(11) & ""&argument(11) & ""&argument(11) & ""&argument(11) & ""&argument(11) & ""&argument(11) & ""&argument(11) & ""&argument(11) & ""&argument(11) & ""&argument(11) & "01100011" & "00000011" & "01110001" & "01110001" & "01100001" & "01100001";
          rdy4400 := eclat_true;
          state := IDLE4401;
        else
          if \$v4327\(0) = '1' then
            
          else
            \$v4327\ := eclat_true;
            \$19763\ := X"0000000" & X"0";
          end if;
          \$19763\ := eclat_if(""&argument(11) & X"0000000" & X"0" & 
                      work.Int.add(\$19763\, X"0000000" & X"1"));
          \$18442_cy\ := \$19763\;
          if \$v4328\(0) = '1' then
            
          else
            \$v4328\ := eclat_true;
            \$18462\ := eclat_false & eclat_false & eclat_false & eclat_false;
          end if;
          \$v5918\ := work.Bool.lnot(""&\$18462\(2));
          if \$v5918\(0) = '1' then
            case state_var5922 is
            when \$18466_LOOP666\ =>
              \$v4581\ := work.Int.ge(\$18466_loop666_arg\(0 to 15), 
                                      work.Int.add(\$18466_loop666_arg\(48 to 63), X"000" & X"1"));
              if \$v4581\(0) = '1' then
                \$18466_loop666_result\ := eclat_unit;
                \$18780\ := \$18466_loop666_result\;
                \$v4590\ := \$ram_lock\;
                if \$v4590\(0) = '1' then
                  state_var5922 := Q_WAIT4589;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18765\(0 to 30),16)));
                  \$ram_write\ <= eclat_resize(\$18467_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var5922 := PAUSE_SET4588;
                end if;
              else
                \$v4580\ := \$ram_lock\;
                if \$v4580\(0) = '1' then
                  state_var5922 := Q_WAIT4579;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$18466_loop666_arg\(32 to 47), \$18466_loop666_arg\(0 to 15))));
                  state_var5922 := PAUSE_GET4578;
                end if;
              end if;
            when \$18467_LOOP665\ =>
              \$v4605\ := work.Int.ge(\$18467_loop665_arg\(0 to 15), 
                                      work.Int.add(\$18467_loop665_arg\(80 to 95), X"000" & X"1"));
              if \$v4605\(0) = '1' then
                \$18467_loop665_result\ := \$18467_loop665_arg\(16 to 31);
                state_var5922 := \$18467_LOOP665\;
              else
                \$v4604\ := \$ram_lock\;
                if \$v4604\(0) = '1' then
                  state_var5922 := Q_WAIT4603;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$18467_loop665_arg\(64 to 79), \$18467_loop665_arg\(0 to 15))));
                  state_var5922 := PAUSE_GET4602;
                end if;
              end if;
            when \$18468_WAIT662\ =>
              if \$v4330\(0) = '1' then
                
              else
                \$v4330\ := eclat_true;
                \$18520\ := \$18468_wait662_arg\(1 to 32) & \$18468_wait662_arg\(33 to 64) & X"0" & X"fa0" & X"0" & X"fa0" & X"0" & X"fa0" & 
                work.Int.add(X"0" & X"fa0", X"1770") & eclat_false;
              end if;
              case state_var5923 is
              when \$18521_LOOP666\ =>
                \$v4616\ := work.Int.ge(\$18521_loop666_arg\(0 to 15), 
                                        work.Int.add(\$18521_loop666_arg\(48 to 63), X"000" & X"1"));
                if \$v4616\(0) = '1' then
                  \$18521_loop666_result\ := eclat_unit;
                  \$18756\ := \$18521_loop666_result\;
                  \$v4625\ := \$ram_lock\;
                  if \$v4625\(0) = '1' then
                    state_var5923 := Q_WAIT4624;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18741\(0 to 30),16)));
                    \$ram_write\ <= eclat_resize(\$18522_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var5923 := PAUSE_SET4623;
                  end if;
                else
                  \$v4615\ := \$ram_lock\;
                  if \$v4615\(0) = '1' then
                    state_var5923 := Q_WAIT4614;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$18521_loop666_arg\(32 to 47), \$18521_loop666_arg\(0 to 15))));
                    state_var5923 := PAUSE_GET4613;
                  end if;
                end if;
              when \$18522_LOOP665\ =>
                \$v4640\ := work.Int.ge(\$18522_loop665_arg\(0 to 15), 
                                        work.Int.add(\$18522_loop665_arg\(80 to 95), X"000" & X"1"));
                if \$v4640\(0) = '1' then
                  \$18522_loop665_result\ := \$18522_loop665_arg\(16 to 31);
                  \$18738_next\ := \$18522_loop665_result\;
                  \$18523_aux664_arg\ := work.Int.add(\$18523_aux664_arg\(0 to 15), 
                                                      work.Int.add(eclat_resize(
                                                                   work.Int.lsr(
                                                                   eclat_resize(eclat_resize(\$18737\(0 to 30),16),31), X"0000000" & X"2"),16), X"000" & X"1")) & \$18738_next\ & \$18523_aux664_arg\(32 to 47) & \$18523_aux664_arg\(48 to 63);
                  state_var5923 := \$18523_AUX664\;
                else
                  \$v4639\ := \$ram_lock\;
                  if \$v4639\(0) = '1' then
                    state_var5923 := Q_WAIT4638;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$18522_loop665_arg\(64 to 79), \$18522_loop665_arg\(0 to 15))));
                    state_var5923 := PAUSE_GET4637;
                  end if;
                end if;
              when \$18523_AUX664\ =>
                \$18732\ := work.Print.print_string(clk,of_string("     scan="));
                \$18733\ := work.Int.print(clk,\$18523_aux664_arg\(0 to 15));
                \$18734\ := work.Print.print_string(clk,of_string(" | next="));
                \$18735\ := work.Int.print(clk,\$18523_aux664_arg\(16 to 31));
                \$18736\ := work.Print.print_newline(clk,eclat_unit);
                \$v4644\ := work.Int.ge(\$18523_aux664_arg\(0 to 15), \$18523_aux664_arg\(16 to 31));
                if \$v4644\(0) = '1' then
                  \$18523_aux664_result\ := \$18523_aux664_arg\(16 to 31);
                  state_var5923 := \$18523_AUX664\;
                else
                  \$v4643\ := \$ram_lock\;
                  if \$v4643\(0) = '1' then
                    state_var5923 := Q_WAIT4642;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(\$18523_aux664_arg\(0 to 15)));
                    state_var5923 := PAUSE_GET4641;
                  end if;
                end if;
              when \$18524_LOOP666\ =>
                \$v4651\ := work.Int.ge(\$18524_loop666_arg\(0 to 15), 
                                        work.Int.add(\$18524_loop666_arg\(48 to 63), X"000" & X"1"));
                if \$v4651\(0) = '1' then
                  \$18524_loop666_result\ := eclat_unit;
                  case \$18524_loop666_id\ is
                  when "000000010000" =>
                    \$18723\ := \$18524_loop666_result\;
                    \$v4660\ := \$ram_lock\;
                    if \$v4660\(0) = '1' then
                      state_var5923 := Q_WAIT4659;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18708\(0 to 30),16)));
                      \$ram_write\ <= eclat_resize(\$18525_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                      state_var5923 := PAUSE_SET4658;
                    end if;
                  when "000000010101" =>
                    \$18595\ := \$18524_loop666_result\;
                    \$v4689\ := \$ram_lock\;
                    if \$v4689\(0) = '1' then
                      state_var5923 := Q_WAIT4688;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18577\(0 to 30),16)));
                      \$ram_write\ <= eclat_resize(\$18571_copy_root_in_ram6634345_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                      state_var5923 := PAUSE_SET4687;
                    end if;
                  when "000000010111" =>
                    \$18610\ := \$18524_loop666_result\;
                    \$v4713\ := \$ram_lock\;
                    if \$v4713\(0) = '1' then
                      state_var5923 := Q_WAIT4712;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18565\(0 to 30),16)));
                      \$ram_write\ <= eclat_resize(\$18559_copy_root_in_ram6634347_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                      state_var5923 := PAUSE_SET4711;
                    end if;
                  when "000000011001" =>
                    \$18649\ := \$18524_loop666_result\;
                    \$v4740\ := \$ram_lock\;
                    if \$v4740\(0) = '1' then
                      state_var5923 := Q_WAIT4739;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18631\(0 to 30),16)));
                      \$ram_write\ <= eclat_resize(\$18625_copy_root_in_ram6634345_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                      state_var5923 := PAUSE_SET4738;
                    end if;
                  when "000000011011" =>
                    \$18664\ := \$18524_loop666_result\;
                    \$v4764\ := \$ram_lock\;
                    if \$v4764\(0) = '1' then
                      state_var5923 := Q_WAIT4763;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18619\(0 to 30),16)));
                      \$ram_write\ <= eclat_resize(\$18613_copy_root_in_ram6634346_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                      state_var5923 := PAUSE_SET4762;
                    end if;
                  when "000000011101" =>
                    \$18679\ := \$18524_loop666_result\;
                    \$v4785\ := \$ram_lock\;
                    if \$v4785\(0) = '1' then
                      state_var5923 := Q_WAIT4784;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18468_wait662_arg\(33 to 63),16)));
                      \$ram_write\ <= eclat_resize(\$18532\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                      state_var5923 := PAUSE_SET4783;
                    end if;
                  when "000000011110" =>
                    \$18694\ := \$18524_loop666_result\;
                    \$v4802\ := \$ram_lock\;
                    if \$v4802\(0) = '1' then
                      state_var5923 := Q_WAIT4801;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18468_wait662_arg\(1 to 31),16)));
                      \$ram_write\ <= eclat_resize(\$18520\(112 to 127),31) & eclat_false; \$ram_write_request\ <= '1';
                      state_var5923 := PAUSE_SET4800;
                    end if;
                  when others =>
                    
                  end case;
                else
                  \$v4650\ := \$ram_lock\;
                  if \$v4650\(0) = '1' then
                    state_var5923 := Q_WAIT4649;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$18524_loop666_arg\(32 to 47), \$18524_loop666_arg\(0 to 15))));
                    state_var5923 := PAUSE_GET4648;
                  end if;
                end if;
              when \$18525_LOOP665\ =>
                \$v4675\ := work.Int.ge(\$18525_loop665_arg\(0 to 15), 
                                        work.Int.add(\$18525_loop665_arg\(80 to 95), X"000" & X"1"));
                if \$v4675\(0) = '1' then
                  \$18525_loop665_result\ := \$18525_loop665_arg\(16 to 31);
                  \$18705_next\ := \$18525_loop665_result\;
                  \$18526_aux664_arg\ := work.Int.add(\$18526_aux664_arg\(0 to 15), 
                                                      work.Int.add(eclat_resize(
                                                                   work.Int.lsr(
                                                                   eclat_resize(eclat_resize(\$18704\(0 to 30),16),31), X"0000000" & X"2"),16), X"000" & X"1")) & \$18705_next\ & \$18526_aux664_arg\(32 to 47) & \$18526_aux664_arg\(48 to 63);
                  state_var5923 := \$18526_AUX664\;
                else
                  \$v4674\ := \$ram_lock\;
                  if \$v4674\(0) = '1' then
                    state_var5923 := Q_WAIT4673;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$18525_loop665_arg\(64 to 79), \$18525_loop665_arg\(0 to 15))));
                    state_var5923 := PAUSE_GET4672;
                  end if;
                end if;
              when \$18526_AUX664\ =>
                \$18699\ := work.Print.print_string(clk,of_string("     scan="));
                \$18700\ := work.Int.print(clk,\$18526_aux664_arg\(0 to 15));
                \$18701\ := work.Print.print_string(clk,of_string(" | next="));
                \$18702\ := work.Int.print(clk,\$18526_aux664_arg\(16 to 31));
                \$18703\ := work.Print.print_newline(clk,eclat_unit);
                \$v4679\ := work.Int.ge(\$18526_aux664_arg\(0 to 15), \$18526_aux664_arg\(16 to 31));
                if \$v4679\(0) = '1' then
                  \$18526_aux664_result\ := \$18526_aux664_arg\(16 to 31);
                  \$18545_next\ := \$18526_aux664_result\;
                  \$18546\ := work.Print.print_string(clk,of_string("memory copied in to_space : "));
                  \$18547\ := work.Int.print(clk,work.Int.sub(\$18545_next\, \$18520\(112 to 127)));
                  \$18548\ := work.Print.print_string(clk,of_string(" words"));
                  \$18549\ := work.Print.print_newline(clk,eclat_unit);
                  \$v4680\ := work.Int.gt(work.Int.sub(\$18545_next\, \$18520\(112 to 127)), X"1770");
                  if \$v4680\(0) = '1' then
                    \$18550\ := work.Print.print_string(clk,of_string("fatal error: "));
                    \$18551\ := work.Print.print_string(clk,of_string("Out of memory"));
                    \$18552\ := work.Print.print_newline(clk,eclat_unit);
                    \$18553_forever6704348_id\ := "000000010011";
                    \$18553_forever6704348_arg\ := eclat_unit;
                    state_var5923 := \$18553_FOREVER6704348\;
                  else
                    \$18535\ := \$18532\(0 to 31) & \$18533\(0 to 31) & \$18545_next\;
                    \$18536\ := work.Print.print_newline(clk,eclat_unit);
                    \$18537\ := work.Print.print_newline(clk,eclat_unit);
                    \$18538\ := work.Print.print_string(clk,of_string("[================= GC END ======================]"));
                    \$18539\ := work.Print.print_newline(clk,eclat_unit);
                    \$18540\ := work.Print.print_newline(clk,eclat_unit);
                    result4607 := \$18535\(0 to 31) & \$18535\(32 to 63) & \$18535\(64 to 79) & 
                    work.Int.add(\$18535\(64 to 79), \$18468_wait662_arg\(81 to 96)) & \$18520\(112 to 127) & \$18520\(96 to 111);
                    rdy4608 := eclat_true;
                    state_var5923 := IDLE4609;
                  end if;
                else
                  \$v4678\ := \$ram_lock\;
                  if \$v4678\(0) = '1' then
                    state_var5923 := Q_WAIT4677;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(\$18526_aux664_arg\(0 to 15)));
                    state_var5923 := PAUSE_GET4676;
                  end if;
                end if;
              when \$18553_FOREVER6704348\ =>
                \$18556_forever6704344_id\ := "000000010010";
                \$18556_forever6704344_arg\ := eclat_unit;
                state_var5923 := \$18556_FOREVER6704344\;
              when \$18556_FOREVER6704344\ =>
                \$18556_forever6704344_arg\ := eclat_unit;
                state_var5923 := \$18556_FOREVER6704344\;
              when \$18559_COPY_ROOT_IN_RAM6634347\ =>
                \$v4728\ := work.Int.ge(\$18559_copy_root_in_ram6634347_arg\(0 to 15), \$18559_copy_root_in_ram6634347_arg\(16 to 31));
                if \$v4728\(0) = '1' then
                  \$18559_copy_root_in_ram6634347_result\ := \$18559_copy_root_in_ram6634347_arg\(32 to 47);
                  \$18542_next\ := \$18559_copy_root_in_ram6634347_result\;
                  \$18543\ := work.Print.print_string(clk,of_string("======================================="));
                  \$18544\ := work.Print.print_newline(clk,eclat_unit);
                  \$18526_aux664_id\ := "000000010100";
                  \$18526_aux664_arg\ := \$18520\(112 to 127) & \$18542_next\ & \$18520\(96 to 111) & \$18520\(112 to 127);
                  state_var5923 := \$18526_AUX664\;
                else
                  \$18562\ := work.Print.print_string(clk,of_string("racine:"));
                  \$18563\ := work.Int.print(clk,\$18559_copy_root_in_ram6634347_arg\(0 to 15));
                  \$18564\ := work.Print.print_newline(clk,eclat_unit);
                  \$v4727\ := \$ram_lock\;
                  if \$v4727\(0) = '1' then
                    state_var5923 := Q_WAIT4726;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(\$18559_copy_root_in_ram6634347_arg\(0 to 15)));
                    state_var5923 := PAUSE_GET4725;
                  end if;
                end if;
              when \$18571_COPY_ROOT_IN_RAM6634345\ =>
                \$v4704\ := work.Int.ge(\$18571_copy_root_in_ram6634345_arg\(0 to 15), \$18571_copy_root_in_ram6634345_arg\(16 to 31));
                if \$v4704\(0) = '1' then
                  \$18571_copy_root_in_ram6634345_result\ := \$18571_copy_root_in_ram6634345_arg\(32 to 47);
                  \$18559_copy_root_in_ram6634347_result\ := \$18571_copy_root_in_ram6634345_result\;
                  \$18542_next\ := \$18559_copy_root_in_ram6634347_result\;
                  \$18543\ := work.Print.print_string(clk,of_string("======================================="));
                  \$18544\ := work.Print.print_newline(clk,eclat_unit);
                  \$18526_aux664_id\ := "000000010100";
                  \$18526_aux664_arg\ := \$18520\(112 to 127) & \$18542_next\ & \$18520\(96 to 111) & \$18520\(112 to 127);
                  state_var5923 := \$18526_AUX664\;
                else
                  \$18574\ := work.Print.print_string(clk,of_string("racine:"));
                  \$18575\ := work.Int.print(clk,\$18571_copy_root_in_ram6634345_arg\(0 to 15));
                  \$18576\ := work.Print.print_newline(clk,eclat_unit);
                  \$v4703\ := \$ram_lock\;
                  if \$v4703\(0) = '1' then
                    state_var5923 := Q_WAIT4702;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(\$18571_copy_root_in_ram6634345_arg\(0 to 15)));
                    state_var5923 := PAUSE_GET4701;
                  end if;
                end if;
              when \$18613_COPY_ROOT_IN_RAM6634346\ =>
                \$v4779\ := work.Int.ge(\$18613_copy_root_in_ram6634346_arg\(0 to 15), \$18613_copy_root_in_ram6634346_arg\(16 to 31));
                if \$v4779\(0) = '1' then
                  \$18613_copy_root_in_ram6634346_result\ := \$18613_copy_root_in_ram6634346_arg\(32 to 47);
                  \$18534_next\ := \$18613_copy_root_in_ram6634346_result\;
                  \$v4731\ := \$global_end_lock\;
                  if \$v4731\(0) = '1' then
                    state_var5923 := Q_WAIT4730;
                  else
                    acquire(\$global_end_lock\);
                    \$global_end_ptr\ <= 0;
                    state_var5923 := PAUSE_GET4729;
                  end if;
                else
                  \$18616\ := work.Print.print_string(clk,of_string("racine:"));
                  \$18617\ := work.Int.print(clk,\$18613_copy_root_in_ram6634346_arg\(0 to 15));
                  \$18618\ := work.Print.print_newline(clk,eclat_unit);
                  \$v4778\ := \$ram_lock\;
                  if \$v4778\(0) = '1' then
                    state_var5923 := Q_WAIT4777;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(\$18613_copy_root_in_ram6634346_arg\(0 to 15)));
                    state_var5923 := PAUSE_GET4776;
                  end if;
                end if;
              when \$18625_COPY_ROOT_IN_RAM6634345\ =>
                \$v4755\ := work.Int.ge(\$18625_copy_root_in_ram6634345_arg\(0 to 15), \$18625_copy_root_in_ram6634345_arg\(16 to 31));
                if \$v4755\(0) = '1' then
                  \$18625_copy_root_in_ram6634345_result\ := \$18625_copy_root_in_ram6634345_arg\(32 to 47);
                  \$18613_copy_root_in_ram6634346_result\ := \$18625_copy_root_in_ram6634345_result\;
                  \$18534_next\ := \$18613_copy_root_in_ram6634346_result\;
                  \$v4731\ := \$global_end_lock\;
                  if \$v4731\(0) = '1' then
                    state_var5923 := Q_WAIT4730;
                  else
                    acquire(\$global_end_lock\);
                    \$global_end_ptr\ <= 0;
                    state_var5923 := PAUSE_GET4729;
                  end if;
                else
                  \$18628\ := work.Print.print_string(clk,of_string("racine:"));
                  \$18629\ := work.Int.print(clk,\$18625_copy_root_in_ram6634345_arg\(0 to 15));
                  \$18630\ := work.Print.print_newline(clk,eclat_unit);
                  \$v4754\ := \$ram_lock\;
                  if \$v4754\(0) = '1' then
                    state_var5923 := Q_WAIT4753;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(\$18625_copy_root_in_ram6634345_arg\(0 to 15)));
                    state_var5923 := PAUSE_GET4752;
                  end if;
                end if;
              when PAUSE_GET4613 =>
                \$18761\ := \$ram_value\;
                release(\$ram_lock\);
                \$v4612\ := \$ram_lock\;
                if \$v4612\(0) = '1' then
                  state_var5923 := Q_WAIT4611;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$18521_loop666_arg\(16 to 31), \$18521_loop666_arg\(0 to 15))));
                  \$ram_write\ <= \$18761\; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4610;
                end if;
              when PAUSE_GET4629 =>
                \$18745_hd\ := \$ram_value\;
                release(\$ram_lock\);
                \$18746\ := work.Print.print_string(clk,of_string("bloc "));
                \$18747\ := work.Int.print(clk,eclat_resize(\$18741\(0 to 30),16));
                \$18748\ := work.Print.print_string(clk,of_string(" of size "));
                \$18749\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                            work.Int.lsr(
                                                            \$18745_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$18750\ := work.Print.print_string(clk,of_string(" from "));
                \$18751\ := work.Int.print(clk,eclat_resize(\$18741\(0 to 30),16));
                \$18752\ := work.Print.print_string(clk,of_string(" to "));
                \$18753\ := work.Int.print(clk,\$18522_loop665_arg\(16 to 31));
                \$18754\ := work.Print.print_newline(clk,eclat_unit);
                \$v4628\ := \$ram_lock\;
                if \$v4628\(0) = '1' then
                  state_var5923 := Q_WAIT4627;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18522_loop665_arg\(16 to 31)));
                  \$ram_write\ <= \$18745_hd\; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4626;
                end if;
              when PAUSE_GET4633 =>
                \$18744_w\ := \$ram_value\;
                release(\$ram_lock\);
                \$v4632\ := eclat_if(work.Bool.lnot(""&\$18744_w\(31)) & 
                            eclat_if(work.Int.le(\$18522_loop665_arg\(48 to 63), eclat_resize(\$18744_w\(0 to 30),16)) & 
                            work.Int.lt(eclat_resize(\$18744_w\(0 to 30),16), 
                                        work.Int.add(\$18522_loop665_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false);
                if \$v4632\(0) = '1' then
                  \$18742\ := \$18744_w\ & \$18522_loop665_arg\(16 to 31);
                  \$v4619\ := \$ram_lock\;
                  if \$v4619\(0) = '1' then
                    state_var5923 := Q_WAIT4618;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            \$18522_loop665_arg\(64 to 79), \$18522_loop665_arg\(0 to 15))));
                    \$ram_write\ <= \$18742\(0 to 31); \$ram_write_request\ <= '1';
                    state_var5923 := PAUSE_SET4617;
                  end if;
                else
                  \$v4631\ := \$ram_lock\;
                  if \$v4631\(0) = '1' then
                    state_var5923 := Q_WAIT4630;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18741\(0 to 30),16)));
                    state_var5923 := PAUSE_GET4629;
                  end if;
                end if;
              when PAUSE_GET4637 =>
                \$18741\ := \$ram_value\;
                release(\$ram_lock\);
                \$v4636\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$18741\(31)) & 
                                           eclat_if(work.Int.le(\$18522_loop665_arg\(32 to 47), eclat_resize(\$18741\(0 to 30),16)) & 
                                           work.Int.lt(eclat_resize(\$18741\(0 to 30),16), 
                                                       work.Int.add(\$18522_loop665_arg\(32 to 47), X"1770")) & eclat_false) & eclat_false));
                if \$v4636\(0) = '1' then
                  \$18742\ := \$18741\ & \$18522_loop665_arg\(16 to 31);
                  \$v4619\ := \$ram_lock\;
                  if \$v4619\(0) = '1' then
                    state_var5923 := Q_WAIT4618;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            \$18522_loop665_arg\(64 to 79), \$18522_loop665_arg\(0 to 15))));
                    \$ram_write\ <= \$18742\(0 to 31); \$ram_write_request\ <= '1';
                    state_var5923 := PAUSE_SET4617;
                  end if;
                else
                  \$v4635\ := \$ram_lock\;
                  if \$v4635\(0) = '1' then
                    state_var5923 := Q_WAIT4634;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18741\(0 to 30),16), X"000" & X"1")));
                    state_var5923 := PAUSE_GET4633;
                  end if;
                end if;
              when PAUSE_GET4641 =>
                \$18737\ := \$ram_value\;
                release(\$ram_lock\);
                \$18522_loop665_id\ := "000000001111";
                \$18522_loop665_arg\ := X"000" & X"1" & \$18523_aux664_arg\(16 to 31) & \$18523_aux664_arg\(32 to 47) & \$18523_aux664_arg\(48 to 63) & \$18523_aux664_arg\(0 to 15) & eclat_resize(
                work.Int.lsr(eclat_resize(eclat_resize(\$18737\(0 to 30),16),31), X"0000000" & X"2"),16);
                state_var5923 := \$18522_LOOP665\;
              when PAUSE_GET4648 =>
                \$18728\ := \$ram_value\;
                release(\$ram_lock\);
                \$v4647\ := \$ram_lock\;
                if \$v4647\(0) = '1' then
                  state_var5923 := Q_WAIT4646;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$18524_loop666_arg\(16 to 31), \$18524_loop666_arg\(0 to 15))));
                  \$ram_write\ <= \$18728\; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4645;
                end if;
              when PAUSE_GET4664 =>
                \$18712_hd\ := \$ram_value\;
                release(\$ram_lock\);
                \$18713\ := work.Print.print_string(clk,of_string("bloc "));
                \$18714\ := work.Int.print(clk,eclat_resize(\$18708\(0 to 30),16));
                \$18715\ := work.Print.print_string(clk,of_string(" of size "));
                \$18716\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                            work.Int.lsr(
                                                            \$18712_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$18717\ := work.Print.print_string(clk,of_string(" from "));
                \$18718\ := work.Int.print(clk,eclat_resize(\$18708\(0 to 30),16));
                \$18719\ := work.Print.print_string(clk,of_string(" to "));
                \$18720\ := work.Int.print(clk,\$18525_loop665_arg\(16 to 31));
                \$18721\ := work.Print.print_newline(clk,eclat_unit);
                \$v4663\ := \$ram_lock\;
                if \$v4663\(0) = '1' then
                  state_var5923 := Q_WAIT4662;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18525_loop665_arg\(16 to 31)));
                  \$ram_write\ <= \$18712_hd\; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4661;
                end if;
              when PAUSE_GET4668 =>
                \$18711_w\ := \$ram_value\;
                release(\$ram_lock\);
                \$v4667\ := eclat_if(work.Bool.lnot(""&\$18711_w\(31)) & 
                            eclat_if(work.Int.le(\$18525_loop665_arg\(48 to 63), eclat_resize(\$18711_w\(0 to 30),16)) & 
                            work.Int.lt(eclat_resize(\$18711_w\(0 to 30),16), 
                                        work.Int.add(\$18525_loop665_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false);
                if \$v4667\(0) = '1' then
                  \$18709\ := \$18711_w\ & \$18525_loop665_arg\(16 to 31);
                  \$v4654\ := \$ram_lock\;
                  if \$v4654\(0) = '1' then
                    state_var5923 := Q_WAIT4653;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            \$18525_loop665_arg\(64 to 79), \$18525_loop665_arg\(0 to 15))));
                    \$ram_write\ <= \$18709\(0 to 31); \$ram_write_request\ <= '1';
                    state_var5923 := PAUSE_SET4652;
                  end if;
                else
                  \$v4666\ := \$ram_lock\;
                  if \$v4666\(0) = '1' then
                    state_var5923 := Q_WAIT4665;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18708\(0 to 30),16)));
                    state_var5923 := PAUSE_GET4664;
                  end if;
                end if;
              when PAUSE_GET4672 =>
                \$18708\ := \$ram_value\;
                release(\$ram_lock\);
                \$v4671\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$18708\(31)) & 
                                           eclat_if(work.Int.le(\$18525_loop665_arg\(32 to 47), eclat_resize(\$18708\(0 to 30),16)) & 
                                           work.Int.lt(eclat_resize(\$18708\(0 to 30),16), 
                                                       work.Int.add(\$18525_loop665_arg\(32 to 47), X"1770")) & eclat_false) & eclat_false));
                if \$v4671\(0) = '1' then
                  \$18709\ := \$18708\ & \$18525_loop665_arg\(16 to 31);
                  \$v4654\ := \$ram_lock\;
                  if \$v4654\(0) = '1' then
                    state_var5923 := Q_WAIT4653;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            \$18525_loop665_arg\(64 to 79), \$18525_loop665_arg\(0 to 15))));
                    \$ram_write\ <= \$18709\(0 to 31); \$ram_write_request\ <= '1';
                    state_var5923 := PAUSE_SET4652;
                  end if;
                else
                  \$v4670\ := \$ram_lock\;
                  if \$v4670\(0) = '1' then
                    state_var5923 := Q_WAIT4669;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18708\(0 to 30),16), X"000" & X"1")));
                    state_var5923 := PAUSE_GET4668;
                  end if;
                end if;
              when PAUSE_GET4676 =>
                \$18704\ := \$ram_value\;
                release(\$ram_lock\);
                \$18525_loop665_id\ := "000000010001";
                \$18525_loop665_arg\ := X"000" & X"1" & \$18526_aux664_arg\(16 to 31) & \$18526_aux664_arg\(32 to 47) & \$18526_aux664_arg\(48 to 63) & \$18526_aux664_arg\(0 to 15) & eclat_resize(
                work.Int.lsr(eclat_resize(eclat_resize(\$18704\(0 to 30),16),31), X"0000000" & X"2"),16);
                state_var5923 := \$18525_LOOP665\;
              when PAUSE_GET4693 =>
                \$18584_hd\ := \$ram_value\;
                release(\$ram_lock\);
                \$18585\ := work.Print.print_string(clk,of_string("bloc "));
                \$18586\ := work.Int.print(clk,eclat_resize(\$18577\(0 to 30),16));
                \$18587\ := work.Print.print_string(clk,of_string(" of size "));
                \$18588\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                            work.Int.lsr(
                                                            \$18584_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$18589\ := work.Print.print_string(clk,of_string(" from "));
                \$18590\ := work.Int.print(clk,eclat_resize(\$18577\(0 to 30),16));
                \$18591\ := work.Print.print_string(clk,of_string(" to "));
                \$18592\ := work.Int.print(clk,\$18571_copy_root_in_ram6634345_arg\(32 to 47));
                \$18593\ := work.Print.print_newline(clk,eclat_unit);
                \$v4692\ := \$ram_lock\;
                if \$v4692\(0) = '1' then
                  state_var5923 := Q_WAIT4691;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18571_copy_root_in_ram6634345_arg\(32 to 47)));
                  \$ram_write\ <= \$18584_hd\; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4690;
                end if;
              when PAUSE_GET4697 =>
                \$18583_w\ := \$ram_value\;
                release(\$ram_lock\);
                \$v4696\ := eclat_if(work.Bool.lnot(""&\$18583_w\(31)) & 
                            eclat_if(work.Int.le(\$18571_copy_root_in_ram6634345_arg\(64 to 79), eclat_resize(\$18583_w\(0 to 30),16)) & 
                            work.Int.lt(eclat_resize(\$18583_w\(0 to 30),16), 
                                        work.Int.add(\$18571_copy_root_in_ram6634345_arg\(64 to 79), X"1770")) & eclat_false) & eclat_false);
                if \$v4696\(0) = '1' then
                  \$18578\ := \$18583_w\ & \$18571_copy_root_in_ram6634345_arg\(32 to 47);
                  \$v4683\ := \$ram_lock\;
                  if \$v4683\(0) = '1' then
                    state_var5923 := Q_WAIT4682;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18571_copy_root_in_ram6634345_arg\(0 to 15)));
                    \$ram_write\ <= \$18578\(0 to 31); \$ram_write_request\ <= '1';
                    state_var5923 := PAUSE_SET4681;
                  end if;
                else
                  \$v4695\ := \$ram_lock\;
                  if \$v4695\(0) = '1' then
                    state_var5923 := Q_WAIT4694;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18577\(0 to 30),16)));
                    state_var5923 := PAUSE_GET4693;
                  end if;
                end if;
              when PAUSE_GET4701 =>
                \$18577\ := \$ram_value\;
                release(\$ram_lock\);
                \$v4700\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$18577\(31)) & 
                                           eclat_if(work.Int.le(\$18571_copy_root_in_ram6634345_arg\(48 to 63), eclat_resize(\$18577\(0 to 30),16)) & 
                                           work.Int.lt(eclat_resize(\$18577\(0 to 30),16), 
                                                       work.Int.add(\$18571_copy_root_in_ram6634345_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false));
                if \$v4700\(0) = '1' then
                  \$18578\ := \$18577\ & \$18571_copy_root_in_ram6634345_arg\(32 to 47);
                  \$v4683\ := \$ram_lock\;
                  if \$v4683\(0) = '1' then
                    state_var5923 := Q_WAIT4682;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18571_copy_root_in_ram6634345_arg\(0 to 15)));
                    \$ram_write\ <= \$18578\(0 to 31); \$ram_write_request\ <= '1';
                    state_var5923 := PAUSE_SET4681;
                  end if;
                else
                  \$v4699\ := \$ram_lock\;
                  if \$v4699\(0) = '1' then
                    state_var5923 := Q_WAIT4698;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18577\(0 to 30),16), X"000" & X"1")));
                    state_var5923 := PAUSE_GET4697;
                  end if;
                end if;
              when PAUSE_GET4717 =>
                \$18599_hd\ := \$ram_value\;
                release(\$ram_lock\);
                \$18600\ := work.Print.print_string(clk,of_string("bloc "));
                \$18601\ := work.Int.print(clk,eclat_resize(\$18565\(0 to 30),16));
                \$18602\ := work.Print.print_string(clk,of_string(" of size "));
                \$18603\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                            work.Int.lsr(
                                                            \$18599_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$18604\ := work.Print.print_string(clk,of_string(" from "));
                \$18605\ := work.Int.print(clk,eclat_resize(\$18565\(0 to 30),16));
                \$18606\ := work.Print.print_string(clk,of_string(" to "));
                \$18607\ := work.Int.print(clk,\$18559_copy_root_in_ram6634347_arg\(32 to 47));
                \$18608\ := work.Print.print_newline(clk,eclat_unit);
                \$v4716\ := \$ram_lock\;
                if \$v4716\(0) = '1' then
                  state_var5923 := Q_WAIT4715;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18559_copy_root_in_ram6634347_arg\(32 to 47)));
                  \$ram_write\ <= \$18599_hd\; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4714;
                end if;
              when PAUSE_GET4721 =>
                \$18598_w\ := \$ram_value\;
                release(\$ram_lock\);
                \$v4720\ := eclat_if(work.Bool.lnot(""&\$18598_w\(31)) & 
                            eclat_if(work.Int.le(\$18559_copy_root_in_ram6634347_arg\(64 to 79), eclat_resize(\$18598_w\(0 to 30),16)) & 
                            work.Int.lt(eclat_resize(\$18598_w\(0 to 30),16), 
                                        work.Int.add(\$18559_copy_root_in_ram6634347_arg\(64 to 79), X"1770")) & eclat_false) & eclat_false);
                if \$v4720\(0) = '1' then
                  \$18566\ := \$18598_w\ & \$18559_copy_root_in_ram6634347_arg\(32 to 47);
                  \$v4707\ := \$ram_lock\;
                  if \$v4707\(0) = '1' then
                    state_var5923 := Q_WAIT4706;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18559_copy_root_in_ram6634347_arg\(0 to 15)));
                    \$ram_write\ <= \$18566\(0 to 31); \$ram_write_request\ <= '1';
                    state_var5923 := PAUSE_SET4705;
                  end if;
                else
                  \$v4719\ := \$ram_lock\;
                  if \$v4719\(0) = '1' then
                    state_var5923 := Q_WAIT4718;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18565\(0 to 30),16)));
                    state_var5923 := PAUSE_GET4717;
                  end if;
                end if;
              when PAUSE_GET4725 =>
                \$18565\ := \$ram_value\;
                release(\$ram_lock\);
                \$v4724\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$18565\(31)) & 
                                           eclat_if(work.Int.le(\$18559_copy_root_in_ram6634347_arg\(48 to 63), eclat_resize(\$18565\(0 to 30),16)) & 
                                           work.Int.lt(eclat_resize(\$18565\(0 to 30),16), 
                                                       work.Int.add(\$18559_copy_root_in_ram6634347_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false));
                if \$v4724\(0) = '1' then
                  \$18566\ := \$18565\ & \$18559_copy_root_in_ram6634347_arg\(32 to 47);
                  \$v4707\ := \$ram_lock\;
                  if \$v4707\(0) = '1' then
                    state_var5923 := Q_WAIT4706;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18559_copy_root_in_ram6634347_arg\(0 to 15)));
                    \$ram_write\ <= \$18566\(0 to 31); \$ram_write_request\ <= '1';
                    state_var5923 := PAUSE_SET4705;
                  end if;
                else
                  \$v4723\ := \$ram_lock\;
                  if \$v4723\(0) = '1' then
                    state_var5923 := Q_WAIT4722;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18565\(0 to 30),16), X"000" & X"1")));
                    state_var5923 := PAUSE_GET4721;
                  end if;
                end if;
              when PAUSE_GET4729 =>
                \$18541\ := \$global_end_value\;
                release(\$global_end_lock\);
                \$18559_copy_root_in_ram6634347_id\ := "000000011000";
                \$18559_copy_root_in_ram6634347_arg\ := X"3e80" & \$18541\ & \$18534_next\ & \$18520\(96 to 111) & \$18520\(112 to 127);
                state_var5923 := \$18559_COPY_ROOT_IN_RAM6634347\;
              when PAUSE_GET4744 =>
                \$18638_hd\ := \$ram_value\;
                release(\$ram_lock\);
                \$18639\ := work.Print.print_string(clk,of_string("bloc "));
                \$18640\ := work.Int.print(clk,eclat_resize(\$18631\(0 to 30),16));
                \$18641\ := work.Print.print_string(clk,of_string(" of size "));
                \$18642\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                            work.Int.lsr(
                                                            \$18638_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$18643\ := work.Print.print_string(clk,of_string(" from "));
                \$18644\ := work.Int.print(clk,eclat_resize(\$18631\(0 to 30),16));
                \$18645\ := work.Print.print_string(clk,of_string(" to "));
                \$18646\ := work.Int.print(clk,\$18625_copy_root_in_ram6634345_arg\(32 to 47));
                \$18647\ := work.Print.print_newline(clk,eclat_unit);
                \$v4743\ := \$ram_lock\;
                if \$v4743\(0) = '1' then
                  state_var5923 := Q_WAIT4742;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18625_copy_root_in_ram6634345_arg\(32 to 47)));
                  \$ram_write\ <= \$18638_hd\; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4741;
                end if;
              when PAUSE_GET4748 =>
                \$18637_w\ := \$ram_value\;
                release(\$ram_lock\);
                \$v4747\ := eclat_if(work.Bool.lnot(""&\$18637_w\(31)) & 
                            eclat_if(work.Int.le(\$18625_copy_root_in_ram6634345_arg\(64 to 79), eclat_resize(\$18637_w\(0 to 30),16)) & 
                            work.Int.lt(eclat_resize(\$18637_w\(0 to 30),16), 
                                        work.Int.add(\$18625_copy_root_in_ram6634345_arg\(64 to 79), X"1770")) & eclat_false) & eclat_false);
                if \$v4747\(0) = '1' then
                  \$18632\ := \$18637_w\ & \$18625_copy_root_in_ram6634345_arg\(32 to 47);
                  \$v4734\ := \$ram_lock\;
                  if \$v4734\(0) = '1' then
                    state_var5923 := Q_WAIT4733;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18625_copy_root_in_ram6634345_arg\(0 to 15)));
                    \$ram_write\ <= \$18632\(0 to 31); \$ram_write_request\ <= '1';
                    state_var5923 := PAUSE_SET4732;
                  end if;
                else
                  \$v4746\ := \$ram_lock\;
                  if \$v4746\(0) = '1' then
                    state_var5923 := Q_WAIT4745;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18631\(0 to 30),16)));
                    state_var5923 := PAUSE_GET4744;
                  end if;
                end if;
              when PAUSE_GET4752 =>
                \$18631\ := \$ram_value\;
                release(\$ram_lock\);
                \$v4751\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$18631\(31)) & 
                                           eclat_if(work.Int.le(\$18625_copy_root_in_ram6634345_arg\(48 to 63), eclat_resize(\$18631\(0 to 30),16)) & 
                                           work.Int.lt(eclat_resize(\$18631\(0 to 30),16), 
                                                       work.Int.add(\$18625_copy_root_in_ram6634345_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false));
                if \$v4751\(0) = '1' then
                  \$18632\ := \$18631\ & \$18625_copy_root_in_ram6634345_arg\(32 to 47);
                  \$v4734\ := \$ram_lock\;
                  if \$v4734\(0) = '1' then
                    state_var5923 := Q_WAIT4733;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18625_copy_root_in_ram6634345_arg\(0 to 15)));
                    \$ram_write\ <= \$18632\(0 to 31); \$ram_write_request\ <= '1';
                    state_var5923 := PAUSE_SET4732;
                  end if;
                else
                  \$v4750\ := \$ram_lock\;
                  if \$v4750\(0) = '1' then
                    state_var5923 := Q_WAIT4749;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18631\(0 to 30),16), X"000" & X"1")));
                    state_var5923 := PAUSE_GET4748;
                  end if;
                end if;
              when PAUSE_GET4768 =>
                \$18653_hd\ := \$ram_value\;
                release(\$ram_lock\);
                \$18654\ := work.Print.print_string(clk,of_string("bloc "));
                \$18655\ := work.Int.print(clk,eclat_resize(\$18619\(0 to 30),16));
                \$18656\ := work.Print.print_string(clk,of_string(" of size "));
                \$18657\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                            work.Int.lsr(
                                                            \$18653_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$18658\ := work.Print.print_string(clk,of_string(" from "));
                \$18659\ := work.Int.print(clk,eclat_resize(\$18619\(0 to 30),16));
                \$18660\ := work.Print.print_string(clk,of_string(" to "));
                \$18661\ := work.Int.print(clk,\$18613_copy_root_in_ram6634346_arg\(32 to 47));
                \$18662\ := work.Print.print_newline(clk,eclat_unit);
                \$v4767\ := \$ram_lock\;
                if \$v4767\(0) = '1' then
                  state_var5923 := Q_WAIT4766;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18613_copy_root_in_ram6634346_arg\(32 to 47)));
                  \$ram_write\ <= \$18653_hd\; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4765;
                end if;
              when PAUSE_GET4772 =>
                \$18652_w\ := \$ram_value\;
                release(\$ram_lock\);
                \$v4771\ := eclat_if(work.Bool.lnot(""&\$18652_w\(31)) & 
                            eclat_if(work.Int.le(\$18613_copy_root_in_ram6634346_arg\(64 to 79), eclat_resize(\$18652_w\(0 to 30),16)) & 
                            work.Int.lt(eclat_resize(\$18652_w\(0 to 30),16), 
                                        work.Int.add(\$18613_copy_root_in_ram6634346_arg\(64 to 79), X"1770")) & eclat_false) & eclat_false);
                if \$v4771\(0) = '1' then
                  \$18620\ := \$18652_w\ & \$18613_copy_root_in_ram6634346_arg\(32 to 47);
                  \$v4758\ := \$ram_lock\;
                  if \$v4758\(0) = '1' then
                    state_var5923 := Q_WAIT4757;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18613_copy_root_in_ram6634346_arg\(0 to 15)));
                    \$ram_write\ <= \$18620\(0 to 31); \$ram_write_request\ <= '1';
                    state_var5923 := PAUSE_SET4756;
                  end if;
                else
                  \$v4770\ := \$ram_lock\;
                  if \$v4770\(0) = '1' then
                    state_var5923 := Q_WAIT4769;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18619\(0 to 30),16)));
                    state_var5923 := PAUSE_GET4768;
                  end if;
                end if;
              when PAUSE_GET4776 =>
                \$18619\ := \$ram_value\;
                release(\$ram_lock\);
                \$v4775\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$18619\(31)) & 
                                           eclat_if(work.Int.le(\$18613_copy_root_in_ram6634346_arg\(48 to 63), eclat_resize(\$18619\(0 to 30),16)) & 
                                           work.Int.lt(eclat_resize(\$18619\(0 to 30),16), 
                                                       work.Int.add(\$18613_copy_root_in_ram6634346_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false));
                if \$v4775\(0) = '1' then
                  \$18620\ := \$18619\ & \$18613_copy_root_in_ram6634346_arg\(32 to 47);
                  \$v4758\ := \$ram_lock\;
                  if \$v4758\(0) = '1' then
                    state_var5923 := Q_WAIT4757;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18613_copy_root_in_ram6634346_arg\(0 to 15)));
                    \$ram_write\ <= \$18620\(0 to 31); \$ram_write_request\ <= '1';
                    state_var5923 := PAUSE_SET4756;
                  end if;
                else
                  \$v4774\ := \$ram_lock\;
                  if \$v4774\(0) = '1' then
                    state_var5923 := Q_WAIT4773;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18619\(0 to 30),16), X"000" & X"1")));
                    state_var5923 := PAUSE_GET4772;
                  end if;
                end if;
              when PAUSE_GET4789 =>
                \$18668_hd\ := \$ram_value\;
                release(\$ram_lock\);
                \$18669\ := work.Print.print_string(clk,of_string("bloc "));
                \$18670\ := work.Int.print(clk,eclat_resize(\$18468_wait662_arg\(33 to 63),16));
                \$18671\ := work.Print.print_string(clk,of_string(" of size "));
                \$18672\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                            work.Int.lsr(
                                                            \$18668_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$18673\ := work.Print.print_string(clk,of_string(" from "));
                \$18674\ := work.Int.print(clk,eclat_resize(\$18468_wait662_arg\(33 to 63),16));
                \$18675\ := work.Print.print_string(clk,of_string(" to "));
                \$18676\ := work.Int.print(clk,\$18532\(32 to 47));
                \$18677\ := work.Print.print_newline(clk,eclat_unit);
                \$v4788\ := \$ram_lock\;
                if \$v4788\(0) = '1' then
                  state_var5923 := Q_WAIT4787;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18532\(32 to 47)));
                  \$ram_write\ <= \$18668_hd\; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4786;
                end if;
              when PAUSE_GET4793 =>
                \$18667_w\ := \$ram_value\;
                release(\$ram_lock\);
                \$v4792\ := eclat_if(work.Bool.lnot(""&\$18667_w\(31)) & 
                            eclat_if(work.Int.le(\$18520\(112 to 127), eclat_resize(\$18667_w\(0 to 30),16)) & 
                            work.Int.lt(eclat_resize(\$18667_w\(0 to 30),16), 
                                        work.Int.add(\$18520\(112 to 127), X"1770")) & eclat_false) & eclat_false);
                if \$v4792\(0) = '1' then
                  \$18533\ := \$18667_w\ & \$18532\(32 to 47);
                  \$18613_copy_root_in_ram6634346_id\ := "000000011100";
                  \$18613_copy_root_in_ram6634346_arg\ := X"0" & X"3e8" & \$18468_wait662_arg\(65 to 80) & \$18533\(32 to 47) & \$18520\(96 to 111) & \$18520\(112 to 127);
                  state_var5923 := \$18613_COPY_ROOT_IN_RAM6634346\;
                else
                  \$v4791\ := \$ram_lock\;
                  if \$v4791\(0) = '1' then
                    state_var5923 := Q_WAIT4790;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18468_wait662_arg\(33 to 63),16)));
                    state_var5923 := PAUSE_GET4789;
                  end if;
                end if;
              when PAUSE_GET4806 =>
                \$18683_hd\ := \$ram_value\;
                release(\$ram_lock\);
                \$18684\ := work.Print.print_string(clk,of_string("bloc "));
                \$18685\ := work.Int.print(clk,eclat_resize(\$18468_wait662_arg\(1 to 31),16));
                \$18686\ := work.Print.print_string(clk,of_string(" of size "));
                \$18687\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                            work.Int.lsr(
                                                            \$18683_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$18688\ := work.Print.print_string(clk,of_string(" from "));
                \$18689\ := work.Int.print(clk,eclat_resize(\$18468_wait662_arg\(1 to 31),16));
                \$18690\ := work.Print.print_string(clk,of_string(" to "));
                \$18691\ := work.Int.print(clk,\$18520\(112 to 127));
                \$18692\ := work.Print.print_newline(clk,eclat_unit);
                \$v4805\ := \$ram_lock\;
                if \$v4805\(0) = '1' then
                  state_var5923 := Q_WAIT4804;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18520\(112 to 127)));
                  \$ram_write\ <= \$18683_hd\; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4803;
                end if;
              when PAUSE_GET4810 =>
                \$18682_w\ := \$ram_value\;
                release(\$ram_lock\);
                \$v4809\ := eclat_if(work.Bool.lnot(""&\$18682_w\(31)) & 
                            eclat_if(work.Int.le(\$18520\(112 to 127), eclat_resize(\$18682_w\(0 to 30),16)) & 
                            work.Int.lt(eclat_resize(\$18682_w\(0 to 30),16), 
                                        work.Int.add(\$18520\(112 to 127), X"1770")) & eclat_false) & eclat_false);
                if \$v4809\(0) = '1' then
                  \$18532\ := \$18682_w\ & \$18520\(112 to 127);
                  \$v4796\ := work.Bool.lnot(eclat_if(work.Bool.lnot(
                                                      ""&\$18468_wait662_arg\(64)) & 
                                             eclat_if(work.Int.le(\$18520\(96 to 111), eclat_resize(\$18468_wait662_arg\(33 to 63),16)) & 
                                             work.Int.lt(eclat_resize(\$18468_wait662_arg\(33 to 63),16), 
                                                         work.Int.add(
                                                         \$18520\(96 to 111), X"1770")) & eclat_false) & eclat_false));
                  if \$v4796\(0) = '1' then
                    \$18533\ := \$18468_wait662_arg\(33 to 64) & \$18532\(32 to 47);
                    \$18613_copy_root_in_ram6634346_id\ := "000000011100";
                    \$18613_copy_root_in_ram6634346_arg\ := X"0" & X"3e8" & \$18468_wait662_arg\(65 to 80) & \$18533\(32 to 47) & \$18520\(96 to 111) & \$18520\(112 to 127);
                    state_var5923 := \$18613_COPY_ROOT_IN_RAM6634346\;
                  else
                    \$v4795\ := \$ram_lock\;
                    if \$v4795\(0) = '1' then
                      state_var5923 := Q_WAIT4794;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                        eclat_resize(\$18468_wait662_arg\(33 to 63),16), X"000" & X"1")));
                      state_var5923 := PAUSE_GET4793;
                    end if;
                  end if;
                else
                  \$v4808\ := \$ram_lock\;
                  if \$v4808\(0) = '1' then
                    state_var5923 := Q_WAIT4807;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18468_wait662_arg\(1 to 31),16)));
                    state_var5923 := PAUSE_GET4806;
                  end if;
                end if;
              when PAUSE_SET4610 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18762\ := eclat_unit;
                \$18521_loop666_arg\ := work.Int.add(\$18521_loop666_arg\(0 to 15), X"000" & X"1") & \$18521_loop666_arg\(16 to 31) & \$18521_loop666_arg\(32 to 47) & \$18521_loop666_arg\(48 to 63);
                state_var5923 := \$18521_LOOP666\;
              when PAUSE_SET4617 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18743\ := eclat_unit;
                \$18522_loop665_arg\ := work.Int.add(\$18522_loop665_arg\(0 to 15), X"000" & X"1") & \$18742\(32 to 47) & \$18522_loop665_arg\(32 to 47) & \$18522_loop665_arg\(48 to 63) & \$18522_loop665_arg\(64 to 79) & \$18522_loop665_arg\(80 to 95);
                state_var5923 := \$18522_LOOP665\;
              when PAUSE_SET4620 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18758\ := eclat_unit;
                \$18742\ := eclat_resize(\$18522_loop665_arg\(16 to 31),31) & eclat_false & 
                work.Int.add(\$18522_loop665_arg\(16 to 31), work.Int.add(
                                                             eclat_resize(
                                                             work.Int.lsr(
                                                             \$18745_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$v4619\ := \$ram_lock\;
                if \$v4619\(0) = '1' then
                  state_var5923 := Q_WAIT4618;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$18522_loop665_arg\(64 to 79), \$18522_loop665_arg\(0 to 15))));
                  \$ram_write\ <= \$18742\(0 to 31); \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4617;
                end if;
              when PAUSE_SET4623 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18757\ := eclat_unit;
                \$v4622\ := \$ram_lock\;
                if \$v4622\(0) = '1' then
                  state_var5923 := Q_WAIT4621;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$18741\(0 to 30),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$18522_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4620;
                end if;
              when PAUSE_SET4626 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18755\ := eclat_unit;
                \$18521_loop666_id\ := "000000001110";
                \$18521_loop666_arg\ := X"000" & X"1" & \$18522_loop665_arg\(16 to 31) & eclat_resize(\$18741\(0 to 30),16) & eclat_resize(
                work.Int.lsr(\$18745_hd\(0 to 30), X"0000000" & X"2"),16);
                state_var5923 := \$18521_LOOP666\;
              when PAUSE_SET4645 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18729\ := eclat_unit;
                \$18524_loop666_arg\ := work.Int.add(\$18524_loop666_arg\(0 to 15), X"000" & X"1") & \$18524_loop666_arg\(16 to 31) & \$18524_loop666_arg\(32 to 47) & \$18524_loop666_arg\(48 to 63);
                state_var5923 := \$18524_LOOP666\;
              when PAUSE_SET4652 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18710\ := eclat_unit;
                \$18525_loop665_arg\ := work.Int.add(\$18525_loop665_arg\(0 to 15), X"000" & X"1") & \$18709\(32 to 47) & \$18525_loop665_arg\(32 to 47) & \$18525_loop665_arg\(48 to 63) & \$18525_loop665_arg\(64 to 79) & \$18525_loop665_arg\(80 to 95);
                state_var5923 := \$18525_LOOP665\;
              when PAUSE_SET4655 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18725\ := eclat_unit;
                \$18709\ := eclat_resize(\$18525_loop665_arg\(16 to 31),31) & eclat_false & 
                work.Int.add(\$18525_loop665_arg\(16 to 31), work.Int.add(
                                                             eclat_resize(
                                                             work.Int.lsr(
                                                             \$18712_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$v4654\ := \$ram_lock\;
                if \$v4654\(0) = '1' then
                  state_var5923 := Q_WAIT4653;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$18525_loop665_arg\(64 to 79), \$18525_loop665_arg\(0 to 15))));
                  \$ram_write\ <= \$18709\(0 to 31); \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4652;
                end if;
              when PAUSE_SET4658 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18724\ := eclat_unit;
                \$v4657\ := \$ram_lock\;
                if \$v4657\(0) = '1' then
                  state_var5923 := Q_WAIT4656;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$18708\(0 to 30),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$18525_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4655;
                end if;
              when PAUSE_SET4661 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18722\ := eclat_unit;
                \$18524_loop666_id\ := "000000010000";
                \$18524_loop666_arg\ := X"000" & X"1" & \$18525_loop665_arg\(16 to 31) & eclat_resize(\$18708\(0 to 30),16) & eclat_resize(
                work.Int.lsr(\$18712_hd\(0 to 30), X"0000000" & X"2"),16);
                state_var5923 := \$18524_LOOP666\;
              when PAUSE_SET4681 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18579\ := eclat_unit;
                \$18580\ := work.Print.print_string(clk,of_string(" next="));
                \$18581\ := work.Int.print(clk,\$18578\(32 to 47));
                \$18582\ := work.Print.print_newline(clk,eclat_unit);
                \$18571_copy_root_in_ram6634345_arg\ := work.Int.add(
                                                        \$18571_copy_root_in_ram6634345_arg\(0 to 15), X"000" & X"1") & \$18571_copy_root_in_ram6634345_arg\(16 to 31) & \$18578\(32 to 47) & \$18571_copy_root_in_ram6634345_arg\(48 to 63) & \$18571_copy_root_in_ram6634345_arg\(64 to 79);
                state_var5923 := \$18571_COPY_ROOT_IN_RAM6634345\;
              when PAUSE_SET4684 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18597\ := eclat_unit;
                \$18578\ := eclat_resize(\$18571_copy_root_in_ram6634345_arg\(32 to 47),31) & eclat_false & 
                work.Int.add(\$18571_copy_root_in_ram6634345_arg\(32 to 47), 
                             work.Int.add(eclat_resize(work.Int.lsr(\$18584_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$v4683\ := \$ram_lock\;
                if \$v4683\(0) = '1' then
                  state_var5923 := Q_WAIT4682;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18571_copy_root_in_ram6634345_arg\(0 to 15)));
                  \$ram_write\ <= \$18578\(0 to 31); \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4681;
                end if;
              when PAUSE_SET4687 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18596\ := eclat_unit;
                \$v4686\ := \$ram_lock\;
                if \$v4686\(0) = '1' then
                  state_var5923 := Q_WAIT4685;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$18577\(0 to 30),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$18571_copy_root_in_ram6634345_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4684;
                end if;
              when PAUSE_SET4690 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18594\ := eclat_unit;
                \$18524_loop666_id\ := "000000010101";
                \$18524_loop666_arg\ := X"000" & X"1" & \$18571_copy_root_in_ram6634345_arg\(32 to 47) & eclat_resize(\$18577\(0 to 30),16) & eclat_resize(
                work.Int.lsr(\$18584_hd\(0 to 30), X"0000000" & X"2"),16);
                state_var5923 := \$18524_LOOP666\;
              when PAUSE_SET4705 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18567\ := eclat_unit;
                \$18568\ := work.Print.print_string(clk,of_string(" next="));
                \$18569\ := work.Int.print(clk,\$18566\(32 to 47));
                \$18570\ := work.Print.print_newline(clk,eclat_unit);
                \$18571_copy_root_in_ram6634345_id\ := "000000010110";
                \$18571_copy_root_in_ram6634345_arg\ := work.Int.add(
                                                        \$18559_copy_root_in_ram6634347_arg\(0 to 15), X"000" & X"1") & \$18559_copy_root_in_ram6634347_arg\(16 to 31) & \$18566\(32 to 47) & \$18559_copy_root_in_ram6634347_arg\(48 to 63) & \$18559_copy_root_in_ram6634347_arg\(64 to 79);
                state_var5923 := \$18571_COPY_ROOT_IN_RAM6634345\;
              when PAUSE_SET4708 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18612\ := eclat_unit;
                \$18566\ := eclat_resize(\$18559_copy_root_in_ram6634347_arg\(32 to 47),31) & eclat_false & 
                work.Int.add(\$18559_copy_root_in_ram6634347_arg\(32 to 47), 
                             work.Int.add(eclat_resize(work.Int.lsr(\$18599_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$v4707\ := \$ram_lock\;
                if \$v4707\(0) = '1' then
                  state_var5923 := Q_WAIT4706;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18559_copy_root_in_ram6634347_arg\(0 to 15)));
                  \$ram_write\ <= \$18566\(0 to 31); \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4705;
                end if;
              when PAUSE_SET4711 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18611\ := eclat_unit;
                \$v4710\ := \$ram_lock\;
                if \$v4710\(0) = '1' then
                  state_var5923 := Q_WAIT4709;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$18565\(0 to 30),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$18559_copy_root_in_ram6634347_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4708;
                end if;
              when PAUSE_SET4714 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18609\ := eclat_unit;
                \$18524_loop666_id\ := "000000010111";
                \$18524_loop666_arg\ := X"000" & X"1" & \$18559_copy_root_in_ram6634347_arg\(32 to 47) & eclat_resize(\$18565\(0 to 30),16) & eclat_resize(
                work.Int.lsr(\$18599_hd\(0 to 30), X"0000000" & X"2"),16);
                state_var5923 := \$18524_LOOP666\;
              when PAUSE_SET4732 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18633\ := eclat_unit;
                \$18634\ := work.Print.print_string(clk,of_string(" next="));
                \$18635\ := work.Int.print(clk,\$18632\(32 to 47));
                \$18636\ := work.Print.print_newline(clk,eclat_unit);
                \$18625_copy_root_in_ram6634345_arg\ := work.Int.add(
                                                        \$18625_copy_root_in_ram6634345_arg\(0 to 15), X"000" & X"1") & \$18625_copy_root_in_ram6634345_arg\(16 to 31) & \$18632\(32 to 47) & \$18625_copy_root_in_ram6634345_arg\(48 to 63) & \$18625_copy_root_in_ram6634345_arg\(64 to 79);
                state_var5923 := \$18625_COPY_ROOT_IN_RAM6634345\;
              when PAUSE_SET4735 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18651\ := eclat_unit;
                \$18632\ := eclat_resize(\$18625_copy_root_in_ram6634345_arg\(32 to 47),31) & eclat_false & 
                work.Int.add(\$18625_copy_root_in_ram6634345_arg\(32 to 47), 
                             work.Int.add(eclat_resize(work.Int.lsr(\$18638_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$v4734\ := \$ram_lock\;
                if \$v4734\(0) = '1' then
                  state_var5923 := Q_WAIT4733;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18625_copy_root_in_ram6634345_arg\(0 to 15)));
                  \$ram_write\ <= \$18632\(0 to 31); \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4732;
                end if;
              when PAUSE_SET4738 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18650\ := eclat_unit;
                \$v4737\ := \$ram_lock\;
                if \$v4737\(0) = '1' then
                  state_var5923 := Q_WAIT4736;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$18631\(0 to 30),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$18625_copy_root_in_ram6634345_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4735;
                end if;
              when PAUSE_SET4741 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18648\ := eclat_unit;
                \$18524_loop666_id\ := "000000011001";
                \$18524_loop666_arg\ := X"000" & X"1" & \$18625_copy_root_in_ram6634345_arg\(32 to 47) & eclat_resize(\$18631\(0 to 30),16) & eclat_resize(
                work.Int.lsr(\$18638_hd\(0 to 30), X"0000000" & X"2"),16);
                state_var5923 := \$18524_LOOP666\;
              when PAUSE_SET4756 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18621\ := eclat_unit;
                \$18622\ := work.Print.print_string(clk,of_string(" next="));
                \$18623\ := work.Int.print(clk,\$18620\(32 to 47));
                \$18624\ := work.Print.print_newline(clk,eclat_unit);
                \$18625_copy_root_in_ram6634345_id\ := "000000011010";
                \$18625_copy_root_in_ram6634345_arg\ := work.Int.add(
                                                        \$18613_copy_root_in_ram6634346_arg\(0 to 15), X"000" & X"1") & \$18613_copy_root_in_ram6634346_arg\(16 to 31) & \$18620\(32 to 47) & \$18613_copy_root_in_ram6634346_arg\(48 to 63) & \$18613_copy_root_in_ram6634346_arg\(64 to 79);
                state_var5923 := \$18625_COPY_ROOT_IN_RAM6634345\;
              when PAUSE_SET4759 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18666\ := eclat_unit;
                \$18620\ := eclat_resize(\$18613_copy_root_in_ram6634346_arg\(32 to 47),31) & eclat_false & 
                work.Int.add(\$18613_copy_root_in_ram6634346_arg\(32 to 47), 
                             work.Int.add(eclat_resize(work.Int.lsr(\$18653_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$v4758\ := \$ram_lock\;
                if \$v4758\(0) = '1' then
                  state_var5923 := Q_WAIT4757;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18613_copy_root_in_ram6634346_arg\(0 to 15)));
                  \$ram_write\ <= \$18620\(0 to 31); \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4756;
                end if;
              when PAUSE_SET4762 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18665\ := eclat_unit;
                \$v4761\ := \$ram_lock\;
                if \$v4761\(0) = '1' then
                  state_var5923 := Q_WAIT4760;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$18619\(0 to 30),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$18613_copy_root_in_ram6634346_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4759;
                end if;
              when PAUSE_SET4765 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18663\ := eclat_unit;
                \$18524_loop666_id\ := "000000011011";
                \$18524_loop666_arg\ := X"000" & X"1" & \$18613_copy_root_in_ram6634346_arg\(32 to 47) & eclat_resize(\$18619\(0 to 30),16) & eclat_resize(
                work.Int.lsr(\$18653_hd\(0 to 30), X"0000000" & X"2"),16);
                state_var5923 := \$18524_LOOP666\;
              when PAUSE_SET4780 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18681\ := eclat_unit;
                \$18533\ := eclat_resize(\$18532\(32 to 47),31) & eclat_false & 
                work.Int.add(\$18532\(32 to 47), work.Int.add(eclat_resize(
                                                              work.Int.lsr(
                                                              \$18668_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$18613_copy_root_in_ram6634346_id\ := "000000011100";
                \$18613_copy_root_in_ram6634346_arg\ := X"0" & X"3e8" & \$18468_wait662_arg\(65 to 80) & \$18533\(32 to 47) & \$18520\(96 to 111) & \$18520\(112 to 127);
                state_var5923 := \$18613_COPY_ROOT_IN_RAM6634346\;
              when PAUSE_SET4783 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18680\ := eclat_unit;
                \$v4782\ := \$ram_lock\;
                if \$v4782\(0) = '1' then
                  state_var5923 := Q_WAIT4781;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$18468_wait662_arg\(33 to 63),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$18532\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4780;
                end if;
              when PAUSE_SET4786 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18678\ := eclat_unit;
                \$18524_loop666_id\ := "000000011101";
                \$18524_loop666_arg\ := X"000" & X"1" & \$18532\(32 to 47) & eclat_resize(\$18468_wait662_arg\(33 to 63),16) & eclat_resize(
                work.Int.lsr(\$18668_hd\(0 to 30), X"0000000" & X"2"),16);
                state_var5923 := \$18524_LOOP666\;
              when PAUSE_SET4797 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18696\ := eclat_unit;
                \$18532\ := eclat_resize(\$18520\(112 to 127),31) & eclat_false & 
                work.Int.add(\$18520\(112 to 127), work.Int.add(eclat_resize(
                                                                work.Int.lsr(
                                                                \$18683_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$v4796\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$18468_wait662_arg\(64)) & 
                                           eclat_if(work.Int.le(\$18520\(96 to 111), eclat_resize(\$18468_wait662_arg\(33 to 63),16)) & 
                                           work.Int.lt(eclat_resize(\$18468_wait662_arg\(33 to 63),16), 
                                                       work.Int.add(\$18520\(96 to 111), X"1770")) & eclat_false) & eclat_false));
                if \$v4796\(0) = '1' then
                  \$18533\ := \$18468_wait662_arg\(33 to 64) & \$18532\(32 to 47);
                  \$18613_copy_root_in_ram6634346_id\ := "000000011100";
                  \$18613_copy_root_in_ram6634346_arg\ := X"0" & X"3e8" & \$18468_wait662_arg\(65 to 80) & \$18533\(32 to 47) & \$18520\(96 to 111) & \$18520\(112 to 127);
                  state_var5923 := \$18613_COPY_ROOT_IN_RAM6634346\;
                else
                  \$v4795\ := \$ram_lock\;
                  if \$v4795\(0) = '1' then
                    state_var5923 := Q_WAIT4794;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18468_wait662_arg\(33 to 63),16), X"000" & X"1")));
                    state_var5923 := PAUSE_GET4793;
                  end if;
                end if;
              when PAUSE_SET4800 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18695\ := eclat_unit;
                \$v4799\ := \$ram_lock\;
                if \$v4799\(0) = '1' then
                  state_var5923 := Q_WAIT4798;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$18468_wait662_arg\(1 to 31),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$18520\(112 to 127),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4797;
                end if;
              when PAUSE_SET4803 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18693\ := eclat_unit;
                \$18524_loop666_id\ := "000000011110";
                \$18524_loop666_arg\ := X"000" & X"1" & \$18520\(112 to 127) & eclat_resize(\$18468_wait662_arg\(1 to 31),16) & eclat_resize(
                work.Int.lsr(\$18683_hd\(0 to 30), X"0000000" & X"2"),16);
                state_var5923 := \$18524_LOOP666\;
              when Q_WAIT4611 =>
                \$v4612\ := \$ram_lock\;
                if \$v4612\(0) = '1' then
                  state_var5923 := Q_WAIT4611;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$18521_loop666_arg\(16 to 31), \$18521_loop666_arg\(0 to 15))));
                  \$ram_write\ <= \$18761\; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4610;
                end if;
              when Q_WAIT4614 =>
                \$v4615\ := \$ram_lock\;
                if \$v4615\(0) = '1' then
                  state_var5923 := Q_WAIT4614;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$18521_loop666_arg\(32 to 47), \$18521_loop666_arg\(0 to 15))));
                  state_var5923 := PAUSE_GET4613;
                end if;
              when Q_WAIT4618 =>
                \$v4619\ := \$ram_lock\;
                if \$v4619\(0) = '1' then
                  state_var5923 := Q_WAIT4618;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$18522_loop665_arg\(64 to 79), \$18522_loop665_arg\(0 to 15))));
                  \$ram_write\ <= \$18742\(0 to 31); \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4617;
                end if;
              when Q_WAIT4621 =>
                \$v4622\ := \$ram_lock\;
                if \$v4622\(0) = '1' then
                  state_var5923 := Q_WAIT4621;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$18741\(0 to 30),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$18522_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4620;
                end if;
              when Q_WAIT4624 =>
                \$v4625\ := \$ram_lock\;
                if \$v4625\(0) = '1' then
                  state_var5923 := Q_WAIT4624;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18741\(0 to 30),16)));
                  \$ram_write\ <= eclat_resize(\$18522_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4623;
                end if;
              when Q_WAIT4627 =>
                \$v4628\ := \$ram_lock\;
                if \$v4628\(0) = '1' then
                  state_var5923 := Q_WAIT4627;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18522_loop665_arg\(16 to 31)));
                  \$ram_write\ <= \$18745_hd\; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4626;
                end if;
              when Q_WAIT4630 =>
                \$v4631\ := \$ram_lock\;
                if \$v4631\(0) = '1' then
                  state_var5923 := Q_WAIT4630;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18741\(0 to 30),16)));
                  state_var5923 := PAUSE_GET4629;
                end if;
              when Q_WAIT4634 =>
                \$v4635\ := \$ram_lock\;
                if \$v4635\(0) = '1' then
                  state_var5923 := Q_WAIT4634;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18741\(0 to 30),16), X"000" & X"1")));
                  state_var5923 := PAUSE_GET4633;
                end if;
              when Q_WAIT4638 =>
                \$v4639\ := \$ram_lock\;
                if \$v4639\(0) = '1' then
                  state_var5923 := Q_WAIT4638;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$18522_loop665_arg\(64 to 79), \$18522_loop665_arg\(0 to 15))));
                  state_var5923 := PAUSE_GET4637;
                end if;
              when Q_WAIT4642 =>
                \$v4643\ := \$ram_lock\;
                if \$v4643\(0) = '1' then
                  state_var5923 := Q_WAIT4642;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(\$18523_aux664_arg\(0 to 15)));
                  state_var5923 := PAUSE_GET4641;
                end if;
              when Q_WAIT4646 =>
                \$v4647\ := \$ram_lock\;
                if \$v4647\(0) = '1' then
                  state_var5923 := Q_WAIT4646;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$18524_loop666_arg\(16 to 31), \$18524_loop666_arg\(0 to 15))));
                  \$ram_write\ <= \$18728\; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4645;
                end if;
              when Q_WAIT4649 =>
                \$v4650\ := \$ram_lock\;
                if \$v4650\(0) = '1' then
                  state_var5923 := Q_WAIT4649;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$18524_loop666_arg\(32 to 47), \$18524_loop666_arg\(0 to 15))));
                  state_var5923 := PAUSE_GET4648;
                end if;
              when Q_WAIT4653 =>
                \$v4654\ := \$ram_lock\;
                if \$v4654\(0) = '1' then
                  state_var5923 := Q_WAIT4653;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$18525_loop665_arg\(64 to 79), \$18525_loop665_arg\(0 to 15))));
                  \$ram_write\ <= \$18709\(0 to 31); \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4652;
                end if;
              when Q_WAIT4656 =>
                \$v4657\ := \$ram_lock\;
                if \$v4657\(0) = '1' then
                  state_var5923 := Q_WAIT4656;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$18708\(0 to 30),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$18525_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4655;
                end if;
              when Q_WAIT4659 =>
                \$v4660\ := \$ram_lock\;
                if \$v4660\(0) = '1' then
                  state_var5923 := Q_WAIT4659;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18708\(0 to 30),16)));
                  \$ram_write\ <= eclat_resize(\$18525_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4658;
                end if;
              when Q_WAIT4662 =>
                \$v4663\ := \$ram_lock\;
                if \$v4663\(0) = '1' then
                  state_var5923 := Q_WAIT4662;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18525_loop665_arg\(16 to 31)));
                  \$ram_write\ <= \$18712_hd\; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4661;
                end if;
              when Q_WAIT4665 =>
                \$v4666\ := \$ram_lock\;
                if \$v4666\(0) = '1' then
                  state_var5923 := Q_WAIT4665;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18708\(0 to 30),16)));
                  state_var5923 := PAUSE_GET4664;
                end if;
              when Q_WAIT4669 =>
                \$v4670\ := \$ram_lock\;
                if \$v4670\(0) = '1' then
                  state_var5923 := Q_WAIT4669;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18708\(0 to 30),16), X"000" & X"1")));
                  state_var5923 := PAUSE_GET4668;
                end if;
              when Q_WAIT4673 =>
                \$v4674\ := \$ram_lock\;
                if \$v4674\(0) = '1' then
                  state_var5923 := Q_WAIT4673;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$18525_loop665_arg\(64 to 79), \$18525_loop665_arg\(0 to 15))));
                  state_var5923 := PAUSE_GET4672;
                end if;
              when Q_WAIT4677 =>
                \$v4678\ := \$ram_lock\;
                if \$v4678\(0) = '1' then
                  state_var5923 := Q_WAIT4677;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(\$18526_aux664_arg\(0 to 15)));
                  state_var5923 := PAUSE_GET4676;
                end if;
              when Q_WAIT4682 =>
                \$v4683\ := \$ram_lock\;
                if \$v4683\(0) = '1' then
                  state_var5923 := Q_WAIT4682;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18571_copy_root_in_ram6634345_arg\(0 to 15)));
                  \$ram_write\ <= \$18578\(0 to 31); \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4681;
                end if;
              when Q_WAIT4685 =>
                \$v4686\ := \$ram_lock\;
                if \$v4686\(0) = '1' then
                  state_var5923 := Q_WAIT4685;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$18577\(0 to 30),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$18571_copy_root_in_ram6634345_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4684;
                end if;
              when Q_WAIT4688 =>
                \$v4689\ := \$ram_lock\;
                if \$v4689\(0) = '1' then
                  state_var5923 := Q_WAIT4688;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18577\(0 to 30),16)));
                  \$ram_write\ <= eclat_resize(\$18571_copy_root_in_ram6634345_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4687;
                end if;
              when Q_WAIT4691 =>
                \$v4692\ := \$ram_lock\;
                if \$v4692\(0) = '1' then
                  state_var5923 := Q_WAIT4691;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18571_copy_root_in_ram6634345_arg\(32 to 47)));
                  \$ram_write\ <= \$18584_hd\; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4690;
                end if;
              when Q_WAIT4694 =>
                \$v4695\ := \$ram_lock\;
                if \$v4695\(0) = '1' then
                  state_var5923 := Q_WAIT4694;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18577\(0 to 30),16)));
                  state_var5923 := PAUSE_GET4693;
                end if;
              when Q_WAIT4698 =>
                \$v4699\ := \$ram_lock\;
                if \$v4699\(0) = '1' then
                  state_var5923 := Q_WAIT4698;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18577\(0 to 30),16), X"000" & X"1")));
                  state_var5923 := PAUSE_GET4697;
                end if;
              when Q_WAIT4702 =>
                \$v4703\ := \$ram_lock\;
                if \$v4703\(0) = '1' then
                  state_var5923 := Q_WAIT4702;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(\$18571_copy_root_in_ram6634345_arg\(0 to 15)));
                  state_var5923 := PAUSE_GET4701;
                end if;
              when Q_WAIT4706 =>
                \$v4707\ := \$ram_lock\;
                if \$v4707\(0) = '1' then
                  state_var5923 := Q_WAIT4706;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18559_copy_root_in_ram6634347_arg\(0 to 15)));
                  \$ram_write\ <= \$18566\(0 to 31); \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4705;
                end if;
              when Q_WAIT4709 =>
                \$v4710\ := \$ram_lock\;
                if \$v4710\(0) = '1' then
                  state_var5923 := Q_WAIT4709;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$18565\(0 to 30),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$18559_copy_root_in_ram6634347_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4708;
                end if;
              when Q_WAIT4712 =>
                \$v4713\ := \$ram_lock\;
                if \$v4713\(0) = '1' then
                  state_var5923 := Q_WAIT4712;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18565\(0 to 30),16)));
                  \$ram_write\ <= eclat_resize(\$18559_copy_root_in_ram6634347_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4711;
                end if;
              when Q_WAIT4715 =>
                \$v4716\ := \$ram_lock\;
                if \$v4716\(0) = '1' then
                  state_var5923 := Q_WAIT4715;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18559_copy_root_in_ram6634347_arg\(32 to 47)));
                  \$ram_write\ <= \$18599_hd\; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4714;
                end if;
              when Q_WAIT4718 =>
                \$v4719\ := \$ram_lock\;
                if \$v4719\(0) = '1' then
                  state_var5923 := Q_WAIT4718;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18565\(0 to 30),16)));
                  state_var5923 := PAUSE_GET4717;
                end if;
              when Q_WAIT4722 =>
                \$v4723\ := \$ram_lock\;
                if \$v4723\(0) = '1' then
                  state_var5923 := Q_WAIT4722;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18565\(0 to 30),16), X"000" & X"1")));
                  state_var5923 := PAUSE_GET4721;
                end if;
              when Q_WAIT4726 =>
                \$v4727\ := \$ram_lock\;
                if \$v4727\(0) = '1' then
                  state_var5923 := Q_WAIT4726;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(\$18559_copy_root_in_ram6634347_arg\(0 to 15)));
                  state_var5923 := PAUSE_GET4725;
                end if;
              when Q_WAIT4730 =>
                \$v4731\ := \$global_end_lock\;
                if \$v4731\(0) = '1' then
                  state_var5923 := Q_WAIT4730;
                else
                  acquire(\$global_end_lock\);
                  \$global_end_ptr\ <= 0;
                  state_var5923 := PAUSE_GET4729;
                end if;
              when Q_WAIT4733 =>
                \$v4734\ := \$ram_lock\;
                if \$v4734\(0) = '1' then
                  state_var5923 := Q_WAIT4733;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18625_copy_root_in_ram6634345_arg\(0 to 15)));
                  \$ram_write\ <= \$18632\(0 to 31); \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4732;
                end if;
              when Q_WAIT4736 =>
                \$v4737\ := \$ram_lock\;
                if \$v4737\(0) = '1' then
                  state_var5923 := Q_WAIT4736;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$18631\(0 to 30),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$18625_copy_root_in_ram6634345_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4735;
                end if;
              when Q_WAIT4739 =>
                \$v4740\ := \$ram_lock\;
                if \$v4740\(0) = '1' then
                  state_var5923 := Q_WAIT4739;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18631\(0 to 30),16)));
                  \$ram_write\ <= eclat_resize(\$18625_copy_root_in_ram6634345_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4738;
                end if;
              when Q_WAIT4742 =>
                \$v4743\ := \$ram_lock\;
                if \$v4743\(0) = '1' then
                  state_var5923 := Q_WAIT4742;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18625_copy_root_in_ram6634345_arg\(32 to 47)));
                  \$ram_write\ <= \$18638_hd\; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4741;
                end if;
              when Q_WAIT4745 =>
                \$v4746\ := \$ram_lock\;
                if \$v4746\(0) = '1' then
                  state_var5923 := Q_WAIT4745;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18631\(0 to 30),16)));
                  state_var5923 := PAUSE_GET4744;
                end if;
              when Q_WAIT4749 =>
                \$v4750\ := \$ram_lock\;
                if \$v4750\(0) = '1' then
                  state_var5923 := Q_WAIT4749;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18631\(0 to 30),16), X"000" & X"1")));
                  state_var5923 := PAUSE_GET4748;
                end if;
              when Q_WAIT4753 =>
                \$v4754\ := \$ram_lock\;
                if \$v4754\(0) = '1' then
                  state_var5923 := Q_WAIT4753;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(\$18625_copy_root_in_ram6634345_arg\(0 to 15)));
                  state_var5923 := PAUSE_GET4752;
                end if;
              when Q_WAIT4757 =>
                \$v4758\ := \$ram_lock\;
                if \$v4758\(0) = '1' then
                  state_var5923 := Q_WAIT4757;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18613_copy_root_in_ram6634346_arg\(0 to 15)));
                  \$ram_write\ <= \$18620\(0 to 31); \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4756;
                end if;
              when Q_WAIT4760 =>
                \$v4761\ := \$ram_lock\;
                if \$v4761\(0) = '1' then
                  state_var5923 := Q_WAIT4760;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$18619\(0 to 30),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$18613_copy_root_in_ram6634346_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4759;
                end if;
              when Q_WAIT4763 =>
                \$v4764\ := \$ram_lock\;
                if \$v4764\(0) = '1' then
                  state_var5923 := Q_WAIT4763;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18619\(0 to 30),16)));
                  \$ram_write\ <= eclat_resize(\$18613_copy_root_in_ram6634346_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4762;
                end if;
              when Q_WAIT4766 =>
                \$v4767\ := \$ram_lock\;
                if \$v4767\(0) = '1' then
                  state_var5923 := Q_WAIT4766;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18613_copy_root_in_ram6634346_arg\(32 to 47)));
                  \$ram_write\ <= \$18653_hd\; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4765;
                end if;
              when Q_WAIT4769 =>
                \$v4770\ := \$ram_lock\;
                if \$v4770\(0) = '1' then
                  state_var5923 := Q_WAIT4769;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18619\(0 to 30),16)));
                  state_var5923 := PAUSE_GET4768;
                end if;
              when Q_WAIT4773 =>
                \$v4774\ := \$ram_lock\;
                if \$v4774\(0) = '1' then
                  state_var5923 := Q_WAIT4773;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18619\(0 to 30),16), X"000" & X"1")));
                  state_var5923 := PAUSE_GET4772;
                end if;
              when Q_WAIT4777 =>
                \$v4778\ := \$ram_lock\;
                if \$v4778\(0) = '1' then
                  state_var5923 := Q_WAIT4777;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(\$18613_copy_root_in_ram6634346_arg\(0 to 15)));
                  state_var5923 := PAUSE_GET4776;
                end if;
              when Q_WAIT4781 =>
                \$v4782\ := \$ram_lock\;
                if \$v4782\(0) = '1' then
                  state_var5923 := Q_WAIT4781;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$18468_wait662_arg\(33 to 63),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$18532\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4780;
                end if;
              when Q_WAIT4784 =>
                \$v4785\ := \$ram_lock\;
                if \$v4785\(0) = '1' then
                  state_var5923 := Q_WAIT4784;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18468_wait662_arg\(33 to 63),16)));
                  \$ram_write\ <= eclat_resize(\$18532\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4783;
                end if;
              when Q_WAIT4787 =>
                \$v4788\ := \$ram_lock\;
                if \$v4788\(0) = '1' then
                  state_var5923 := Q_WAIT4787;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18532\(32 to 47)));
                  \$ram_write\ <= \$18668_hd\; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4786;
                end if;
              when Q_WAIT4790 =>
                \$v4791\ := \$ram_lock\;
                if \$v4791\(0) = '1' then
                  state_var5923 := Q_WAIT4790;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18468_wait662_arg\(33 to 63),16)));
                  state_var5923 := PAUSE_GET4789;
                end if;
              when Q_WAIT4794 =>
                \$v4795\ := \$ram_lock\;
                if \$v4795\(0) = '1' then
                  state_var5923 := Q_WAIT4794;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18468_wait662_arg\(33 to 63),16), X"000" & X"1")));
                  state_var5923 := PAUSE_GET4793;
                end if;
              when Q_WAIT4798 =>
                \$v4799\ := \$ram_lock\;
                if \$v4799\(0) = '1' then
                  state_var5923 := Q_WAIT4798;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$18468_wait662_arg\(1 to 31),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$18520\(112 to 127),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4797;
                end if;
              when Q_WAIT4801 =>
                \$v4802\ := \$ram_lock\;
                if \$v4802\(0) = '1' then
                  state_var5923 := Q_WAIT4801;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18468_wait662_arg\(1 to 31),16)));
                  \$ram_write\ <= eclat_resize(\$18520\(112 to 127),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4800;
                end if;
              when Q_WAIT4804 =>
                \$v4805\ := \$ram_lock\;
                if \$v4805\(0) = '1' then
                  state_var5923 := Q_WAIT4804;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18520\(112 to 127)));
                  \$ram_write\ <= \$18683_hd\; \$ram_write_request\ <= '1';
                  state_var5923 := PAUSE_SET4803;
                end if;
              when Q_WAIT4807 =>
                \$v4808\ := \$ram_lock\;
                if \$v4808\(0) = '1' then
                  state_var5923 := Q_WAIT4807;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18468_wait662_arg\(1 to 31),16)));
                  state_var5923 := PAUSE_GET4806;
                end if;
              when Q_WAIT4811 =>
                \$v4812\ := \$ram_lock\;
                if \$v4812\(0) = '1' then
                  state_var5923 := Q_WAIT4811;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18468_wait662_arg\(1 to 31),16), X"000" & X"1")));
                  state_var5923 := PAUSE_GET4810;
                end if;
              when IDLE4609 =>
                rdy4608 := eclat_false;
                \$v4814\ := work.Int.gt(work.Int.add(\$18520\(80 to 95), \$18468_wait662_arg\(81 to 96)), 
                                        work.Int.add(\$18520\(96 to 111), X"1770"));
                if \$v4814\(0) = '1' then
                  \$18527\ := work.Print.print_newline(clk,eclat_unit);
                  \$18528\ := work.Print.print_newline(clk,eclat_unit);
                  \$18529\ := work.Print.print_string(clk,of_string("[================= GC START ======================]"));
                  \$18530\ := work.Print.print_newline(clk,eclat_unit);
                  \$18531\ := work.Print.print_newline(clk,eclat_unit);
                  \$v4813\ := work.Bool.lnot(eclat_if(work.Bool.lnot(
                                                      ""&\$18468_wait662_arg\(32)) & 
                                             eclat_if(work.Int.le(\$18520\(96 to 111), eclat_resize(\$18468_wait662_arg\(1 to 31),16)) & 
                                             work.Int.lt(eclat_resize(\$18468_wait662_arg\(1 to 31),16), 
                                                         work.Int.add(
                                                         \$18520\(96 to 111), X"1770")) & eclat_false) & eclat_false));
                  if \$v4813\(0) = '1' then
                    \$18532\ := \$18468_wait662_arg\(1 to 32) & \$18520\(112 to 127);
                    \$v4796\ := work.Bool.lnot(eclat_if(work.Bool.lnot(
                                                        ""&\$18468_wait662_arg\(64)) & 
                                               eclat_if(work.Int.le(\$18520\(96 to 111), eclat_resize(\$18468_wait662_arg\(33 to 63),16)) & 
                                               work.Int.lt(eclat_resize(\$18468_wait662_arg\(33 to 63),16), 
                                                           work.Int.add(
                                                           \$18520\(96 to 111), X"1770")) & eclat_false) & eclat_false));
                    if \$v4796\(0) = '1' then
                      \$18533\ := \$18468_wait662_arg\(33 to 64) & \$18532\(32 to 47);
                      \$18613_copy_root_in_ram6634346_id\ := "000000011100";
                      \$18613_copy_root_in_ram6634346_arg\ := X"0" & X"3e8" & \$18468_wait662_arg\(65 to 80) & \$18533\(32 to 47) & \$18520\(96 to 111) & \$18520\(112 to 127);
                      state_var5923 := \$18613_COPY_ROOT_IN_RAM6634346\;
                    else
                      \$v4795\ := \$ram_lock\;
                      if \$v4795\(0) = '1' then
                        state_var5923 := Q_WAIT4794;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$18468_wait662_arg\(33 to 63),16), X"000" & X"1")));
                        state_var5923 := PAUSE_GET4793;
                      end if;
                    end if;
                  else
                    \$v4812\ := \$ram_lock\;
                    if \$v4812\(0) = '1' then
                      state_var5923 := Q_WAIT4811;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                        eclat_resize(\$18468_wait662_arg\(1 to 31),16), X"000" & X"1")));
                      state_var5923 := PAUSE_GET4810;
                    end if;
                  end if;
                else
                  result4607 := \$18468_wait662_arg\(1 to 32) & \$18468_wait662_arg\(33 to 64) & \$18520\(80 to 95) & 
                  work.Int.add(\$18520\(80 to 95), \$18468_wait662_arg\(81 to 96)) & \$18520\(96 to 111) & \$18520\(112 to 127);
                  rdy4608 := eclat_true;
                  state_var5923 := IDLE4609;
                end if;
              end case;
              
              if rdy4608(0) = '1' then
                
              else
                result4607 := \$18520\(0 to 31) & \$18520\(32 to 63) & \$18520\(64 to 79) & \$18520\(80 to 95) & \$18520\(96 to 111) & \$18520\(112 to 127);
              end if;
              \$18520\ := result4607 & rdy4608;
              \$18519\ := \$18520\;
              \$v4606\ := ""&\$18519\(128);
              if \$v4606\(0) = '1' then
                \$18468_wait662_result\ := \$18519\(0 to 31) & \$18519\(32 to 63) & \$18519\(64 to 79);
                \$18512\ := \$18468_wait662_result\;
                \$18513\ := work.Print.print_string(clk,of_string("size:"));
                \$18514\ := work.Int.print(clk,eclat_if(work.Int.eq(\$18469_make_block579_arg\(112 to 127), X"000" & X"0") & X"000" & X"1" & \$18469_make_block579_arg\(112 to 127)));
                \$18515\ := work.Print.print_newline(clk,eclat_unit);
                \$v4818\ := \$ram_lock\;
                if \$v4818\(0) = '1' then
                  state_var5922 := Q_WAIT4817;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18512\(64 to 79)));
                  \$ram_write\ <= work.Int.lor(work.Int.lsl(eclat_resize(\$18469_make_block579_arg\(80 to 111),31), X"000000" & X"18"), 
                                               work.Int.lsl(eclat_resize(
                                                            eclat_if(
                                                            work.Int.eq(
                                                            \$18469_make_block579_arg\(112 to 127), X"000" & X"0") & X"000" & X"1" & \$18469_make_block579_arg\(112 to 127)),31), X"0000000" & X"2")) & eclat_true; \$ram_write_request\ <= '1';
                  state_var5922 := PAUSE_SET4816;
                end if;
              else
                \$18468_wait662_arg\ := eclat_unit & \$18468_wait662_arg\(1 to 32) & \$18468_wait662_arg\(33 to 64) & \$18468_wait662_arg\(65 to 80) & \$18468_wait662_arg\(81 to 96);
                state_var5922 := \$18468_WAIT662\;
              end if;
            when \$18469_MAKE_BLOCK579\ =>
              \$18508\ := work.Print.print_string(clk,of_string("GC-ALLOC:(size="));
              \$18509\ := work.Int.print(clk,work.Int.add(eclat_if(work.Int.eq(
                                                                   \$18469_make_block579_arg\(112 to 127), X"000" & X"0") & X"000" & X"1" & \$18469_make_block579_arg\(112 to 127)), X"000" & X"1"));
              \$18510\ := work.Print.print_string(clk,of_string(")"));
              \$18511\ := work.Print.print_newline(clk,eclat_unit);
              \$18468_wait662_id\ := "000000011111";
              \$18468_wait662_arg\ := eclat_unit & \$18469_make_block579_arg\(16 to 47) & \$18469_make_block579_arg\(48 to 79) & \$18469_make_block579_arg\(0 to 15) & 
              work.Int.add(eclat_if(work.Int.eq(\$18469_make_block579_arg\(112 to 127), X"000" & X"0") & X"000" & X"1" & \$18469_make_block579_arg\(112 to 127)), X"000" & X"1");
              state_var5922 := \$18468_WAIT662\;
            when PAUSE_GET4578 =>
              \$18785\ := \$ram_value\;
              release(\$ram_lock\);
              \$v4577\ := \$ram_lock\;
              if \$v4577\(0) = '1' then
                state_var5922 := Q_WAIT4576;
              else
                acquire(\$ram_lock\);
                \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                        \$18466_loop666_arg\(16 to 31), \$18466_loop666_arg\(0 to 15))));
                \$ram_write\ <= \$18785\; \$ram_write_request\ <= '1';
                state_var5922 := PAUSE_SET4575;
              end if;
            when PAUSE_GET4594 =>
              \$18769_hd\ := \$ram_value\;
              release(\$ram_lock\);
              \$18770\ := work.Print.print_string(clk,of_string("bloc "));
              \$18771\ := work.Int.print(clk,eclat_resize(\$18765\(0 to 30),16));
              \$18772\ := work.Print.print_string(clk,of_string(" of size "));
              \$18773\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                          work.Int.lsr(
                                                          \$18769_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
              \$18774\ := work.Print.print_string(clk,of_string(" from "));
              \$18775\ := work.Int.print(clk,eclat_resize(\$18765\(0 to 30),16));
              \$18776\ := work.Print.print_string(clk,of_string(" to "));
              \$18777\ := work.Int.print(clk,\$18467_loop665_arg\(16 to 31));
              \$18778\ := work.Print.print_newline(clk,eclat_unit);
              \$v4593\ := \$ram_lock\;
              if \$v4593\(0) = '1' then
                state_var5922 := Q_WAIT4592;
              else
                acquire(\$ram_lock\);
                \$ram_ptr_write\ <= to_integer(unsigned(\$18467_loop665_arg\(16 to 31)));
                \$ram_write\ <= \$18769_hd\; \$ram_write_request\ <= '1';
                state_var5922 := PAUSE_SET4591;
              end if;
            when PAUSE_GET4598 =>
              \$18768_w\ := \$ram_value\;
              release(\$ram_lock\);
              \$v4597\ := eclat_if(work.Bool.lnot(""&\$18768_w\(31)) & 
                          eclat_if(work.Int.le(\$18467_loop665_arg\(48 to 63), eclat_resize(\$18768_w\(0 to 30),16)) & 
                          work.Int.lt(eclat_resize(\$18768_w\(0 to 30),16), 
                                      work.Int.add(\$18467_loop665_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false);
              if \$v4597\(0) = '1' then
                \$18766\ := \$18768_w\ & \$18467_loop665_arg\(16 to 31);
                \$v4584\ := \$ram_lock\;
                if \$v4584\(0) = '1' then
                  state_var5922 := Q_WAIT4583;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$18467_loop665_arg\(64 to 79), \$18467_loop665_arg\(0 to 15))));
                  \$ram_write\ <= \$18766\(0 to 31); \$ram_write_request\ <= '1';
                  state_var5922 := PAUSE_SET4582;
                end if;
              else
                \$v4596\ := \$ram_lock\;
                if \$v4596\(0) = '1' then
                  state_var5922 := Q_WAIT4595;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18765\(0 to 30),16)));
                  state_var5922 := PAUSE_GET4594;
                end if;
              end if;
            when PAUSE_GET4602 =>
              \$18765\ := \$ram_value\;
              release(\$ram_lock\);
              \$v4601\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$18765\(31)) & 
                                         eclat_if(work.Int.le(\$18467_loop665_arg\(32 to 47), eclat_resize(\$18765\(0 to 30),16)) & 
                                         work.Int.lt(eclat_resize(\$18765\(0 to 30),16), 
                                                     work.Int.add(\$18467_loop665_arg\(32 to 47), X"1770")) & eclat_false) & eclat_false));
              if \$v4601\(0) = '1' then
                \$18766\ := \$18765\ & \$18467_loop665_arg\(16 to 31);
                \$v4584\ := \$ram_lock\;
                if \$v4584\(0) = '1' then
                  state_var5922 := Q_WAIT4583;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$18467_loop665_arg\(64 to 79), \$18467_loop665_arg\(0 to 15))));
                  \$ram_write\ <= \$18766\(0 to 31); \$ram_write_request\ <= '1';
                  state_var5922 := PAUSE_SET4582;
                end if;
              else
                \$v4600\ := \$ram_lock\;
                if \$v4600\(0) = '1' then
                  state_var5922 := Q_WAIT4599;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18765\(0 to 30),16), X"000" & X"1")));
                  state_var5922 := PAUSE_GET4598;
                end if;
              end if;
            when PAUSE_SET4575 =>
              \$ram_write_request\ <= '0';
              release(\$ram_lock\);
              \$18786\ := eclat_unit;
              \$18466_loop666_arg\ := work.Int.add(\$18466_loop666_arg\(0 to 15), X"000" & X"1") & \$18466_loop666_arg\(16 to 31) & \$18466_loop666_arg\(32 to 47) & \$18466_loop666_arg\(48 to 63);
              state_var5922 := \$18466_LOOP666\;
            when PAUSE_SET4582 =>
              \$ram_write_request\ <= '0';
              release(\$ram_lock\);
              \$18767\ := eclat_unit;
              \$18467_loop665_arg\ := work.Int.add(\$18467_loop665_arg\(0 to 15), X"000" & X"1") & \$18766\(32 to 47) & \$18467_loop665_arg\(32 to 47) & \$18467_loop665_arg\(48 to 63) & \$18467_loop665_arg\(64 to 79) & \$18467_loop665_arg\(80 to 95);
              state_var5922 := \$18467_LOOP665\;
            when PAUSE_SET4585 =>
              \$ram_write_request\ <= '0';
              release(\$ram_lock\);
              \$18782\ := eclat_unit;
              \$18766\ := eclat_resize(\$18467_loop665_arg\(16 to 31),31) & eclat_false & 
              work.Int.add(\$18467_loop665_arg\(16 to 31), work.Int.add(
                                                           eclat_resize(
                                                           work.Int.lsr(
                                                           \$18769_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
              \$v4584\ := \$ram_lock\;
              if \$v4584\(0) = '1' then
                state_var5922 := Q_WAIT4583;
              else
                acquire(\$ram_lock\);
                \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                        \$18467_loop665_arg\(64 to 79), \$18467_loop665_arg\(0 to 15))));
                \$ram_write\ <= \$18766\(0 to 31); \$ram_write_request\ <= '1';
                state_var5922 := PAUSE_SET4582;
              end if;
            when PAUSE_SET4588 =>
              \$ram_write_request\ <= '0';
              release(\$ram_lock\);
              \$18781\ := eclat_unit;
              \$v4587\ := \$ram_lock\;
              if \$v4587\(0) = '1' then
                state_var5922 := Q_WAIT4586;
              else
                acquire(\$ram_lock\);
                \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                        eclat_resize(\$18765\(0 to 30),16), X"000" & X"1")));
                \$ram_write\ <= eclat_resize(\$18467_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                state_var5922 := PAUSE_SET4585;
              end if;
            when PAUSE_SET4591 =>
              \$ram_write_request\ <= '0';
              release(\$ram_lock\);
              \$18779\ := eclat_unit;
              \$18466_loop666_id\ := "000000001101";
              \$18466_loop666_arg\ := X"000" & X"1" & \$18467_loop665_arg\(16 to 31) & eclat_resize(\$18765\(0 to 30),16) & eclat_resize(
              work.Int.lsr(\$18769_hd\(0 to 30), X"0000000" & X"2"),16);
              state_var5922 := \$18466_LOOP666\;
            when PAUSE_SET4816 =>
              \$ram_write_request\ <= '0';
              release(\$ram_lock\);
              \$18516\ := eclat_unit;
              \$18469_make_block579_result\ := \$18512\(0 to 31) & \$18512\(32 to 63) & eclat_resize(\$18512\(64 to 79),31) & eclat_false;
              state_var5922 := \$18469_MAKE_BLOCK579\;
            when PAUSE_SET4819 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18505\ := eclat_unit;
              result4572 := eclat_unit;
              rdy4573 := eclat_true;
              state_var5922 := IDLE4574;
            when PAUSE_SET4822 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18504\ := eclat_unit;
              \$v4821\ := \$code_lock\;
              if \$v4821\(0) = '1' then
                state_var5922 := Q_WAIT4820;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 34;\$code_write\ <= "000"& X"00000" & X"8f"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4819;
              end if;
            when PAUSE_SET4825 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18503\ := eclat_unit;
              \$v4824\ := \$code_lock\;
              if \$v4824\(0) = '1' then
                state_var5922 := Q_WAIT4823;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 33;\$code_write\ <= "000"& X"000000" & X"1"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4822;
              end if;
            when PAUSE_SET4828 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18502\ := eclat_unit;
              \$v4827\ := \$code_lock\;
              if \$v4827\(0) = '1' then
                state_var5922 := Q_WAIT4826;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 32;\$code_write\ <= "000"& X"00000" & X"13"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4825;
              end if;
            when PAUSE_SET4831 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18501\ := eclat_unit;
              \$v4830\ := \$code_lock\;
              if \$v4830\(0) = '1' then
                state_var5922 := Q_WAIT4829;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 31;\$code_write\ <= "000"& X"000000" & X"0"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4828;
              end if;
            when PAUSE_SET4834 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18500\ := eclat_unit;
              \$v4833\ := \$code_lock\;
              if \$v4833\(0) = '1' then
                state_var5922 := Q_WAIT4832;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 30;\$code_write\ <= "000"& X"00000" & X"5d"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4831;
              end if;
            when PAUSE_SET4837 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18499\ := eclat_unit;
              \$v4836\ := \$code_lock\;
              if \$v4836\(0) = '1' then
                state_var5922 := Q_WAIT4835;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 29;\$code_write\ <= "000"& X"00000" & X"21"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4834;
              end if;
            when PAUSE_SET4840 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18498\ := eclat_unit;
              \$v4839\ := \$code_lock\;
              if \$v4839\(0) = '1' then
                state_var5922 := Q_WAIT4838;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 28;\$code_write\ <= "000"& X"000000" & X"b"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4837;
              end if;
            when PAUSE_SET4843 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18497\ := eclat_unit;
              \$v4842\ := \$code_lock\;
              if \$v4842\(0) = '1' then
                state_var5922 := Q_WAIT4841;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 27;\$code_write\ <= "000"& X"000000" & X"b"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4840;
              end if;
            when PAUSE_SET4846 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18496\ := eclat_unit;
              \$v4845\ := \$code_lock\;
              if \$v4845\(0) = '1' then
                state_var5922 := Q_WAIT4844;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 26;\$code_write\ <= "000"& X"00000" & X"67"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4843;
              end if;
            when PAUSE_SET4849 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18495\ := eclat_unit;
              \$v4848\ := \$code_lock\;
              if \$v4848\(0) = '1' then
                state_var5922 := Q_WAIT4847;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 25;\$code_write\ <= work.Int.neg(
                                                         "000"& X"00000" & X"17"); \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4846;
              end if;
            when PAUSE_SET4852 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18494\ := eclat_unit;
              \$v4851\ := \$code_lock\;
              if \$v4851\(0) = '1' then
                state_var5922 := Q_WAIT4850;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 24;\$code_write\ <= "000"& X"000000" & X"0"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4849;
              end if;
            when PAUSE_SET4855 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18493\ := eclat_unit;
              \$v4854\ := \$code_lock\;
              if \$v4854\(0) = '1' then
                state_var5922 := Q_WAIT4853;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 23;\$code_write\ <= "000"& X"000000" & X"1"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4852;
              end if;
            when PAUSE_SET4858 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18492\ := eclat_unit;
              \$v4857\ := \$code_lock\;
              if \$v4857\(0) = '1' then
                state_var5922 := Q_WAIT4856;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 22;\$code_write\ <= "000"& X"00000" & X"2c"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4855;
              end if;
            when PAUSE_SET4861 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18491\ := eclat_unit;
              \$v4860\ := \$code_lock\;
              if \$v4860\(0) = '1' then
                state_var5922 := Q_WAIT4859;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 21;\$code_write\ <= "000"& X"000000" & X"1"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4858;
              end if;
            when PAUSE_SET4864 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18490\ := eclat_unit;
              \$v4863\ := \$code_lock\;
              if \$v4863\(0) = '1' then
                state_var5922 := Q_WAIT4862;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 20;\$code_write\ <= "000"& X"00000" & X"28"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4861;
              end if;
            when PAUSE_SET4867 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18489\ := eclat_unit;
              \$v4866\ := \$code_lock\;
              if \$v4866\(0) = '1' then
                state_var5922 := Q_WAIT4865;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 19;\$code_write\ <= "000"& X"00000" & X"6e"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4864;
              end if;
            when PAUSE_SET4870 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18488\ := eclat_unit;
              \$v4869\ := \$code_lock\;
              if \$v4869\(0) = '1' then
                state_var5922 := Q_WAIT4868;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 18;\$code_write\ <= "000"& X"00000" & X"21"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4867;
              end if;
            when PAUSE_SET4873 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18487\ := eclat_unit;
              \$v4872\ := \$code_lock\;
              if \$v4872\(0) = '1' then
                state_var5922 := Q_WAIT4871;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 17;\$code_write\ <= "000"& X"00000" & X"32"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4870;
              end if;
            when PAUSE_SET4876 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18486\ := eclat_unit;
              \$v4875\ := \$code_lock\;
              if \$v4875\(0) = '1' then
                state_var5922 := Q_WAIT4874;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 16;\$code_write\ <= work.Int.neg(
                                                         "000"& X"000000" & X"1"); \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4873;
              end if;
            when PAUSE_SET4879 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18485\ := eclat_unit;
              \$v4878\ := \$code_lock\;
              if \$v4878\(0) = '1' then
                state_var5922 := Q_WAIT4877;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 15;\$code_write\ <= "000"& X"00000" & X"7f"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4876;
              end if;
            when PAUSE_SET4882 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18484\ := eclat_unit;
              \$v4881\ := \$code_lock\;
              if \$v4881\(0) = '1' then
                state_var5922 := Q_WAIT4880;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 14;\$code_write\ <= "000"& X"000000" & X"b"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4879;
              end if;
            when PAUSE_SET4885 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18483\ := eclat_unit;
              \$v4884\ := \$code_lock\;
              if \$v4884\(0) = '1' then
                state_var5922 := Q_WAIT4883;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 13;\$code_write\ <= "000"& X"00000" & X"21"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4882;
              end if;
            when PAUSE_SET4888 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18482\ := eclat_unit;
              \$v4887\ := \$code_lock\;
              if \$v4887\(0) = '1' then
                state_var5922 := Q_WAIT4886;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 12;\$code_write\ <= "000"& X"00000" & X"32"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4885;
              end if;
            when PAUSE_SET4891 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18481\ := eclat_unit;
              \$v4890\ := \$code_lock\;
              if \$v4890\(0) = '1' then
                state_var5922 := Q_WAIT4889;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 11;\$code_write\ <= work.Int.neg(
                                                         "000"& X"000000" & X"2"); \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4888;
              end if;
            when PAUSE_SET4894 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18480\ := eclat_unit;
              \$v4893\ := \$code_lock\;
              if \$v4893\(0) = '1' then
                state_var5922 := Q_WAIT4892;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 10;\$code_write\ <= "000"& X"00000" & X"7f"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4891;
              end if;
            when PAUSE_SET4897 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18479\ := eclat_unit;
              \$v4896\ := \$code_lock\;
              if \$v4896\(0) = '1' then
                state_var5922 := Q_WAIT4895;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 9;\$code_write\ <= "000"& X"000000" & X"0"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4894;
              end if;
            when PAUSE_SET4900 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18478\ := eclat_unit;
              \$v4899\ := \$code_lock\;
              if \$v4899\(0) = '1' then
                state_var5922 := Q_WAIT4898;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 8;\$code_write\ <= "000"& X"000000" & X"1"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4897;
              end if;
            when PAUSE_SET4903 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18477\ := eclat_unit;
              \$v4902\ := \$code_lock\;
              if \$v4902\(0) = '1' then
                state_var5922 := Q_WAIT4901;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 7;\$code_write\ <= "000"& X"00000" & X"28"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4900;
              end if;
            when PAUSE_SET4906 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18476\ := eclat_unit;
              \$v4905\ := \$code_lock\;
              if \$v4905\(0) = '1' then
                state_var5922 := Q_WAIT4904;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 6;\$code_write\ <= "000"& X"00000" & X"64"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4903;
              end if;
            when PAUSE_SET4909 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18475\ := eclat_unit;
              \$v4908\ := \$code_lock\;
              if \$v4908\(0) = '1' then
                state_var5922 := Q_WAIT4907;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 5;\$code_write\ <= "000"& X"000000" & X"4"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4906;
              end if;
            when PAUSE_SET4912 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18474\ := eclat_unit;
              \$v4911\ := \$code_lock\;
              if \$v4911\(0) = '1' then
                state_var5922 := Q_WAIT4910;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 4;\$code_write\ <= "000"& X"000000" & X"2"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4909;
              end if;
            when PAUSE_SET4915 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18473\ := eclat_unit;
              \$v4914\ := \$code_lock\;
              if \$v4914\(0) = '1' then
                state_var5922 := Q_WAIT4913;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 3;\$code_write\ <= "000"& X"00000" & X"86"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4912;
              end if;
            when PAUSE_SET4918 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18472\ := eclat_unit;
              \$v4917\ := \$code_lock\;
              if \$v4917\(0) = '1' then
                state_var5922 := Q_WAIT4916;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 2;\$code_write\ <= "000"& X"000000" & X"0"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4915;
              end if;
            when PAUSE_SET4921 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$18471\ := eclat_unit;
              \$v4920\ := \$code_lock\;
              if \$v4920\(0) = '1' then
                state_var5922 := Q_WAIT4919;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 1;\$code_write\ <= "000"& X"00000" & X"15"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4918;
              end if;
            when PAUSE_SET4924 =>
              \$global_end_write_request\ <= '0';
              release(\$global_end_lock\);
              \$18470\ := eclat_unit;
              \$v4923\ := \$code_lock\;
              if \$v4923\(0) = '1' then
                state_var5922 := Q_WAIT4922;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 0;\$code_write\ <= "000"& X"00000" & X"54"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4921;
              end if;
            when Q_WAIT4576 =>
              \$v4577\ := \$ram_lock\;
              if \$v4577\(0) = '1' then
                state_var5922 := Q_WAIT4576;
              else
                acquire(\$ram_lock\);
                \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                        \$18466_loop666_arg\(16 to 31), \$18466_loop666_arg\(0 to 15))));
                \$ram_write\ <= \$18785\; \$ram_write_request\ <= '1';
                state_var5922 := PAUSE_SET4575;
              end if;
            when Q_WAIT4579 =>
              \$v4580\ := \$ram_lock\;
              if \$v4580\(0) = '1' then
                state_var5922 := Q_WAIT4579;
              else
                acquire(\$ram_lock\);
                \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$18466_loop666_arg\(32 to 47), \$18466_loop666_arg\(0 to 15))));
                state_var5922 := PAUSE_GET4578;
              end if;
            when Q_WAIT4583 =>
              \$v4584\ := \$ram_lock\;
              if \$v4584\(0) = '1' then
                state_var5922 := Q_WAIT4583;
              else
                acquire(\$ram_lock\);
                \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                        \$18467_loop665_arg\(64 to 79), \$18467_loop665_arg\(0 to 15))));
                \$ram_write\ <= \$18766\(0 to 31); \$ram_write_request\ <= '1';
                state_var5922 := PAUSE_SET4582;
              end if;
            when Q_WAIT4586 =>
              \$v4587\ := \$ram_lock\;
              if \$v4587\(0) = '1' then
                state_var5922 := Q_WAIT4586;
              else
                acquire(\$ram_lock\);
                \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                        eclat_resize(\$18765\(0 to 30),16), X"000" & X"1")));
                \$ram_write\ <= eclat_resize(\$18467_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                state_var5922 := PAUSE_SET4585;
              end if;
            when Q_WAIT4589 =>
              \$v4590\ := \$ram_lock\;
              if \$v4590\(0) = '1' then
                state_var5922 := Q_WAIT4589;
              else
                acquire(\$ram_lock\);
                \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18765\(0 to 30),16)));
                \$ram_write\ <= eclat_resize(\$18467_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                state_var5922 := PAUSE_SET4588;
              end if;
            when Q_WAIT4592 =>
              \$v4593\ := \$ram_lock\;
              if \$v4593\(0) = '1' then
                state_var5922 := Q_WAIT4592;
              else
                acquire(\$ram_lock\);
                \$ram_ptr_write\ <= to_integer(unsigned(\$18467_loop665_arg\(16 to 31)));
                \$ram_write\ <= \$18769_hd\; \$ram_write_request\ <= '1';
                state_var5922 := PAUSE_SET4591;
              end if;
            when Q_WAIT4595 =>
              \$v4596\ := \$ram_lock\;
              if \$v4596\(0) = '1' then
                state_var5922 := Q_WAIT4595;
              else
                acquire(\$ram_lock\);
                \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18765\(0 to 30),16)));
                state_var5922 := PAUSE_GET4594;
              end if;
            when Q_WAIT4599 =>
              \$v4600\ := \$ram_lock\;
              if \$v4600\(0) = '1' then
                state_var5922 := Q_WAIT4599;
              else
                acquire(\$ram_lock\);
                \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18765\(0 to 30),16), X"000" & X"1")));
                state_var5922 := PAUSE_GET4598;
              end if;
            when Q_WAIT4603 =>
              \$v4604\ := \$ram_lock\;
              if \$v4604\(0) = '1' then
                state_var5922 := Q_WAIT4603;
              else
                acquire(\$ram_lock\);
                \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$18467_loop665_arg\(64 to 79), \$18467_loop665_arg\(0 to 15))));
                state_var5922 := PAUSE_GET4602;
              end if;
            when Q_WAIT4817 =>
              \$v4818\ := \$ram_lock\;
              if \$v4818\(0) = '1' then
                state_var5922 := Q_WAIT4817;
              else
                acquire(\$ram_lock\);
                \$ram_ptr_write\ <= to_integer(unsigned(\$18512\(64 to 79)));
                \$ram_write\ <= work.Int.lor(work.Int.lsl(eclat_resize(\$18469_make_block579_arg\(80 to 111),31), X"000000" & X"18"), 
                                             work.Int.lsl(eclat_resize(
                                                          eclat_if(work.Int.eq(
                                                                   \$18469_make_block579_arg\(112 to 127), X"000" & X"0") & X"000" & X"1" & \$18469_make_block579_arg\(112 to 127)),31), X"0000000" & X"2")) & eclat_true; \$ram_write_request\ <= '1';
                state_var5922 := PAUSE_SET4816;
              end if;
            when Q_WAIT4820 =>
              \$v4821\ := \$code_lock\;
              if \$v4821\(0) = '1' then
                state_var5922 := Q_WAIT4820;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 34;\$code_write\ <= "000"& X"00000" & X"8f"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4819;
              end if;
            when Q_WAIT4823 =>
              \$v4824\ := \$code_lock\;
              if \$v4824\(0) = '1' then
                state_var5922 := Q_WAIT4823;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 33;\$code_write\ <= "000"& X"000000" & X"1"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4822;
              end if;
            when Q_WAIT4826 =>
              \$v4827\ := \$code_lock\;
              if \$v4827\(0) = '1' then
                state_var5922 := Q_WAIT4826;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 32;\$code_write\ <= "000"& X"00000" & X"13"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4825;
              end if;
            when Q_WAIT4829 =>
              \$v4830\ := \$code_lock\;
              if \$v4830\(0) = '1' then
                state_var5922 := Q_WAIT4829;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 31;\$code_write\ <= "000"& X"000000" & X"0"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4828;
              end if;
            when Q_WAIT4832 =>
              \$v4833\ := \$code_lock\;
              if \$v4833\(0) = '1' then
                state_var5922 := Q_WAIT4832;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 30;\$code_write\ <= "000"& X"00000" & X"5d"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4831;
              end if;
            when Q_WAIT4835 =>
              \$v4836\ := \$code_lock\;
              if \$v4836\(0) = '1' then
                state_var5922 := Q_WAIT4835;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 29;\$code_write\ <= "000"& X"00000" & X"21"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4834;
              end if;
            when Q_WAIT4838 =>
              \$v4839\ := \$code_lock\;
              if \$v4839\(0) = '1' then
                state_var5922 := Q_WAIT4838;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 28;\$code_write\ <= "000"& X"000000" & X"b"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4837;
              end if;
            when Q_WAIT4841 =>
              \$v4842\ := \$code_lock\;
              if \$v4842\(0) = '1' then
                state_var5922 := Q_WAIT4841;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 27;\$code_write\ <= "000"& X"000000" & X"b"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4840;
              end if;
            when Q_WAIT4844 =>
              \$v4845\ := \$code_lock\;
              if \$v4845\(0) = '1' then
                state_var5922 := Q_WAIT4844;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 26;\$code_write\ <= "000"& X"00000" & X"67"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4843;
              end if;
            when Q_WAIT4847 =>
              \$v4848\ := \$code_lock\;
              if \$v4848\(0) = '1' then
                state_var5922 := Q_WAIT4847;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 25;\$code_write\ <= work.Int.neg(
                                                         "000"& X"00000" & X"17"); \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4846;
              end if;
            when Q_WAIT4850 =>
              \$v4851\ := \$code_lock\;
              if \$v4851\(0) = '1' then
                state_var5922 := Q_WAIT4850;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 24;\$code_write\ <= "000"& X"000000" & X"0"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4849;
              end if;
            when Q_WAIT4853 =>
              \$v4854\ := \$code_lock\;
              if \$v4854\(0) = '1' then
                state_var5922 := Q_WAIT4853;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 23;\$code_write\ <= "000"& X"000000" & X"1"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4852;
              end if;
            when Q_WAIT4856 =>
              \$v4857\ := \$code_lock\;
              if \$v4857\(0) = '1' then
                state_var5922 := Q_WAIT4856;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 22;\$code_write\ <= "000"& X"00000" & X"2c"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4855;
              end if;
            when Q_WAIT4859 =>
              \$v4860\ := \$code_lock\;
              if \$v4860\(0) = '1' then
                state_var5922 := Q_WAIT4859;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 21;\$code_write\ <= "000"& X"000000" & X"1"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4858;
              end if;
            when Q_WAIT4862 =>
              \$v4863\ := \$code_lock\;
              if \$v4863\(0) = '1' then
                state_var5922 := Q_WAIT4862;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 20;\$code_write\ <= "000"& X"00000" & X"28"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4861;
              end if;
            when Q_WAIT4865 =>
              \$v4866\ := \$code_lock\;
              if \$v4866\(0) = '1' then
                state_var5922 := Q_WAIT4865;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 19;\$code_write\ <= "000"& X"00000" & X"6e"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4864;
              end if;
            when Q_WAIT4868 =>
              \$v4869\ := \$code_lock\;
              if \$v4869\(0) = '1' then
                state_var5922 := Q_WAIT4868;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 18;\$code_write\ <= "000"& X"00000" & X"21"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4867;
              end if;
            when Q_WAIT4871 =>
              \$v4872\ := \$code_lock\;
              if \$v4872\(0) = '1' then
                state_var5922 := Q_WAIT4871;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 17;\$code_write\ <= "000"& X"00000" & X"32"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4870;
              end if;
            when Q_WAIT4874 =>
              \$v4875\ := \$code_lock\;
              if \$v4875\(0) = '1' then
                state_var5922 := Q_WAIT4874;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 16;\$code_write\ <= work.Int.neg(
                                                         "000"& X"000000" & X"1"); \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4873;
              end if;
            when Q_WAIT4877 =>
              \$v4878\ := \$code_lock\;
              if \$v4878\(0) = '1' then
                state_var5922 := Q_WAIT4877;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 15;\$code_write\ <= "000"& X"00000" & X"7f"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4876;
              end if;
            when Q_WAIT4880 =>
              \$v4881\ := \$code_lock\;
              if \$v4881\(0) = '1' then
                state_var5922 := Q_WAIT4880;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 14;\$code_write\ <= "000"& X"000000" & X"b"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4879;
              end if;
            when Q_WAIT4883 =>
              \$v4884\ := \$code_lock\;
              if \$v4884\(0) = '1' then
                state_var5922 := Q_WAIT4883;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 13;\$code_write\ <= "000"& X"00000" & X"21"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4882;
              end if;
            when Q_WAIT4886 =>
              \$v4887\ := \$code_lock\;
              if \$v4887\(0) = '1' then
                state_var5922 := Q_WAIT4886;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 12;\$code_write\ <= "000"& X"00000" & X"32"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4885;
              end if;
            when Q_WAIT4889 =>
              \$v4890\ := \$code_lock\;
              if \$v4890\(0) = '1' then
                state_var5922 := Q_WAIT4889;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 11;\$code_write\ <= work.Int.neg(
                                                         "000"& X"000000" & X"2"); \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4888;
              end if;
            when Q_WAIT4892 =>
              \$v4893\ := \$code_lock\;
              if \$v4893\(0) = '1' then
                state_var5922 := Q_WAIT4892;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 10;\$code_write\ <= "000"& X"00000" & X"7f"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4891;
              end if;
            when Q_WAIT4895 =>
              \$v4896\ := \$code_lock\;
              if \$v4896\(0) = '1' then
                state_var5922 := Q_WAIT4895;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 9;\$code_write\ <= "000"& X"000000" & X"0"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4894;
              end if;
            when Q_WAIT4898 =>
              \$v4899\ := \$code_lock\;
              if \$v4899\(0) = '1' then
                state_var5922 := Q_WAIT4898;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 8;\$code_write\ <= "000"& X"000000" & X"1"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4897;
              end if;
            when Q_WAIT4901 =>
              \$v4902\ := \$code_lock\;
              if \$v4902\(0) = '1' then
                state_var5922 := Q_WAIT4901;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 7;\$code_write\ <= "000"& X"00000" & X"28"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4900;
              end if;
            when Q_WAIT4904 =>
              \$v4905\ := \$code_lock\;
              if \$v4905\(0) = '1' then
                state_var5922 := Q_WAIT4904;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 6;\$code_write\ <= "000"& X"00000" & X"64"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4903;
              end if;
            when Q_WAIT4907 =>
              \$v4908\ := \$code_lock\;
              if \$v4908\(0) = '1' then
                state_var5922 := Q_WAIT4907;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 5;\$code_write\ <= "000"& X"000000" & X"4"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4906;
              end if;
            when Q_WAIT4910 =>
              \$v4911\ := \$code_lock\;
              if \$v4911\(0) = '1' then
                state_var5922 := Q_WAIT4910;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 4;\$code_write\ <= "000"& X"000000" & X"2"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4909;
              end if;
            when Q_WAIT4913 =>
              \$v4914\ := \$code_lock\;
              if \$v4914\(0) = '1' then
                state_var5922 := Q_WAIT4913;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 3;\$code_write\ <= "000"& X"00000" & X"86"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4912;
              end if;
            when Q_WAIT4916 =>
              \$v4917\ := \$code_lock\;
              if \$v4917\(0) = '1' then
                state_var5922 := Q_WAIT4916;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 2;\$code_write\ <= "000"& X"000000" & X"0"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4915;
              end if;
            when Q_WAIT4919 =>
              \$v4920\ := \$code_lock\;
              if \$v4920\(0) = '1' then
                state_var5922 := Q_WAIT4919;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 1;\$code_write\ <= "000"& X"00000" & X"15"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4918;
              end if;
            when Q_WAIT4922 =>
              \$v4923\ := \$code_lock\;
              if \$v4923\(0) = '1' then
                state_var5922 := Q_WAIT4922;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 0;\$code_write\ <= "000"& X"00000" & X"54"; \$code_write_request\ <= '1';
                state_var5922 := PAUSE_SET4921;
              end if;
            when Q_WAIT4925 =>
              \$v4926\ := \$global_end_lock\;
              if \$v4926\(0) = '1' then
                state_var5922 := Q_WAIT4925;
              else
                acquire(\$global_end_lock\);
                \$global_end_ptr_write\ <= 0;\$global_end_write\ <= work.Int.add(
                                                                    X"3e80", X"000" & X"c"); \$global_end_write_request\ <= '1';
                state_var5922 := PAUSE_SET4924;
              end if;
            when IDLE4574 =>
              rdy4573 := eclat_false;
              \$v4926\ := \$global_end_lock\;
              if \$v4926\(0) = '1' then
                state_var5922 := Q_WAIT4925;
              else
                acquire(\$global_end_lock\);
                \$global_end_ptr_write\ <= 0;\$global_end_write\ <= work.Int.add(
                                                                    X"3e80", X"000" & X"c"); \$global_end_write_request\ <= '1';
                state_var5922 := PAUSE_SET4924;
              end if;
            end case;
            
            if rdy4573(0) = '1' then
              
            else
              result4572 := eclat_unit;
            end if;
            \$18463\ := result4572 & rdy4573;
            if \$v4332\(0) = '1' then
              
            else
              \$v4332\ := eclat_true;
              \$18465\ := eclat_false;
            end if;
            \$18465\ := work.Bool.land(eclat_if(\$18465\ & eclat_true & ""&\$18463\(1)), 
                                       work.Bool.lnot(eclat_false));
            \$18464_rdy\ := \$18465\;
            \$18462\ := eclat_false & eclat_true & \$18464_rdy\ & ""&\$18462\(3);
          else
            if \$v4333\(0) = '1' then
              
            else
              \$v4333\ := eclat_true;
              \$18788\ := X"000" & X"0" & "000"& X"000000" & X"1" & eclat_true & X"0" & X"3e8" & "000"& X"000000" & X"1" & eclat_true & "00000000" & X"000" & X"0" & eclat_false & eclat_false & eclat_true;
            end if;
            \$v5917\ := work.Bool.lnot(""&\$18462\(2));
            if \$v5917\(0) = '1' then
              \$18788\ := \$18788\(0 to 121) & eclat_true;
            else
              case state_var5920 is
              when \$18790_LOOP666\ =>
                \$v4937\ := work.Int.ge(\$18790_loop666_arg\(0 to 15), 
                                        work.Int.add(\$18790_loop666_arg\(48 to 63), X"000" & X"1"));
                if \$v4937\(0) = '1' then
                  \$18790_loop666_result\ := eclat_unit;
                  \$19756\ := \$18790_loop666_result\;
                  \$v4946\ := \$ram_lock\;
                  if \$v4946\(0) = '1' then
                    state_var5920 := Q_WAIT4945;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$19741\(0 to 30),16)));
                    \$ram_write\ <= eclat_resize(\$18791_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET4944;
                  end if;
                else
                  \$v4936\ := \$ram_lock\;
                  if \$v4936\(0) = '1' then
                    state_var5920 := Q_WAIT4935;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$18790_loop666_arg\(32 to 47), \$18790_loop666_arg\(0 to 15))));
                    state_var5920 := PAUSE_GET4934;
                  end if;
                end if;
              when \$18791_LOOP665\ =>
                \$v4961\ := work.Int.ge(\$18791_loop665_arg\(0 to 15), 
                                        work.Int.add(\$18791_loop665_arg\(80 to 95), X"000" & X"1"));
                if \$v4961\(0) = '1' then
                  \$18791_loop665_result\ := \$18791_loop665_arg\(16 to 31);
                  state_var5920 := \$18791_LOOP665\;
                else
                  \$v4960\ := \$ram_lock\;
                  if \$v4960\(0) = '1' then
                    state_var5920 := Q_WAIT4959;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$18791_loop665_arg\(64 to 79), \$18791_loop665_arg\(0 to 15))));
                    state_var5920 := PAUSE_GET4958;
                  end if;
                end if;
              when \$18792_WAIT662\ =>
                if \$v4335\(0) = '1' then
                  
                else
                  \$v4335\ := eclat_true;
                  \$19493\ := \$18792_wait662_arg\(1 to 32) & \$18792_wait662_arg\(33 to 64) & X"0" & X"fa0" & X"0" & X"fa0" & X"0" & X"fa0" & 
                  work.Int.add(X"0" & X"fa0", X"1770") & eclat_false;
                end if;
                case state_var5921 is
                when \$19494_LOOP666\ =>
                  \$v4972\ := work.Int.ge(\$19494_loop666_arg\(0 to 15), 
                                          work.Int.add(\$19494_loop666_arg\(48 to 63), X"000" & X"1"));
                  if \$v4972\(0) = '1' then
                    \$19494_loop666_result\ := eclat_unit;
                    \$19732\ := \$19494_loop666_result\;
                    \$v4981\ := \$ram_lock\;
                    if \$v4981\(0) = '1' then
                      state_var5921 := Q_WAIT4980;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$19717\(0 to 30),16)));
                      \$ram_write\ <= eclat_resize(\$19495_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                      state_var5921 := PAUSE_SET4979;
                    end if;
                  else
                    \$v4971\ := \$ram_lock\;
                    if \$v4971\(0) = '1' then
                      state_var5921 := Q_WAIT4970;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                        \$19494_loop666_arg\(32 to 47), \$19494_loop666_arg\(0 to 15))));
                      state_var5921 := PAUSE_GET4969;
                    end if;
                  end if;
                when \$19495_LOOP665\ =>
                  \$v4996\ := work.Int.ge(\$19495_loop665_arg\(0 to 15), 
                                          work.Int.add(\$19495_loop665_arg\(80 to 95), X"000" & X"1"));
                  if \$v4996\(0) = '1' then
                    \$19495_loop665_result\ := \$19495_loop665_arg\(16 to 31);
                    \$19714_next\ := \$19495_loop665_result\;
                    \$19496_aux664_arg\ := work.Int.add(\$19496_aux664_arg\(0 to 15), 
                                                        work.Int.add(
                                                        eclat_resize(
                                                        work.Int.lsr(
                                                        eclat_resize(eclat_resize(\$19713\(0 to 30),16),31), X"0000000" & X"2"),16), X"000" & X"1")) & \$19714_next\ & \$19496_aux664_arg\(32 to 47) & \$19496_aux664_arg\(48 to 63);
                    state_var5921 := \$19496_AUX664\;
                  else
                    \$v4995\ := \$ram_lock\;
                    if \$v4995\(0) = '1' then
                      state_var5921 := Q_WAIT4994;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                        \$19495_loop665_arg\(64 to 79), \$19495_loop665_arg\(0 to 15))));
                      state_var5921 := PAUSE_GET4993;
                    end if;
                  end if;
                when \$19496_AUX664\ =>
                  \$19708\ := work.Print.print_string(clk,of_string("     scan="));
                  \$19709\ := work.Int.print(clk,\$19496_aux664_arg\(0 to 15));
                  \$19710\ := work.Print.print_string(clk,of_string(" | next="));
                  \$19711\ := work.Int.print(clk,\$19496_aux664_arg\(16 to 31));
                  \$19712\ := work.Print.print_newline(clk,eclat_unit);
                  \$v5000\ := work.Int.ge(\$19496_aux664_arg\(0 to 15), \$19496_aux664_arg\(16 to 31));
                  if \$v5000\(0) = '1' then
                    \$19496_aux664_result\ := \$19496_aux664_arg\(16 to 31);
                    state_var5921 := \$19496_AUX664\;
                  else
                    \$v4999\ := \$ram_lock\;
                    if \$v4999\(0) = '1' then
                      state_var5921 := Q_WAIT4998;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(\$19496_aux664_arg\(0 to 15)));
                      state_var5921 := PAUSE_GET4997;
                    end if;
                  end if;
                when \$19497_LOOP666\ =>
                  \$v5007\ := work.Int.ge(\$19497_loop666_arg\(0 to 15), 
                                          work.Int.add(\$19497_loop666_arg\(48 to 63), X"000" & X"1"));
                  if \$v5007\(0) = '1' then
                    \$19497_loop666_result\ := eclat_unit;
                    case \$19497_loop666_id\ is
                    when "000000100011" =>
                      \$19699\ := \$19497_loop666_result\;
                      \$v5016\ := \$ram_lock\;
                      if \$v5016\(0) = '1' then
                        state_var5921 := Q_WAIT5015;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$19684\(0 to 30),16)));
                        \$ram_write\ <= eclat_resize(\$19498_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                        state_var5921 := PAUSE_SET5014;
                      end if;
                    when "000000101001" =>
                      \$19571\ := \$19497_loop666_result\;
                      \$v5045\ := \$ram_lock\;
                      if \$v5045\(0) = '1' then
                        state_var5921 := Q_WAIT5044;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$19553\(0 to 30),16)));
                        \$ram_write\ <= eclat_resize(\$19547_copy_root_in_ram6634352_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                        state_var5921 := PAUSE_SET5043;
                      end if;
                    when "000000101011" =>
                      \$19586\ := \$19497_loop666_result\;
                      \$v5069\ := \$ram_lock\;
                      if \$v5069\(0) = '1' then
                        state_var5921 := Q_WAIT5068;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$19541\(0 to 30),16)));
                        \$ram_write\ <= eclat_resize(\$19535_copy_root_in_ram6634354_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                        state_var5921 := PAUSE_SET5067;
                      end if;
                    when "000000101101" =>
                      \$19625\ := \$19497_loop666_result\;
                      \$v5096\ := \$ram_lock\;
                      if \$v5096\(0) = '1' then
                        state_var5921 := Q_WAIT5095;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$19607\(0 to 30),16)));
                        \$ram_write\ <= eclat_resize(\$19601_copy_root_in_ram6634352_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                        state_var5921 := PAUSE_SET5094;
                      end if;
                    when "000000101111" =>
                      \$19640\ := \$19497_loop666_result\;
                      \$v5120\ := \$ram_lock\;
                      if \$v5120\(0) = '1' then
                        state_var5921 := Q_WAIT5119;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$19595\(0 to 30),16)));
                        \$ram_write\ <= eclat_resize(\$19589_copy_root_in_ram6634353_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                        state_var5921 := PAUSE_SET5118;
                      end if;
                    when "000000110001" =>
                      \$19655\ := \$19497_loop666_result\;
                      \$v5141\ := \$ram_lock\;
                      if \$v5141\(0) = '1' then
                        state_var5921 := Q_WAIT5140;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18792_wait662_arg\(33 to 63),16)));
                        \$ram_write\ <= eclat_resize(\$19505\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                        state_var5921 := PAUSE_SET5139;
                      end if;
                    when "000000110010" =>
                      \$19670\ := \$19497_loop666_result\;
                      \$v5158\ := \$ram_lock\;
                      if \$v5158\(0) = '1' then
                        state_var5921 := Q_WAIT5157;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18792_wait662_arg\(1 to 31),16)));
                        \$ram_write\ <= eclat_resize(\$19493\(112 to 127),31) & eclat_false; \$ram_write_request\ <= '1';
                        state_var5921 := PAUSE_SET5156;
                      end if;
                    when others =>
                      
                    end case;
                  else
                    \$v5006\ := \$ram_lock\;
                    if \$v5006\(0) = '1' then
                      state_var5921 := Q_WAIT5005;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                        \$19497_loop666_arg\(32 to 47), \$19497_loop666_arg\(0 to 15))));
                      state_var5921 := PAUSE_GET5004;
                    end if;
                  end if;
                when \$19498_LOOP665\ =>
                  \$v5031\ := work.Int.ge(\$19498_loop665_arg\(0 to 15), 
                                          work.Int.add(\$19498_loop665_arg\(80 to 95), X"000" & X"1"));
                  if \$v5031\(0) = '1' then
                    \$19498_loop665_result\ := \$19498_loop665_arg\(16 to 31);
                    \$19681_next\ := \$19498_loop665_result\;
                    \$19499_aux664_arg\ := work.Int.add(\$19499_aux664_arg\(0 to 15), 
                                                        work.Int.add(
                                                        eclat_resize(
                                                        work.Int.lsr(
                                                        eclat_resize(eclat_resize(\$19680\(0 to 30),16),31), X"0000000" & X"2"),16), X"000" & X"1")) & \$19681_next\ & \$19499_aux664_arg\(32 to 47) & \$19499_aux664_arg\(48 to 63);
                    state_var5921 := \$19499_AUX664\;
                  else
                    \$v5030\ := \$ram_lock\;
                    if \$v5030\(0) = '1' then
                      state_var5921 := Q_WAIT5029;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                        \$19498_loop665_arg\(64 to 79), \$19498_loop665_arg\(0 to 15))));
                      state_var5921 := PAUSE_GET5028;
                    end if;
                  end if;
                when \$19499_AUX664\ =>
                  \$19675\ := work.Print.print_string(clk,of_string("     scan="));
                  \$19676\ := work.Int.print(clk,\$19499_aux664_arg\(0 to 15));
                  \$19677\ := work.Print.print_string(clk,of_string(" | next="));
                  \$19678\ := work.Int.print(clk,\$19499_aux664_arg\(16 to 31));
                  \$19679\ := work.Print.print_newline(clk,eclat_unit);
                  \$v5035\ := work.Int.ge(\$19499_aux664_arg\(0 to 15), \$19499_aux664_arg\(16 to 31));
                  if \$v5035\(0) = '1' then
                    \$19499_aux664_result\ := \$19499_aux664_arg\(16 to 31);
                    \$19518_next\ := \$19499_aux664_result\;
                    \$19519\ := work.Print.print_string(clk,of_string("memory copied in to_space : "));
                    \$19520\ := work.Int.print(clk,work.Int.sub(\$19518_next\, \$19493\(112 to 127)));
                    \$19521\ := work.Print.print_string(clk,of_string(" words"));
                    \$19522\ := work.Print.print_newline(clk,eclat_unit);
                    \$v5036\ := work.Int.gt(work.Int.sub(\$19518_next\, \$19493\(112 to 127)), X"1770");
                    if \$v5036\(0) = '1' then
                      \$19523\ := work.Print.print_string(clk,of_string("fatal error: "));
                      \$19524\ := work.Print.print_string(clk,of_string("Out of memory"));
                      \$19525\ := work.Print.print_newline(clk,eclat_unit);
                      \$19526_forever6704355_id\ := "000000100111";
                      \$19526_forever6704355_arg\ := eclat_unit;
                      state_var5921 := \$19526_FOREVER6704355\;
                    else
                      \$19508\ := \$19505\(0 to 31) & \$19506\(0 to 31) & \$19518_next\;
                      \$19509\ := work.Print.print_newline(clk,eclat_unit);
                      \$19510\ := work.Print.print_newline(clk,eclat_unit);
                      \$19511\ := work.Print.print_string(clk,of_string("[================= GC END ======================]"));
                      \$19512\ := work.Print.print_newline(clk,eclat_unit);
                      \$19513\ := work.Print.print_newline(clk,eclat_unit);
                      result4963 := \$19508\(0 to 31) & \$19508\(32 to 63) & \$19508\(64 to 79) & 
                      work.Int.add(\$19508\(64 to 79), \$18792_wait662_arg\(81 to 96)) & \$19493\(112 to 127) & \$19493\(96 to 111);
                      rdy4964 := eclat_true;
                      state_var5921 := IDLE4965;
                    end if;
                  else
                    \$v5034\ := \$ram_lock\;
                    if \$v5034\(0) = '1' then
                      state_var5921 := Q_WAIT5033;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(\$19499_aux664_arg\(0 to 15)));
                      state_var5921 := PAUSE_GET5032;
                    end if;
                  end if;
                when \$19526_FOREVER6704355\ =>
                  \$19529_forever6704351_id\ := "000000100110";
                  \$19529_forever6704351_arg\ := eclat_unit;
                  state_var5921 := \$19529_FOREVER6704351\;
                when \$19529_FOREVER6704351\ =>
                  \$19532_forever6704350_id\ := "000000100101";
                  \$19532_forever6704350_arg\ := eclat_unit;
                  state_var5921 := \$19532_FOREVER6704350\;
                when \$19532_FOREVER6704350\ =>
                  \$19532_forever6704350_arg\ := eclat_unit;
                  state_var5921 := \$19532_FOREVER6704350\;
                when \$19535_COPY_ROOT_IN_RAM6634354\ =>
                  \$v5084\ := work.Int.ge(\$19535_copy_root_in_ram6634354_arg\(0 to 15), \$19535_copy_root_in_ram6634354_arg\(16 to 31));
                  if \$v5084\(0) = '1' then
                    \$19535_copy_root_in_ram6634354_result\ := \$19535_copy_root_in_ram6634354_arg\(32 to 47);
                    \$19515_next\ := \$19535_copy_root_in_ram6634354_result\;
                    \$19516\ := work.Print.print_string(clk,of_string("======================================="));
                    \$19517\ := work.Print.print_newline(clk,eclat_unit);
                    \$19499_aux664_id\ := "000000101000";
                    \$19499_aux664_arg\ := \$19493\(112 to 127) & \$19515_next\ & \$19493\(96 to 111) & \$19493\(112 to 127);
                    state_var5921 := \$19499_AUX664\;
                  else
                    \$19538\ := work.Print.print_string(clk,of_string("racine:"));
                    \$19539\ := work.Int.print(clk,\$19535_copy_root_in_ram6634354_arg\(0 to 15));
                    \$19540\ := work.Print.print_newline(clk,eclat_unit);
                    \$v5083\ := \$ram_lock\;
                    if \$v5083\(0) = '1' then
                      state_var5921 := Q_WAIT5082;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(\$19535_copy_root_in_ram6634354_arg\(0 to 15)));
                      state_var5921 := PAUSE_GET5081;
                    end if;
                  end if;
                when \$19547_COPY_ROOT_IN_RAM6634352\ =>
                  \$v5060\ := work.Int.ge(\$19547_copy_root_in_ram6634352_arg\(0 to 15), \$19547_copy_root_in_ram6634352_arg\(16 to 31));
                  if \$v5060\(0) = '1' then
                    \$19547_copy_root_in_ram6634352_result\ := \$19547_copy_root_in_ram6634352_arg\(32 to 47);
                    \$19535_copy_root_in_ram6634354_result\ := \$19547_copy_root_in_ram6634352_result\;
                    \$19515_next\ := \$19535_copy_root_in_ram6634354_result\;
                    \$19516\ := work.Print.print_string(clk,of_string("======================================="));
                    \$19517\ := work.Print.print_newline(clk,eclat_unit);
                    \$19499_aux664_id\ := "000000101000";
                    \$19499_aux664_arg\ := \$19493\(112 to 127) & \$19515_next\ & \$19493\(96 to 111) & \$19493\(112 to 127);
                    state_var5921 := \$19499_AUX664\;
                  else
                    \$19550\ := work.Print.print_string(clk,of_string("racine:"));
                    \$19551\ := work.Int.print(clk,\$19547_copy_root_in_ram6634352_arg\(0 to 15));
                    \$19552\ := work.Print.print_newline(clk,eclat_unit);
                    \$v5059\ := \$ram_lock\;
                    if \$v5059\(0) = '1' then
                      state_var5921 := Q_WAIT5058;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(\$19547_copy_root_in_ram6634352_arg\(0 to 15)));
                      state_var5921 := PAUSE_GET5057;
                    end if;
                  end if;
                when \$19589_COPY_ROOT_IN_RAM6634353\ =>
                  \$v5135\ := work.Int.ge(\$19589_copy_root_in_ram6634353_arg\(0 to 15), \$19589_copy_root_in_ram6634353_arg\(16 to 31));
                  if \$v5135\(0) = '1' then
                    \$19589_copy_root_in_ram6634353_result\ := \$19589_copy_root_in_ram6634353_arg\(32 to 47);
                    \$19507_next\ := \$19589_copy_root_in_ram6634353_result\;
                    \$v5087\ := \$global_end_lock\;
                    if \$v5087\(0) = '1' then
                      state_var5921 := Q_WAIT5086;
                    else
                      acquire(\$global_end_lock\);
                      \$global_end_ptr\ <= 0;
                      state_var5921 := PAUSE_GET5085;
                    end if;
                  else
                    \$19592\ := work.Print.print_string(clk,of_string("racine:"));
                    \$19593\ := work.Int.print(clk,\$19589_copy_root_in_ram6634353_arg\(0 to 15));
                    \$19594\ := work.Print.print_newline(clk,eclat_unit);
                    \$v5134\ := \$ram_lock\;
                    if \$v5134\(0) = '1' then
                      state_var5921 := Q_WAIT5133;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(\$19589_copy_root_in_ram6634353_arg\(0 to 15)));
                      state_var5921 := PAUSE_GET5132;
                    end if;
                  end if;
                when \$19601_COPY_ROOT_IN_RAM6634352\ =>
                  \$v5111\ := work.Int.ge(\$19601_copy_root_in_ram6634352_arg\(0 to 15), \$19601_copy_root_in_ram6634352_arg\(16 to 31));
                  if \$v5111\(0) = '1' then
                    \$19601_copy_root_in_ram6634352_result\ := \$19601_copy_root_in_ram6634352_arg\(32 to 47);
                    \$19589_copy_root_in_ram6634353_result\ := \$19601_copy_root_in_ram6634352_result\;
                    \$19507_next\ := \$19589_copy_root_in_ram6634353_result\;
                    \$v5087\ := \$global_end_lock\;
                    if \$v5087\(0) = '1' then
                      state_var5921 := Q_WAIT5086;
                    else
                      acquire(\$global_end_lock\);
                      \$global_end_ptr\ <= 0;
                      state_var5921 := PAUSE_GET5085;
                    end if;
                  else
                    \$19604\ := work.Print.print_string(clk,of_string("racine:"));
                    \$19605\ := work.Int.print(clk,\$19601_copy_root_in_ram6634352_arg\(0 to 15));
                    \$19606\ := work.Print.print_newline(clk,eclat_unit);
                    \$v5110\ := \$ram_lock\;
                    if \$v5110\(0) = '1' then
                      state_var5921 := Q_WAIT5109;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(\$19601_copy_root_in_ram6634352_arg\(0 to 15)));
                      state_var5921 := PAUSE_GET5108;
                    end if;
                  end if;
                when PAUSE_GET4969 =>
                  \$19737\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v4968\ := \$ram_lock\;
                  if \$v4968\(0) = '1' then
                    state_var5921 := Q_WAIT4967;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            \$19494_loop666_arg\(16 to 31), \$19494_loop666_arg\(0 to 15))));
                    \$ram_write\ <= \$19737\; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET4966;
                  end if;
                when PAUSE_GET4985 =>
                  \$19721_hd\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$19722\ := work.Print.print_string(clk,of_string("bloc "));
                  \$19723\ := work.Int.print(clk,eclat_resize(\$19717\(0 to 30),16));
                  \$19724\ := work.Print.print_string(clk,of_string(" of size "));
                  \$19725\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                              work.Int.lsr(
                                                              \$19721_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$19726\ := work.Print.print_string(clk,of_string(" from "));
                  \$19727\ := work.Int.print(clk,eclat_resize(\$19717\(0 to 30),16));
                  \$19728\ := work.Print.print_string(clk,of_string(" to "));
                  \$19729\ := work.Int.print(clk,\$19495_loop665_arg\(16 to 31));
                  \$19730\ := work.Print.print_newline(clk,eclat_unit);
                  \$v4984\ := \$ram_lock\;
                  if \$v4984\(0) = '1' then
                    state_var5921 := Q_WAIT4983;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19495_loop665_arg\(16 to 31)));
                    \$ram_write\ <= \$19721_hd\; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET4982;
                  end if;
                when PAUSE_GET4989 =>
                  \$19720_w\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v4988\ := eclat_if(work.Bool.lnot(""&\$19720_w\(31)) & 
                              eclat_if(work.Int.le(\$19495_loop665_arg\(48 to 63), eclat_resize(\$19720_w\(0 to 30),16)) & 
                              work.Int.lt(eclat_resize(\$19720_w\(0 to 30),16), 
                                          work.Int.add(\$19495_loop665_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false);
                  if \$v4988\(0) = '1' then
                    \$19718\ := \$19720_w\ & \$19495_loop665_arg\(16 to 31);
                    \$v4975\ := \$ram_lock\;
                    if \$v4975\(0) = '1' then
                      state_var5921 := Q_WAIT4974;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                              \$19495_loop665_arg\(64 to 79), \$19495_loop665_arg\(0 to 15))));
                      \$ram_write\ <= \$19718\(0 to 31); \$ram_write_request\ <= '1';
                      state_var5921 := PAUSE_SET4973;
                    end if;
                  else
                    \$v4987\ := \$ram_lock\;
                    if \$v4987\(0) = '1' then
                      state_var5921 := Q_WAIT4986;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$19717\(0 to 30),16)));
                      state_var5921 := PAUSE_GET4985;
                    end if;
                  end if;
                when PAUSE_GET4993 =>
                  \$19717\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v4992\ := work.Bool.lnot(eclat_if(work.Bool.lnot(
                                                      ""&\$19717\(31)) & 
                                             eclat_if(work.Int.le(\$19495_loop665_arg\(32 to 47), eclat_resize(\$19717\(0 to 30),16)) & 
                                             work.Int.lt(eclat_resize(\$19717\(0 to 30),16), 
                                                         work.Int.add(
                                                         \$19495_loop665_arg\(32 to 47), X"1770")) & eclat_false) & eclat_false));
                  if \$v4992\(0) = '1' then
                    \$19718\ := \$19717\ & \$19495_loop665_arg\(16 to 31);
                    \$v4975\ := \$ram_lock\;
                    if \$v4975\(0) = '1' then
                      state_var5921 := Q_WAIT4974;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                              \$19495_loop665_arg\(64 to 79), \$19495_loop665_arg\(0 to 15))));
                      \$ram_write\ <= \$19718\(0 to 31); \$ram_write_request\ <= '1';
                      state_var5921 := PAUSE_SET4973;
                    end if;
                  else
                    \$v4991\ := \$ram_lock\;
                    if \$v4991\(0) = '1' then
                      state_var5921 := Q_WAIT4990;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                        eclat_resize(\$19717\(0 to 30),16), X"000" & X"1")));
                      state_var5921 := PAUSE_GET4989;
                    end if;
                  end if;
                when PAUSE_GET4997 =>
                  \$19713\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$19495_loop665_id\ := "000000100010";
                  \$19495_loop665_arg\ := X"000" & X"1" & \$19496_aux664_arg\(16 to 31) & \$19496_aux664_arg\(32 to 47) & \$19496_aux664_arg\(48 to 63) & \$19496_aux664_arg\(0 to 15) & eclat_resize(
                  work.Int.lsr(eclat_resize(eclat_resize(\$19713\(0 to 30),16),31), X"0000000" & X"2"),16);
                  state_var5921 := \$19495_LOOP665\;
                when PAUSE_GET5004 =>
                  \$19704\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v5003\ := \$ram_lock\;
                  if \$v5003\(0) = '1' then
                    state_var5921 := Q_WAIT5002;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            \$19497_loop666_arg\(16 to 31), \$19497_loop666_arg\(0 to 15))));
                    \$ram_write\ <= \$19704\; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5001;
                  end if;
                when PAUSE_GET5020 =>
                  \$19688_hd\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$19689\ := work.Print.print_string(clk,of_string("bloc "));
                  \$19690\ := work.Int.print(clk,eclat_resize(\$19684\(0 to 30),16));
                  \$19691\ := work.Print.print_string(clk,of_string(" of size "));
                  \$19692\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                              work.Int.lsr(
                                                              \$19688_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$19693\ := work.Print.print_string(clk,of_string(" from "));
                  \$19694\ := work.Int.print(clk,eclat_resize(\$19684\(0 to 30),16));
                  \$19695\ := work.Print.print_string(clk,of_string(" to "));
                  \$19696\ := work.Int.print(clk,\$19498_loop665_arg\(16 to 31));
                  \$19697\ := work.Print.print_newline(clk,eclat_unit);
                  \$v5019\ := \$ram_lock\;
                  if \$v5019\(0) = '1' then
                    state_var5921 := Q_WAIT5018;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19498_loop665_arg\(16 to 31)));
                    \$ram_write\ <= \$19688_hd\; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5017;
                  end if;
                when PAUSE_GET5024 =>
                  \$19687_w\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v5023\ := eclat_if(work.Bool.lnot(""&\$19687_w\(31)) & 
                              eclat_if(work.Int.le(\$19498_loop665_arg\(48 to 63), eclat_resize(\$19687_w\(0 to 30),16)) & 
                              work.Int.lt(eclat_resize(\$19687_w\(0 to 30),16), 
                                          work.Int.add(\$19498_loop665_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false);
                  if \$v5023\(0) = '1' then
                    \$19685\ := \$19687_w\ & \$19498_loop665_arg\(16 to 31);
                    \$v5010\ := \$ram_lock\;
                    if \$v5010\(0) = '1' then
                      state_var5921 := Q_WAIT5009;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                              \$19498_loop665_arg\(64 to 79), \$19498_loop665_arg\(0 to 15))));
                      \$ram_write\ <= \$19685\(0 to 31); \$ram_write_request\ <= '1';
                      state_var5921 := PAUSE_SET5008;
                    end if;
                  else
                    \$v5022\ := \$ram_lock\;
                    if \$v5022\(0) = '1' then
                      state_var5921 := Q_WAIT5021;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$19684\(0 to 30),16)));
                      state_var5921 := PAUSE_GET5020;
                    end if;
                  end if;
                when PAUSE_GET5028 =>
                  \$19684\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v5027\ := work.Bool.lnot(eclat_if(work.Bool.lnot(
                                                      ""&\$19684\(31)) & 
                                             eclat_if(work.Int.le(\$19498_loop665_arg\(32 to 47), eclat_resize(\$19684\(0 to 30),16)) & 
                                             work.Int.lt(eclat_resize(\$19684\(0 to 30),16), 
                                                         work.Int.add(
                                                         \$19498_loop665_arg\(32 to 47), X"1770")) & eclat_false) & eclat_false));
                  if \$v5027\(0) = '1' then
                    \$19685\ := \$19684\ & \$19498_loop665_arg\(16 to 31);
                    \$v5010\ := \$ram_lock\;
                    if \$v5010\(0) = '1' then
                      state_var5921 := Q_WAIT5009;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                              \$19498_loop665_arg\(64 to 79), \$19498_loop665_arg\(0 to 15))));
                      \$ram_write\ <= \$19685\(0 to 31); \$ram_write_request\ <= '1';
                      state_var5921 := PAUSE_SET5008;
                    end if;
                  else
                    \$v5026\ := \$ram_lock\;
                    if \$v5026\(0) = '1' then
                      state_var5921 := Q_WAIT5025;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                        eclat_resize(\$19684\(0 to 30),16), X"000" & X"1")));
                      state_var5921 := PAUSE_GET5024;
                    end if;
                  end if;
                when PAUSE_GET5032 =>
                  \$19680\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$19498_loop665_id\ := "000000100100";
                  \$19498_loop665_arg\ := X"000" & X"1" & \$19499_aux664_arg\(16 to 31) & \$19499_aux664_arg\(32 to 47) & \$19499_aux664_arg\(48 to 63) & \$19499_aux664_arg\(0 to 15) & eclat_resize(
                  work.Int.lsr(eclat_resize(eclat_resize(\$19680\(0 to 30),16),31), X"0000000" & X"2"),16);
                  state_var5921 := \$19498_LOOP665\;
                when PAUSE_GET5049 =>
                  \$19560_hd\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$19561\ := work.Print.print_string(clk,of_string("bloc "));
                  \$19562\ := work.Int.print(clk,eclat_resize(\$19553\(0 to 30),16));
                  \$19563\ := work.Print.print_string(clk,of_string(" of size "));
                  \$19564\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                              work.Int.lsr(
                                                              \$19560_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$19565\ := work.Print.print_string(clk,of_string(" from "));
                  \$19566\ := work.Int.print(clk,eclat_resize(\$19553\(0 to 30),16));
                  \$19567\ := work.Print.print_string(clk,of_string(" to "));
                  \$19568\ := work.Int.print(clk,\$19547_copy_root_in_ram6634352_arg\(32 to 47));
                  \$19569\ := work.Print.print_newline(clk,eclat_unit);
                  \$v5048\ := \$ram_lock\;
                  if \$v5048\(0) = '1' then
                    state_var5921 := Q_WAIT5047;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19547_copy_root_in_ram6634352_arg\(32 to 47)));
                    \$ram_write\ <= \$19560_hd\; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5046;
                  end if;
                when PAUSE_GET5053 =>
                  \$19559_w\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v5052\ := eclat_if(work.Bool.lnot(""&\$19559_w\(31)) & 
                              eclat_if(work.Int.le(\$19547_copy_root_in_ram6634352_arg\(64 to 79), eclat_resize(\$19559_w\(0 to 30),16)) & 
                              work.Int.lt(eclat_resize(\$19559_w\(0 to 30),16), 
                                          work.Int.add(\$19547_copy_root_in_ram6634352_arg\(64 to 79), X"1770")) & eclat_false) & eclat_false);
                  if \$v5052\(0) = '1' then
                    \$19554\ := \$19559_w\ & \$19547_copy_root_in_ram6634352_arg\(32 to 47);
                    \$v5039\ := \$ram_lock\;
                    if \$v5039\(0) = '1' then
                      state_var5921 := Q_WAIT5038;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(\$19547_copy_root_in_ram6634352_arg\(0 to 15)));
                      \$ram_write\ <= \$19554\(0 to 31); \$ram_write_request\ <= '1';
                      state_var5921 := PAUSE_SET5037;
                    end if;
                  else
                    \$v5051\ := \$ram_lock\;
                    if \$v5051\(0) = '1' then
                      state_var5921 := Q_WAIT5050;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$19553\(0 to 30),16)));
                      state_var5921 := PAUSE_GET5049;
                    end if;
                  end if;
                when PAUSE_GET5057 =>
                  \$19553\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v5056\ := work.Bool.lnot(eclat_if(work.Bool.lnot(
                                                      ""&\$19553\(31)) & 
                                             eclat_if(work.Int.le(\$19547_copy_root_in_ram6634352_arg\(48 to 63), eclat_resize(\$19553\(0 to 30),16)) & 
                                             work.Int.lt(eclat_resize(\$19553\(0 to 30),16), 
                                                         work.Int.add(
                                                         \$19547_copy_root_in_ram6634352_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false));
                  if \$v5056\(0) = '1' then
                    \$19554\ := \$19553\ & \$19547_copy_root_in_ram6634352_arg\(32 to 47);
                    \$v5039\ := \$ram_lock\;
                    if \$v5039\(0) = '1' then
                      state_var5921 := Q_WAIT5038;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(\$19547_copy_root_in_ram6634352_arg\(0 to 15)));
                      \$ram_write\ <= \$19554\(0 to 31); \$ram_write_request\ <= '1';
                      state_var5921 := PAUSE_SET5037;
                    end if;
                  else
                    \$v5055\ := \$ram_lock\;
                    if \$v5055\(0) = '1' then
                      state_var5921 := Q_WAIT5054;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                        eclat_resize(\$19553\(0 to 30),16), X"000" & X"1")));
                      state_var5921 := PAUSE_GET5053;
                    end if;
                  end if;
                when PAUSE_GET5073 =>
                  \$19575_hd\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$19576\ := work.Print.print_string(clk,of_string("bloc "));
                  \$19577\ := work.Int.print(clk,eclat_resize(\$19541\(0 to 30),16));
                  \$19578\ := work.Print.print_string(clk,of_string(" of size "));
                  \$19579\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                              work.Int.lsr(
                                                              \$19575_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$19580\ := work.Print.print_string(clk,of_string(" from "));
                  \$19581\ := work.Int.print(clk,eclat_resize(\$19541\(0 to 30),16));
                  \$19582\ := work.Print.print_string(clk,of_string(" to "));
                  \$19583\ := work.Int.print(clk,\$19535_copy_root_in_ram6634354_arg\(32 to 47));
                  \$19584\ := work.Print.print_newline(clk,eclat_unit);
                  \$v5072\ := \$ram_lock\;
                  if \$v5072\(0) = '1' then
                    state_var5921 := Q_WAIT5071;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19535_copy_root_in_ram6634354_arg\(32 to 47)));
                    \$ram_write\ <= \$19575_hd\; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5070;
                  end if;
                when PAUSE_GET5077 =>
                  \$19574_w\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v5076\ := eclat_if(work.Bool.lnot(""&\$19574_w\(31)) & 
                              eclat_if(work.Int.le(\$19535_copy_root_in_ram6634354_arg\(64 to 79), eclat_resize(\$19574_w\(0 to 30),16)) & 
                              work.Int.lt(eclat_resize(\$19574_w\(0 to 30),16), 
                                          work.Int.add(\$19535_copy_root_in_ram6634354_arg\(64 to 79), X"1770")) & eclat_false) & eclat_false);
                  if \$v5076\(0) = '1' then
                    \$19542\ := \$19574_w\ & \$19535_copy_root_in_ram6634354_arg\(32 to 47);
                    \$v5063\ := \$ram_lock\;
                    if \$v5063\(0) = '1' then
                      state_var5921 := Q_WAIT5062;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(\$19535_copy_root_in_ram6634354_arg\(0 to 15)));
                      \$ram_write\ <= \$19542\(0 to 31); \$ram_write_request\ <= '1';
                      state_var5921 := PAUSE_SET5061;
                    end if;
                  else
                    \$v5075\ := \$ram_lock\;
                    if \$v5075\(0) = '1' then
                      state_var5921 := Q_WAIT5074;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$19541\(0 to 30),16)));
                      state_var5921 := PAUSE_GET5073;
                    end if;
                  end if;
                when PAUSE_GET5081 =>
                  \$19541\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v5080\ := work.Bool.lnot(eclat_if(work.Bool.lnot(
                                                      ""&\$19541\(31)) & 
                                             eclat_if(work.Int.le(\$19535_copy_root_in_ram6634354_arg\(48 to 63), eclat_resize(\$19541\(0 to 30),16)) & 
                                             work.Int.lt(eclat_resize(\$19541\(0 to 30),16), 
                                                         work.Int.add(
                                                         \$19535_copy_root_in_ram6634354_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false));
                  if \$v5080\(0) = '1' then
                    \$19542\ := \$19541\ & \$19535_copy_root_in_ram6634354_arg\(32 to 47);
                    \$v5063\ := \$ram_lock\;
                    if \$v5063\(0) = '1' then
                      state_var5921 := Q_WAIT5062;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(\$19535_copy_root_in_ram6634354_arg\(0 to 15)));
                      \$ram_write\ <= \$19542\(0 to 31); \$ram_write_request\ <= '1';
                      state_var5921 := PAUSE_SET5061;
                    end if;
                  else
                    \$v5079\ := \$ram_lock\;
                    if \$v5079\(0) = '1' then
                      state_var5921 := Q_WAIT5078;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                        eclat_resize(\$19541\(0 to 30),16), X"000" & X"1")));
                      state_var5921 := PAUSE_GET5077;
                    end if;
                  end if;
                when PAUSE_GET5085 =>
                  \$19514\ := \$global_end_value\;
                  release(\$global_end_lock\);
                  \$19535_copy_root_in_ram6634354_id\ := "000000101100";
                  \$19535_copy_root_in_ram6634354_arg\ := X"3e80" & \$19514\ & \$19507_next\ & \$19493\(96 to 111) & \$19493\(112 to 127);
                  state_var5921 := \$19535_COPY_ROOT_IN_RAM6634354\;
                when PAUSE_GET5100 =>
                  \$19614_hd\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$19615\ := work.Print.print_string(clk,of_string("bloc "));
                  \$19616\ := work.Int.print(clk,eclat_resize(\$19607\(0 to 30),16));
                  \$19617\ := work.Print.print_string(clk,of_string(" of size "));
                  \$19618\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                              work.Int.lsr(
                                                              \$19614_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$19619\ := work.Print.print_string(clk,of_string(" from "));
                  \$19620\ := work.Int.print(clk,eclat_resize(\$19607\(0 to 30),16));
                  \$19621\ := work.Print.print_string(clk,of_string(" to "));
                  \$19622\ := work.Int.print(clk,\$19601_copy_root_in_ram6634352_arg\(32 to 47));
                  \$19623\ := work.Print.print_newline(clk,eclat_unit);
                  \$v5099\ := \$ram_lock\;
                  if \$v5099\(0) = '1' then
                    state_var5921 := Q_WAIT5098;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19601_copy_root_in_ram6634352_arg\(32 to 47)));
                    \$ram_write\ <= \$19614_hd\; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5097;
                  end if;
                when PAUSE_GET5104 =>
                  \$19613_w\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v5103\ := eclat_if(work.Bool.lnot(""&\$19613_w\(31)) & 
                              eclat_if(work.Int.le(\$19601_copy_root_in_ram6634352_arg\(64 to 79), eclat_resize(\$19613_w\(0 to 30),16)) & 
                              work.Int.lt(eclat_resize(\$19613_w\(0 to 30),16), 
                                          work.Int.add(\$19601_copy_root_in_ram6634352_arg\(64 to 79), X"1770")) & eclat_false) & eclat_false);
                  if \$v5103\(0) = '1' then
                    \$19608\ := \$19613_w\ & \$19601_copy_root_in_ram6634352_arg\(32 to 47);
                    \$v5090\ := \$ram_lock\;
                    if \$v5090\(0) = '1' then
                      state_var5921 := Q_WAIT5089;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(\$19601_copy_root_in_ram6634352_arg\(0 to 15)));
                      \$ram_write\ <= \$19608\(0 to 31); \$ram_write_request\ <= '1';
                      state_var5921 := PAUSE_SET5088;
                    end if;
                  else
                    \$v5102\ := \$ram_lock\;
                    if \$v5102\(0) = '1' then
                      state_var5921 := Q_WAIT5101;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$19607\(0 to 30),16)));
                      state_var5921 := PAUSE_GET5100;
                    end if;
                  end if;
                when PAUSE_GET5108 =>
                  \$19607\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v5107\ := work.Bool.lnot(eclat_if(work.Bool.lnot(
                                                      ""&\$19607\(31)) & 
                                             eclat_if(work.Int.le(\$19601_copy_root_in_ram6634352_arg\(48 to 63), eclat_resize(\$19607\(0 to 30),16)) & 
                                             work.Int.lt(eclat_resize(\$19607\(0 to 30),16), 
                                                         work.Int.add(
                                                         \$19601_copy_root_in_ram6634352_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false));
                  if \$v5107\(0) = '1' then
                    \$19608\ := \$19607\ & \$19601_copy_root_in_ram6634352_arg\(32 to 47);
                    \$v5090\ := \$ram_lock\;
                    if \$v5090\(0) = '1' then
                      state_var5921 := Q_WAIT5089;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(\$19601_copy_root_in_ram6634352_arg\(0 to 15)));
                      \$ram_write\ <= \$19608\(0 to 31); \$ram_write_request\ <= '1';
                      state_var5921 := PAUSE_SET5088;
                    end if;
                  else
                    \$v5106\ := \$ram_lock\;
                    if \$v5106\(0) = '1' then
                      state_var5921 := Q_WAIT5105;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                        eclat_resize(\$19607\(0 to 30),16), X"000" & X"1")));
                      state_var5921 := PAUSE_GET5104;
                    end if;
                  end if;
                when PAUSE_GET5124 =>
                  \$19629_hd\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$19630\ := work.Print.print_string(clk,of_string("bloc "));
                  \$19631\ := work.Int.print(clk,eclat_resize(\$19595\(0 to 30),16));
                  \$19632\ := work.Print.print_string(clk,of_string(" of size "));
                  \$19633\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                              work.Int.lsr(
                                                              \$19629_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$19634\ := work.Print.print_string(clk,of_string(" from "));
                  \$19635\ := work.Int.print(clk,eclat_resize(\$19595\(0 to 30),16));
                  \$19636\ := work.Print.print_string(clk,of_string(" to "));
                  \$19637\ := work.Int.print(clk,\$19589_copy_root_in_ram6634353_arg\(32 to 47));
                  \$19638\ := work.Print.print_newline(clk,eclat_unit);
                  \$v5123\ := \$ram_lock\;
                  if \$v5123\(0) = '1' then
                    state_var5921 := Q_WAIT5122;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19589_copy_root_in_ram6634353_arg\(32 to 47)));
                    \$ram_write\ <= \$19629_hd\; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5121;
                  end if;
                when PAUSE_GET5128 =>
                  \$19628_w\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v5127\ := eclat_if(work.Bool.lnot(""&\$19628_w\(31)) & 
                              eclat_if(work.Int.le(\$19589_copy_root_in_ram6634353_arg\(64 to 79), eclat_resize(\$19628_w\(0 to 30),16)) & 
                              work.Int.lt(eclat_resize(\$19628_w\(0 to 30),16), 
                                          work.Int.add(\$19589_copy_root_in_ram6634353_arg\(64 to 79), X"1770")) & eclat_false) & eclat_false);
                  if \$v5127\(0) = '1' then
                    \$19596\ := \$19628_w\ & \$19589_copy_root_in_ram6634353_arg\(32 to 47);
                    \$v5114\ := \$ram_lock\;
                    if \$v5114\(0) = '1' then
                      state_var5921 := Q_WAIT5113;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(\$19589_copy_root_in_ram6634353_arg\(0 to 15)));
                      \$ram_write\ <= \$19596\(0 to 31); \$ram_write_request\ <= '1';
                      state_var5921 := PAUSE_SET5112;
                    end if;
                  else
                    \$v5126\ := \$ram_lock\;
                    if \$v5126\(0) = '1' then
                      state_var5921 := Q_WAIT5125;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$19595\(0 to 30),16)));
                      state_var5921 := PAUSE_GET5124;
                    end if;
                  end if;
                when PAUSE_GET5132 =>
                  \$19595\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v5131\ := work.Bool.lnot(eclat_if(work.Bool.lnot(
                                                      ""&\$19595\(31)) & 
                                             eclat_if(work.Int.le(\$19589_copy_root_in_ram6634353_arg\(48 to 63), eclat_resize(\$19595\(0 to 30),16)) & 
                                             work.Int.lt(eclat_resize(\$19595\(0 to 30),16), 
                                                         work.Int.add(
                                                         \$19589_copy_root_in_ram6634353_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false));
                  if \$v5131\(0) = '1' then
                    \$19596\ := \$19595\ & \$19589_copy_root_in_ram6634353_arg\(32 to 47);
                    \$v5114\ := \$ram_lock\;
                    if \$v5114\(0) = '1' then
                      state_var5921 := Q_WAIT5113;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(\$19589_copy_root_in_ram6634353_arg\(0 to 15)));
                      \$ram_write\ <= \$19596\(0 to 31); \$ram_write_request\ <= '1';
                      state_var5921 := PAUSE_SET5112;
                    end if;
                  else
                    \$v5130\ := \$ram_lock\;
                    if \$v5130\(0) = '1' then
                      state_var5921 := Q_WAIT5129;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                        eclat_resize(\$19595\(0 to 30),16), X"000" & X"1")));
                      state_var5921 := PAUSE_GET5128;
                    end if;
                  end if;
                when PAUSE_GET5145 =>
                  \$19644_hd\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$19645\ := work.Print.print_string(clk,of_string("bloc "));
                  \$19646\ := work.Int.print(clk,eclat_resize(\$18792_wait662_arg\(33 to 63),16));
                  \$19647\ := work.Print.print_string(clk,of_string(" of size "));
                  \$19648\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                              work.Int.lsr(
                                                              \$19644_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$19649\ := work.Print.print_string(clk,of_string(" from "));
                  \$19650\ := work.Int.print(clk,eclat_resize(\$18792_wait662_arg\(33 to 63),16));
                  \$19651\ := work.Print.print_string(clk,of_string(" to "));
                  \$19652\ := work.Int.print(clk,\$19505\(32 to 47));
                  \$19653\ := work.Print.print_newline(clk,eclat_unit);
                  \$v5144\ := \$ram_lock\;
                  if \$v5144\(0) = '1' then
                    state_var5921 := Q_WAIT5143;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19505\(32 to 47)));
                    \$ram_write\ <= \$19644_hd\; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5142;
                  end if;
                when PAUSE_GET5149 =>
                  \$19643_w\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v5148\ := eclat_if(work.Bool.lnot(""&\$19643_w\(31)) & 
                              eclat_if(work.Int.le(\$19493\(112 to 127), eclat_resize(\$19643_w\(0 to 30),16)) & 
                              work.Int.lt(eclat_resize(\$19643_w\(0 to 30),16), 
                                          work.Int.add(\$19493\(112 to 127), X"1770")) & eclat_false) & eclat_false);
                  if \$v5148\(0) = '1' then
                    \$19506\ := \$19643_w\ & \$19505\(32 to 47);
                    \$19589_copy_root_in_ram6634353_id\ := "000000110000";
                    \$19589_copy_root_in_ram6634353_arg\ := X"0" & X"3e8" & \$18792_wait662_arg\(65 to 80) & \$19506\(32 to 47) & \$19493\(96 to 111) & \$19493\(112 to 127);
                    state_var5921 := \$19589_COPY_ROOT_IN_RAM6634353\;
                  else
                    \$v5147\ := \$ram_lock\;
                    if \$v5147\(0) = '1' then
                      state_var5921 := Q_WAIT5146;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18792_wait662_arg\(33 to 63),16)));
                      state_var5921 := PAUSE_GET5145;
                    end if;
                  end if;
                when PAUSE_GET5162 =>
                  \$19659_hd\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$19660\ := work.Print.print_string(clk,of_string("bloc "));
                  \$19661\ := work.Int.print(clk,eclat_resize(\$18792_wait662_arg\(1 to 31),16));
                  \$19662\ := work.Print.print_string(clk,of_string(" of size "));
                  \$19663\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                              work.Int.lsr(
                                                              \$19659_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$19664\ := work.Print.print_string(clk,of_string(" from "));
                  \$19665\ := work.Int.print(clk,eclat_resize(\$18792_wait662_arg\(1 to 31),16));
                  \$19666\ := work.Print.print_string(clk,of_string(" to "));
                  \$19667\ := work.Int.print(clk,\$19493\(112 to 127));
                  \$19668\ := work.Print.print_newline(clk,eclat_unit);
                  \$v5161\ := \$ram_lock\;
                  if \$v5161\(0) = '1' then
                    state_var5921 := Q_WAIT5160;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19493\(112 to 127)));
                    \$ram_write\ <= \$19659_hd\; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5159;
                  end if;
                when PAUSE_GET5166 =>
                  \$19658_w\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v5165\ := eclat_if(work.Bool.lnot(""&\$19658_w\(31)) & 
                              eclat_if(work.Int.le(\$19493\(112 to 127), eclat_resize(\$19658_w\(0 to 30),16)) & 
                              work.Int.lt(eclat_resize(\$19658_w\(0 to 30),16), 
                                          work.Int.add(\$19493\(112 to 127), X"1770")) & eclat_false) & eclat_false);
                  if \$v5165\(0) = '1' then
                    \$19505\ := \$19658_w\ & \$19493\(112 to 127);
                    \$v5152\ := work.Bool.lnot(eclat_if(work.Bool.lnot(
                                                        ""&\$18792_wait662_arg\(64)) & 
                                               eclat_if(work.Int.le(\$19493\(96 to 111), eclat_resize(\$18792_wait662_arg\(33 to 63),16)) & 
                                               work.Int.lt(eclat_resize(\$18792_wait662_arg\(33 to 63),16), 
                                                           work.Int.add(
                                                           \$19493\(96 to 111), X"1770")) & eclat_false) & eclat_false));
                    if \$v5152\(0) = '1' then
                      \$19506\ := \$18792_wait662_arg\(33 to 64) & \$19505\(32 to 47);
                      \$19589_copy_root_in_ram6634353_id\ := "000000110000";
                      \$19589_copy_root_in_ram6634353_arg\ := X"0" & X"3e8" & \$18792_wait662_arg\(65 to 80) & \$19506\(32 to 47) & \$19493\(96 to 111) & \$19493\(112 to 127);
                      state_var5921 := \$19589_COPY_ROOT_IN_RAM6634353\;
                    else
                      \$v5151\ := \$ram_lock\;
                      if \$v5151\(0) = '1' then
                        state_var5921 := Q_WAIT5150;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$18792_wait662_arg\(33 to 63),16), X"000" & X"1")));
                        state_var5921 := PAUSE_GET5149;
                      end if;
                    end if;
                  else
                    \$v5164\ := \$ram_lock\;
                    if \$v5164\(0) = '1' then
                      state_var5921 := Q_WAIT5163;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18792_wait662_arg\(1 to 31),16)));
                      state_var5921 := PAUSE_GET5162;
                    end if;
                  end if;
                when PAUSE_SET4966 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19738\ := eclat_unit;
                  \$19494_loop666_arg\ := work.Int.add(\$19494_loop666_arg\(0 to 15), X"000" & X"1") & \$19494_loop666_arg\(16 to 31) & \$19494_loop666_arg\(32 to 47) & \$19494_loop666_arg\(48 to 63);
                  state_var5921 := \$19494_LOOP666\;
                when PAUSE_SET4973 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19719\ := eclat_unit;
                  \$19495_loop665_arg\ := work.Int.add(\$19495_loop665_arg\(0 to 15), X"000" & X"1") & \$19718\(32 to 47) & \$19495_loop665_arg\(32 to 47) & \$19495_loop665_arg\(48 to 63) & \$19495_loop665_arg\(64 to 79) & \$19495_loop665_arg\(80 to 95);
                  state_var5921 := \$19495_LOOP665\;
                when PAUSE_SET4976 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19734\ := eclat_unit;
                  \$19718\ := eclat_resize(\$19495_loop665_arg\(16 to 31),31) & eclat_false & 
                  work.Int.add(\$19495_loop665_arg\(16 to 31), work.Int.add(
                                                               eclat_resize(
                                                               work.Int.lsr(
                                                               \$19721_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$v4975\ := \$ram_lock\;
                  if \$v4975\(0) = '1' then
                    state_var5921 := Q_WAIT4974;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            \$19495_loop665_arg\(64 to 79), \$19495_loop665_arg\(0 to 15))));
                    \$ram_write\ <= \$19718\(0 to 31); \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET4973;
                  end if;
                when PAUSE_SET4979 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19733\ := eclat_unit;
                  \$v4978\ := \$ram_lock\;
                  if \$v4978\(0) = '1' then
                    state_var5921 := Q_WAIT4977;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$19717\(0 to 30),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$19495_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET4976;
                  end if;
                when PAUSE_SET4982 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19731\ := eclat_unit;
                  \$19494_loop666_id\ := "000000100001";
                  \$19494_loop666_arg\ := X"000" & X"1" & \$19495_loop665_arg\(16 to 31) & eclat_resize(\$19717\(0 to 30),16) & eclat_resize(
                  work.Int.lsr(\$19721_hd\(0 to 30), X"0000000" & X"2"),16);
                  state_var5921 := \$19494_LOOP666\;
                when PAUSE_SET5001 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19705\ := eclat_unit;
                  \$19497_loop666_arg\ := work.Int.add(\$19497_loop666_arg\(0 to 15), X"000" & X"1") & \$19497_loop666_arg\(16 to 31) & \$19497_loop666_arg\(32 to 47) & \$19497_loop666_arg\(48 to 63);
                  state_var5921 := \$19497_LOOP666\;
                when PAUSE_SET5008 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19686\ := eclat_unit;
                  \$19498_loop665_arg\ := work.Int.add(\$19498_loop665_arg\(0 to 15), X"000" & X"1") & \$19685\(32 to 47) & \$19498_loop665_arg\(32 to 47) & \$19498_loop665_arg\(48 to 63) & \$19498_loop665_arg\(64 to 79) & \$19498_loop665_arg\(80 to 95);
                  state_var5921 := \$19498_LOOP665\;
                when PAUSE_SET5011 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19701\ := eclat_unit;
                  \$19685\ := eclat_resize(\$19498_loop665_arg\(16 to 31),31) & eclat_false & 
                  work.Int.add(\$19498_loop665_arg\(16 to 31), work.Int.add(
                                                               eclat_resize(
                                                               work.Int.lsr(
                                                               \$19688_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$v5010\ := \$ram_lock\;
                  if \$v5010\(0) = '1' then
                    state_var5921 := Q_WAIT5009;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            \$19498_loop665_arg\(64 to 79), \$19498_loop665_arg\(0 to 15))));
                    \$ram_write\ <= \$19685\(0 to 31); \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5008;
                  end if;
                when PAUSE_SET5014 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19700\ := eclat_unit;
                  \$v5013\ := \$ram_lock\;
                  if \$v5013\(0) = '1' then
                    state_var5921 := Q_WAIT5012;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$19684\(0 to 30),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$19498_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5011;
                  end if;
                when PAUSE_SET5017 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19698\ := eclat_unit;
                  \$19497_loop666_id\ := "000000100011";
                  \$19497_loop666_arg\ := X"000" & X"1" & \$19498_loop665_arg\(16 to 31) & eclat_resize(\$19684\(0 to 30),16) & eclat_resize(
                  work.Int.lsr(\$19688_hd\(0 to 30), X"0000000" & X"2"),16);
                  state_var5921 := \$19497_LOOP666\;
                when PAUSE_SET5037 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19555\ := eclat_unit;
                  \$19556\ := work.Print.print_string(clk,of_string(" next="));
                  \$19557\ := work.Int.print(clk,\$19554\(32 to 47));
                  \$19558\ := work.Print.print_newline(clk,eclat_unit);
                  \$19547_copy_root_in_ram6634352_arg\ := work.Int.add(
                                                          \$19547_copy_root_in_ram6634352_arg\(0 to 15), X"000" & X"1") & \$19547_copy_root_in_ram6634352_arg\(16 to 31) & \$19554\(32 to 47) & \$19547_copy_root_in_ram6634352_arg\(48 to 63) & \$19547_copy_root_in_ram6634352_arg\(64 to 79);
                  state_var5921 := \$19547_COPY_ROOT_IN_RAM6634352\;
                when PAUSE_SET5040 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19573\ := eclat_unit;
                  \$19554\ := eclat_resize(\$19547_copy_root_in_ram6634352_arg\(32 to 47),31) & eclat_false & 
                  work.Int.add(\$19547_copy_root_in_ram6634352_arg\(32 to 47), 
                               work.Int.add(eclat_resize(work.Int.lsr(
                                                         \$19560_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$v5039\ := \$ram_lock\;
                  if \$v5039\(0) = '1' then
                    state_var5921 := Q_WAIT5038;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19547_copy_root_in_ram6634352_arg\(0 to 15)));
                    \$ram_write\ <= \$19554\(0 to 31); \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5037;
                  end if;
                when PAUSE_SET5043 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19572\ := eclat_unit;
                  \$v5042\ := \$ram_lock\;
                  if \$v5042\(0) = '1' then
                    state_var5921 := Q_WAIT5041;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$19553\(0 to 30),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$19547_copy_root_in_ram6634352_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5040;
                  end if;
                when PAUSE_SET5046 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19570\ := eclat_unit;
                  \$19497_loop666_id\ := "000000101001";
                  \$19497_loop666_arg\ := X"000" & X"1" & \$19547_copy_root_in_ram6634352_arg\(32 to 47) & eclat_resize(\$19553\(0 to 30),16) & eclat_resize(
                  work.Int.lsr(\$19560_hd\(0 to 30), X"0000000" & X"2"),16);
                  state_var5921 := \$19497_LOOP666\;
                when PAUSE_SET5061 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19543\ := eclat_unit;
                  \$19544\ := work.Print.print_string(clk,of_string(" next="));
                  \$19545\ := work.Int.print(clk,\$19542\(32 to 47));
                  \$19546\ := work.Print.print_newline(clk,eclat_unit);
                  \$19547_copy_root_in_ram6634352_id\ := "000000101010";
                  \$19547_copy_root_in_ram6634352_arg\ := work.Int.add(
                                                          \$19535_copy_root_in_ram6634354_arg\(0 to 15), X"000" & X"1") & \$19535_copy_root_in_ram6634354_arg\(16 to 31) & \$19542\(32 to 47) & \$19535_copy_root_in_ram6634354_arg\(48 to 63) & \$19535_copy_root_in_ram6634354_arg\(64 to 79);
                  state_var5921 := \$19547_COPY_ROOT_IN_RAM6634352\;
                when PAUSE_SET5064 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19588\ := eclat_unit;
                  \$19542\ := eclat_resize(\$19535_copy_root_in_ram6634354_arg\(32 to 47),31) & eclat_false & 
                  work.Int.add(\$19535_copy_root_in_ram6634354_arg\(32 to 47), 
                               work.Int.add(eclat_resize(work.Int.lsr(
                                                         \$19575_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$v5063\ := \$ram_lock\;
                  if \$v5063\(0) = '1' then
                    state_var5921 := Q_WAIT5062;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19535_copy_root_in_ram6634354_arg\(0 to 15)));
                    \$ram_write\ <= \$19542\(0 to 31); \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5061;
                  end if;
                when PAUSE_SET5067 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19587\ := eclat_unit;
                  \$v5066\ := \$ram_lock\;
                  if \$v5066\(0) = '1' then
                    state_var5921 := Q_WAIT5065;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$19541\(0 to 30),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$19535_copy_root_in_ram6634354_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5064;
                  end if;
                when PAUSE_SET5070 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19585\ := eclat_unit;
                  \$19497_loop666_id\ := "000000101011";
                  \$19497_loop666_arg\ := X"000" & X"1" & \$19535_copy_root_in_ram6634354_arg\(32 to 47) & eclat_resize(\$19541\(0 to 30),16) & eclat_resize(
                  work.Int.lsr(\$19575_hd\(0 to 30), X"0000000" & X"2"),16);
                  state_var5921 := \$19497_LOOP666\;
                when PAUSE_SET5088 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19609\ := eclat_unit;
                  \$19610\ := work.Print.print_string(clk,of_string(" next="));
                  \$19611\ := work.Int.print(clk,\$19608\(32 to 47));
                  \$19612\ := work.Print.print_newline(clk,eclat_unit);
                  \$19601_copy_root_in_ram6634352_arg\ := work.Int.add(
                                                          \$19601_copy_root_in_ram6634352_arg\(0 to 15), X"000" & X"1") & \$19601_copy_root_in_ram6634352_arg\(16 to 31) & \$19608\(32 to 47) & \$19601_copy_root_in_ram6634352_arg\(48 to 63) & \$19601_copy_root_in_ram6634352_arg\(64 to 79);
                  state_var5921 := \$19601_COPY_ROOT_IN_RAM6634352\;
                when PAUSE_SET5091 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19627\ := eclat_unit;
                  \$19608\ := eclat_resize(\$19601_copy_root_in_ram6634352_arg\(32 to 47),31) & eclat_false & 
                  work.Int.add(\$19601_copy_root_in_ram6634352_arg\(32 to 47), 
                               work.Int.add(eclat_resize(work.Int.lsr(
                                                         \$19614_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$v5090\ := \$ram_lock\;
                  if \$v5090\(0) = '1' then
                    state_var5921 := Q_WAIT5089;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19601_copy_root_in_ram6634352_arg\(0 to 15)));
                    \$ram_write\ <= \$19608\(0 to 31); \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5088;
                  end if;
                when PAUSE_SET5094 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19626\ := eclat_unit;
                  \$v5093\ := \$ram_lock\;
                  if \$v5093\(0) = '1' then
                    state_var5921 := Q_WAIT5092;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$19607\(0 to 30),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$19601_copy_root_in_ram6634352_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5091;
                  end if;
                when PAUSE_SET5097 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19624\ := eclat_unit;
                  \$19497_loop666_id\ := "000000101101";
                  \$19497_loop666_arg\ := X"000" & X"1" & \$19601_copy_root_in_ram6634352_arg\(32 to 47) & eclat_resize(\$19607\(0 to 30),16) & eclat_resize(
                  work.Int.lsr(\$19614_hd\(0 to 30), X"0000000" & X"2"),16);
                  state_var5921 := \$19497_LOOP666\;
                when PAUSE_SET5112 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19597\ := eclat_unit;
                  \$19598\ := work.Print.print_string(clk,of_string(" next="));
                  \$19599\ := work.Int.print(clk,\$19596\(32 to 47));
                  \$19600\ := work.Print.print_newline(clk,eclat_unit);
                  \$19601_copy_root_in_ram6634352_id\ := "000000101110";
                  \$19601_copy_root_in_ram6634352_arg\ := work.Int.add(
                                                          \$19589_copy_root_in_ram6634353_arg\(0 to 15), X"000" & X"1") & \$19589_copy_root_in_ram6634353_arg\(16 to 31) & \$19596\(32 to 47) & \$19589_copy_root_in_ram6634353_arg\(48 to 63) & \$19589_copy_root_in_ram6634353_arg\(64 to 79);
                  state_var5921 := \$19601_COPY_ROOT_IN_RAM6634352\;
                when PAUSE_SET5115 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19642\ := eclat_unit;
                  \$19596\ := eclat_resize(\$19589_copy_root_in_ram6634353_arg\(32 to 47),31) & eclat_false & 
                  work.Int.add(\$19589_copy_root_in_ram6634353_arg\(32 to 47), 
                               work.Int.add(eclat_resize(work.Int.lsr(
                                                         \$19629_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$v5114\ := \$ram_lock\;
                  if \$v5114\(0) = '1' then
                    state_var5921 := Q_WAIT5113;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19589_copy_root_in_ram6634353_arg\(0 to 15)));
                    \$ram_write\ <= \$19596\(0 to 31); \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5112;
                  end if;
                when PAUSE_SET5118 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19641\ := eclat_unit;
                  \$v5117\ := \$ram_lock\;
                  if \$v5117\(0) = '1' then
                    state_var5921 := Q_WAIT5116;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$19595\(0 to 30),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$19589_copy_root_in_ram6634353_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5115;
                  end if;
                when PAUSE_SET5121 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19639\ := eclat_unit;
                  \$19497_loop666_id\ := "000000101111";
                  \$19497_loop666_arg\ := X"000" & X"1" & \$19589_copy_root_in_ram6634353_arg\(32 to 47) & eclat_resize(\$19595\(0 to 30),16) & eclat_resize(
                  work.Int.lsr(\$19629_hd\(0 to 30), X"0000000" & X"2"),16);
                  state_var5921 := \$19497_LOOP666\;
                when PAUSE_SET5136 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19657\ := eclat_unit;
                  \$19506\ := eclat_resize(\$19505\(32 to 47),31) & eclat_false & 
                  work.Int.add(\$19505\(32 to 47), work.Int.add(eclat_resize(
                                                                work.Int.lsr(
                                                                \$19644_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$19589_copy_root_in_ram6634353_id\ := "000000110000";
                  \$19589_copy_root_in_ram6634353_arg\ := X"0" & X"3e8" & \$18792_wait662_arg\(65 to 80) & \$19506\(32 to 47) & \$19493\(96 to 111) & \$19493\(112 to 127);
                  state_var5921 := \$19589_COPY_ROOT_IN_RAM6634353\;
                when PAUSE_SET5139 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19656\ := eclat_unit;
                  \$v5138\ := \$ram_lock\;
                  if \$v5138\(0) = '1' then
                    state_var5921 := Q_WAIT5137;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$18792_wait662_arg\(33 to 63),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$19505\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5136;
                  end if;
                when PAUSE_SET5142 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19654\ := eclat_unit;
                  \$19497_loop666_id\ := "000000110001";
                  \$19497_loop666_arg\ := X"000" & X"1" & \$19505\(32 to 47) & eclat_resize(\$18792_wait662_arg\(33 to 63),16) & eclat_resize(
                  work.Int.lsr(\$19644_hd\(0 to 30), X"0000000" & X"2"),16);
                  state_var5921 := \$19497_LOOP666\;
                when PAUSE_SET5153 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19672\ := eclat_unit;
                  \$19505\ := eclat_resize(\$19493\(112 to 127),31) & eclat_false & 
                  work.Int.add(\$19493\(112 to 127), work.Int.add(eclat_resize(
                                                                  work.Int.lsr(
                                                                  \$19659_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$v5152\ := work.Bool.lnot(eclat_if(work.Bool.lnot(
                                                      ""&\$18792_wait662_arg\(64)) & 
                                             eclat_if(work.Int.le(\$19493\(96 to 111), eclat_resize(\$18792_wait662_arg\(33 to 63),16)) & 
                                             work.Int.lt(eclat_resize(\$18792_wait662_arg\(33 to 63),16), 
                                                         work.Int.add(
                                                         \$19493\(96 to 111), X"1770")) & eclat_false) & eclat_false));
                  if \$v5152\(0) = '1' then
                    \$19506\ := \$18792_wait662_arg\(33 to 64) & \$19505\(32 to 47);
                    \$19589_copy_root_in_ram6634353_id\ := "000000110000";
                    \$19589_copy_root_in_ram6634353_arg\ := X"0" & X"3e8" & \$18792_wait662_arg\(65 to 80) & \$19506\(32 to 47) & \$19493\(96 to 111) & \$19493\(112 to 127);
                    state_var5921 := \$19589_COPY_ROOT_IN_RAM6634353\;
                  else
                    \$v5151\ := \$ram_lock\;
                    if \$v5151\(0) = '1' then
                      state_var5921 := Q_WAIT5150;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                        eclat_resize(\$18792_wait662_arg\(33 to 63),16), X"000" & X"1")));
                      state_var5921 := PAUSE_GET5149;
                    end if;
                  end if;
                when PAUSE_SET5156 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19671\ := eclat_unit;
                  \$v5155\ := \$ram_lock\;
                  if \$v5155\(0) = '1' then
                    state_var5921 := Q_WAIT5154;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$18792_wait662_arg\(1 to 31),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$19493\(112 to 127),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5153;
                  end if;
                when PAUSE_SET5159 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$19669\ := eclat_unit;
                  \$19497_loop666_id\ := "000000110010";
                  \$19497_loop666_arg\ := X"000" & X"1" & \$19493\(112 to 127) & eclat_resize(\$18792_wait662_arg\(1 to 31),16) & eclat_resize(
                  work.Int.lsr(\$19659_hd\(0 to 30), X"0000000" & X"2"),16);
                  state_var5921 := \$19497_LOOP666\;
                when Q_WAIT4967 =>
                  \$v4968\ := \$ram_lock\;
                  if \$v4968\(0) = '1' then
                    state_var5921 := Q_WAIT4967;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            \$19494_loop666_arg\(16 to 31), \$19494_loop666_arg\(0 to 15))));
                    \$ram_write\ <= \$19737\; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET4966;
                  end if;
                when Q_WAIT4970 =>
                  \$v4971\ := \$ram_lock\;
                  if \$v4971\(0) = '1' then
                    state_var5921 := Q_WAIT4970;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$19494_loop666_arg\(32 to 47), \$19494_loop666_arg\(0 to 15))));
                    state_var5921 := PAUSE_GET4969;
                  end if;
                when Q_WAIT4974 =>
                  \$v4975\ := \$ram_lock\;
                  if \$v4975\(0) = '1' then
                    state_var5921 := Q_WAIT4974;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            \$19495_loop665_arg\(64 to 79), \$19495_loop665_arg\(0 to 15))));
                    \$ram_write\ <= \$19718\(0 to 31); \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET4973;
                  end if;
                when Q_WAIT4977 =>
                  \$v4978\ := \$ram_lock\;
                  if \$v4978\(0) = '1' then
                    state_var5921 := Q_WAIT4977;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$19717\(0 to 30),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$19495_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET4976;
                  end if;
                when Q_WAIT4980 =>
                  \$v4981\ := \$ram_lock\;
                  if \$v4981\(0) = '1' then
                    state_var5921 := Q_WAIT4980;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$19717\(0 to 30),16)));
                    \$ram_write\ <= eclat_resize(\$19495_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET4979;
                  end if;
                when Q_WAIT4983 =>
                  \$v4984\ := \$ram_lock\;
                  if \$v4984\(0) = '1' then
                    state_var5921 := Q_WAIT4983;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19495_loop665_arg\(16 to 31)));
                    \$ram_write\ <= \$19721_hd\; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET4982;
                  end if;
                when Q_WAIT4986 =>
                  \$v4987\ := \$ram_lock\;
                  if \$v4987\(0) = '1' then
                    state_var5921 := Q_WAIT4986;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$19717\(0 to 30),16)));
                    state_var5921 := PAUSE_GET4985;
                  end if;
                when Q_WAIT4990 =>
                  \$v4991\ := \$ram_lock\;
                  if \$v4991\(0) = '1' then
                    state_var5921 := Q_WAIT4990;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19717\(0 to 30),16), X"000" & X"1")));
                    state_var5921 := PAUSE_GET4989;
                  end if;
                when Q_WAIT4994 =>
                  \$v4995\ := \$ram_lock\;
                  if \$v4995\(0) = '1' then
                    state_var5921 := Q_WAIT4994;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$19495_loop665_arg\(64 to 79), \$19495_loop665_arg\(0 to 15))));
                    state_var5921 := PAUSE_GET4993;
                  end if;
                when Q_WAIT4998 =>
                  \$v4999\ := \$ram_lock\;
                  if \$v4999\(0) = '1' then
                    state_var5921 := Q_WAIT4998;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(\$19496_aux664_arg\(0 to 15)));
                    state_var5921 := PAUSE_GET4997;
                  end if;
                when Q_WAIT5002 =>
                  \$v5003\ := \$ram_lock\;
                  if \$v5003\(0) = '1' then
                    state_var5921 := Q_WAIT5002;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            \$19497_loop666_arg\(16 to 31), \$19497_loop666_arg\(0 to 15))));
                    \$ram_write\ <= \$19704\; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5001;
                  end if;
                when Q_WAIT5005 =>
                  \$v5006\ := \$ram_lock\;
                  if \$v5006\(0) = '1' then
                    state_var5921 := Q_WAIT5005;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$19497_loop666_arg\(32 to 47), \$19497_loop666_arg\(0 to 15))));
                    state_var5921 := PAUSE_GET5004;
                  end if;
                when Q_WAIT5009 =>
                  \$v5010\ := \$ram_lock\;
                  if \$v5010\(0) = '1' then
                    state_var5921 := Q_WAIT5009;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            \$19498_loop665_arg\(64 to 79), \$19498_loop665_arg\(0 to 15))));
                    \$ram_write\ <= \$19685\(0 to 31); \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5008;
                  end if;
                when Q_WAIT5012 =>
                  \$v5013\ := \$ram_lock\;
                  if \$v5013\(0) = '1' then
                    state_var5921 := Q_WAIT5012;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$19684\(0 to 30),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$19498_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5011;
                  end if;
                when Q_WAIT5015 =>
                  \$v5016\ := \$ram_lock\;
                  if \$v5016\(0) = '1' then
                    state_var5921 := Q_WAIT5015;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$19684\(0 to 30),16)));
                    \$ram_write\ <= eclat_resize(\$19498_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5014;
                  end if;
                when Q_WAIT5018 =>
                  \$v5019\ := \$ram_lock\;
                  if \$v5019\(0) = '1' then
                    state_var5921 := Q_WAIT5018;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19498_loop665_arg\(16 to 31)));
                    \$ram_write\ <= \$19688_hd\; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5017;
                  end if;
                when Q_WAIT5021 =>
                  \$v5022\ := \$ram_lock\;
                  if \$v5022\(0) = '1' then
                    state_var5921 := Q_WAIT5021;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$19684\(0 to 30),16)));
                    state_var5921 := PAUSE_GET5020;
                  end if;
                when Q_WAIT5025 =>
                  \$v5026\ := \$ram_lock\;
                  if \$v5026\(0) = '1' then
                    state_var5921 := Q_WAIT5025;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19684\(0 to 30),16), X"000" & X"1")));
                    state_var5921 := PAUSE_GET5024;
                  end if;
                when Q_WAIT5029 =>
                  \$v5030\ := \$ram_lock\;
                  if \$v5030\(0) = '1' then
                    state_var5921 := Q_WAIT5029;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$19498_loop665_arg\(64 to 79), \$19498_loop665_arg\(0 to 15))));
                    state_var5921 := PAUSE_GET5028;
                  end if;
                when Q_WAIT5033 =>
                  \$v5034\ := \$ram_lock\;
                  if \$v5034\(0) = '1' then
                    state_var5921 := Q_WAIT5033;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(\$19499_aux664_arg\(0 to 15)));
                    state_var5921 := PAUSE_GET5032;
                  end if;
                when Q_WAIT5038 =>
                  \$v5039\ := \$ram_lock\;
                  if \$v5039\(0) = '1' then
                    state_var5921 := Q_WAIT5038;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19547_copy_root_in_ram6634352_arg\(0 to 15)));
                    \$ram_write\ <= \$19554\(0 to 31); \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5037;
                  end if;
                when Q_WAIT5041 =>
                  \$v5042\ := \$ram_lock\;
                  if \$v5042\(0) = '1' then
                    state_var5921 := Q_WAIT5041;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$19553\(0 to 30),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$19547_copy_root_in_ram6634352_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5040;
                  end if;
                when Q_WAIT5044 =>
                  \$v5045\ := \$ram_lock\;
                  if \$v5045\(0) = '1' then
                    state_var5921 := Q_WAIT5044;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$19553\(0 to 30),16)));
                    \$ram_write\ <= eclat_resize(\$19547_copy_root_in_ram6634352_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5043;
                  end if;
                when Q_WAIT5047 =>
                  \$v5048\ := \$ram_lock\;
                  if \$v5048\(0) = '1' then
                    state_var5921 := Q_WAIT5047;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19547_copy_root_in_ram6634352_arg\(32 to 47)));
                    \$ram_write\ <= \$19560_hd\; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5046;
                  end if;
                when Q_WAIT5050 =>
                  \$v5051\ := \$ram_lock\;
                  if \$v5051\(0) = '1' then
                    state_var5921 := Q_WAIT5050;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$19553\(0 to 30),16)));
                    state_var5921 := PAUSE_GET5049;
                  end if;
                when Q_WAIT5054 =>
                  \$v5055\ := \$ram_lock\;
                  if \$v5055\(0) = '1' then
                    state_var5921 := Q_WAIT5054;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19553\(0 to 30),16), X"000" & X"1")));
                    state_var5921 := PAUSE_GET5053;
                  end if;
                when Q_WAIT5058 =>
                  \$v5059\ := \$ram_lock\;
                  if \$v5059\(0) = '1' then
                    state_var5921 := Q_WAIT5058;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(\$19547_copy_root_in_ram6634352_arg\(0 to 15)));
                    state_var5921 := PAUSE_GET5057;
                  end if;
                when Q_WAIT5062 =>
                  \$v5063\ := \$ram_lock\;
                  if \$v5063\(0) = '1' then
                    state_var5921 := Q_WAIT5062;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19535_copy_root_in_ram6634354_arg\(0 to 15)));
                    \$ram_write\ <= \$19542\(0 to 31); \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5061;
                  end if;
                when Q_WAIT5065 =>
                  \$v5066\ := \$ram_lock\;
                  if \$v5066\(0) = '1' then
                    state_var5921 := Q_WAIT5065;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$19541\(0 to 30),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$19535_copy_root_in_ram6634354_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5064;
                  end if;
                when Q_WAIT5068 =>
                  \$v5069\ := \$ram_lock\;
                  if \$v5069\(0) = '1' then
                    state_var5921 := Q_WAIT5068;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$19541\(0 to 30),16)));
                    \$ram_write\ <= eclat_resize(\$19535_copy_root_in_ram6634354_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5067;
                  end if;
                when Q_WAIT5071 =>
                  \$v5072\ := \$ram_lock\;
                  if \$v5072\(0) = '1' then
                    state_var5921 := Q_WAIT5071;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19535_copy_root_in_ram6634354_arg\(32 to 47)));
                    \$ram_write\ <= \$19575_hd\; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5070;
                  end if;
                when Q_WAIT5074 =>
                  \$v5075\ := \$ram_lock\;
                  if \$v5075\(0) = '1' then
                    state_var5921 := Q_WAIT5074;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$19541\(0 to 30),16)));
                    state_var5921 := PAUSE_GET5073;
                  end if;
                when Q_WAIT5078 =>
                  \$v5079\ := \$ram_lock\;
                  if \$v5079\(0) = '1' then
                    state_var5921 := Q_WAIT5078;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19541\(0 to 30),16), X"000" & X"1")));
                    state_var5921 := PAUSE_GET5077;
                  end if;
                when Q_WAIT5082 =>
                  \$v5083\ := \$ram_lock\;
                  if \$v5083\(0) = '1' then
                    state_var5921 := Q_WAIT5082;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(\$19535_copy_root_in_ram6634354_arg\(0 to 15)));
                    state_var5921 := PAUSE_GET5081;
                  end if;
                when Q_WAIT5086 =>
                  \$v5087\ := \$global_end_lock\;
                  if \$v5087\(0) = '1' then
                    state_var5921 := Q_WAIT5086;
                  else
                    acquire(\$global_end_lock\);
                    \$global_end_ptr\ <= 0;
                    state_var5921 := PAUSE_GET5085;
                  end if;
                when Q_WAIT5089 =>
                  \$v5090\ := \$ram_lock\;
                  if \$v5090\(0) = '1' then
                    state_var5921 := Q_WAIT5089;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19601_copy_root_in_ram6634352_arg\(0 to 15)));
                    \$ram_write\ <= \$19608\(0 to 31); \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5088;
                  end if;
                when Q_WAIT5092 =>
                  \$v5093\ := \$ram_lock\;
                  if \$v5093\(0) = '1' then
                    state_var5921 := Q_WAIT5092;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$19607\(0 to 30),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$19601_copy_root_in_ram6634352_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5091;
                  end if;
                when Q_WAIT5095 =>
                  \$v5096\ := \$ram_lock\;
                  if \$v5096\(0) = '1' then
                    state_var5921 := Q_WAIT5095;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$19607\(0 to 30),16)));
                    \$ram_write\ <= eclat_resize(\$19601_copy_root_in_ram6634352_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5094;
                  end if;
                when Q_WAIT5098 =>
                  \$v5099\ := \$ram_lock\;
                  if \$v5099\(0) = '1' then
                    state_var5921 := Q_WAIT5098;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19601_copy_root_in_ram6634352_arg\(32 to 47)));
                    \$ram_write\ <= \$19614_hd\; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5097;
                  end if;
                when Q_WAIT5101 =>
                  \$v5102\ := \$ram_lock\;
                  if \$v5102\(0) = '1' then
                    state_var5921 := Q_WAIT5101;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$19607\(0 to 30),16)));
                    state_var5921 := PAUSE_GET5100;
                  end if;
                when Q_WAIT5105 =>
                  \$v5106\ := \$ram_lock\;
                  if \$v5106\(0) = '1' then
                    state_var5921 := Q_WAIT5105;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19607\(0 to 30),16), X"000" & X"1")));
                    state_var5921 := PAUSE_GET5104;
                  end if;
                when Q_WAIT5109 =>
                  \$v5110\ := \$ram_lock\;
                  if \$v5110\(0) = '1' then
                    state_var5921 := Q_WAIT5109;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(\$19601_copy_root_in_ram6634352_arg\(0 to 15)));
                    state_var5921 := PAUSE_GET5108;
                  end if;
                when Q_WAIT5113 =>
                  \$v5114\ := \$ram_lock\;
                  if \$v5114\(0) = '1' then
                    state_var5921 := Q_WAIT5113;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19589_copy_root_in_ram6634353_arg\(0 to 15)));
                    \$ram_write\ <= \$19596\(0 to 31); \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5112;
                  end if;
                when Q_WAIT5116 =>
                  \$v5117\ := \$ram_lock\;
                  if \$v5117\(0) = '1' then
                    state_var5921 := Q_WAIT5116;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$19595\(0 to 30),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$19589_copy_root_in_ram6634353_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5115;
                  end if;
                when Q_WAIT5119 =>
                  \$v5120\ := \$ram_lock\;
                  if \$v5120\(0) = '1' then
                    state_var5921 := Q_WAIT5119;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$19595\(0 to 30),16)));
                    \$ram_write\ <= eclat_resize(\$19589_copy_root_in_ram6634353_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5118;
                  end if;
                when Q_WAIT5122 =>
                  \$v5123\ := \$ram_lock\;
                  if \$v5123\(0) = '1' then
                    state_var5921 := Q_WAIT5122;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19589_copy_root_in_ram6634353_arg\(32 to 47)));
                    \$ram_write\ <= \$19629_hd\; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5121;
                  end if;
                when Q_WAIT5125 =>
                  \$v5126\ := \$ram_lock\;
                  if \$v5126\(0) = '1' then
                    state_var5921 := Q_WAIT5125;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$19595\(0 to 30),16)));
                    state_var5921 := PAUSE_GET5124;
                  end if;
                when Q_WAIT5129 =>
                  \$v5130\ := \$ram_lock\;
                  if \$v5130\(0) = '1' then
                    state_var5921 := Q_WAIT5129;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19595\(0 to 30),16), X"000" & X"1")));
                    state_var5921 := PAUSE_GET5128;
                  end if;
                when Q_WAIT5133 =>
                  \$v5134\ := \$ram_lock\;
                  if \$v5134\(0) = '1' then
                    state_var5921 := Q_WAIT5133;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(\$19589_copy_root_in_ram6634353_arg\(0 to 15)));
                    state_var5921 := PAUSE_GET5132;
                  end if;
                when Q_WAIT5137 =>
                  \$v5138\ := \$ram_lock\;
                  if \$v5138\(0) = '1' then
                    state_var5921 := Q_WAIT5137;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$18792_wait662_arg\(33 to 63),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$19505\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5136;
                  end if;
                when Q_WAIT5140 =>
                  \$v5141\ := \$ram_lock\;
                  if \$v5141\(0) = '1' then
                    state_var5921 := Q_WAIT5140;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18792_wait662_arg\(33 to 63),16)));
                    \$ram_write\ <= eclat_resize(\$19505\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5139;
                  end if;
                when Q_WAIT5143 =>
                  \$v5144\ := \$ram_lock\;
                  if \$v5144\(0) = '1' then
                    state_var5921 := Q_WAIT5143;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19505\(32 to 47)));
                    \$ram_write\ <= \$19644_hd\; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5142;
                  end if;
                when Q_WAIT5146 =>
                  \$v5147\ := \$ram_lock\;
                  if \$v5147\(0) = '1' then
                    state_var5921 := Q_WAIT5146;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18792_wait662_arg\(33 to 63),16)));
                    state_var5921 := PAUSE_GET5145;
                  end if;
                when Q_WAIT5150 =>
                  \$v5151\ := \$ram_lock\;
                  if \$v5151\(0) = '1' then
                    state_var5921 := Q_WAIT5150;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18792_wait662_arg\(33 to 63),16), X"000" & X"1")));
                    state_var5921 := PAUSE_GET5149;
                  end if;
                when Q_WAIT5154 =>
                  \$v5155\ := \$ram_lock\;
                  if \$v5155\(0) = '1' then
                    state_var5921 := Q_WAIT5154;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$18792_wait662_arg\(1 to 31),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$19493\(112 to 127),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5153;
                  end if;
                when Q_WAIT5157 =>
                  \$v5158\ := \$ram_lock\;
                  if \$v5158\(0) = '1' then
                    state_var5921 := Q_WAIT5157;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18792_wait662_arg\(1 to 31),16)));
                    \$ram_write\ <= eclat_resize(\$19493\(112 to 127),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5156;
                  end if;
                when Q_WAIT5160 =>
                  \$v5161\ := \$ram_lock\;
                  if \$v5161\(0) = '1' then
                    state_var5921 := Q_WAIT5160;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19493\(112 to 127)));
                    \$ram_write\ <= \$19659_hd\; \$ram_write_request\ <= '1';
                    state_var5921 := PAUSE_SET5159;
                  end if;
                when Q_WAIT5163 =>
                  \$v5164\ := \$ram_lock\;
                  if \$v5164\(0) = '1' then
                    state_var5921 := Q_WAIT5163;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18792_wait662_arg\(1 to 31),16)));
                    state_var5921 := PAUSE_GET5162;
                  end if;
                when Q_WAIT5167 =>
                  \$v5168\ := \$ram_lock\;
                  if \$v5168\(0) = '1' then
                    state_var5921 := Q_WAIT5167;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18792_wait662_arg\(1 to 31),16), X"000" & X"1")));
                    state_var5921 := PAUSE_GET5166;
                  end if;
                when IDLE4965 =>
                  rdy4964 := eclat_false;
                  \$v5170\ := work.Int.gt(work.Int.add(\$19493\(80 to 95), \$18792_wait662_arg\(81 to 96)), 
                                          work.Int.add(\$19493\(96 to 111), X"1770"));
                  if \$v5170\(0) = '1' then
                    \$19500\ := work.Print.print_newline(clk,eclat_unit);
                    \$19501\ := work.Print.print_newline(clk,eclat_unit);
                    \$19502\ := work.Print.print_string(clk,of_string("[================= GC START ======================]"));
                    \$19503\ := work.Print.print_newline(clk,eclat_unit);
                    \$19504\ := work.Print.print_newline(clk,eclat_unit);
                    \$v5169\ := work.Bool.lnot(eclat_if(work.Bool.lnot(
                                                        ""&\$18792_wait662_arg\(32)) & 
                                               eclat_if(work.Int.le(\$19493\(96 to 111), eclat_resize(\$18792_wait662_arg\(1 to 31),16)) & 
                                               work.Int.lt(eclat_resize(\$18792_wait662_arg\(1 to 31),16), 
                                                           work.Int.add(
                                                           \$19493\(96 to 111), X"1770")) & eclat_false) & eclat_false));
                    if \$v5169\(0) = '1' then
                      \$19505\ := \$18792_wait662_arg\(1 to 32) & \$19493\(112 to 127);
                      \$v5152\ := work.Bool.lnot(eclat_if(work.Bool.lnot(
                                                          ""&\$18792_wait662_arg\(64)) & 
                                                 eclat_if(work.Int.le(
                                                          \$19493\(96 to 111), eclat_resize(\$18792_wait662_arg\(33 to 63),16)) & 
                                                 work.Int.lt(eclat_resize(\$18792_wait662_arg\(33 to 63),16), 
                                                             work.Int.add(
                                                             \$19493\(96 to 111), X"1770")) & eclat_false) & eclat_false));
                      if \$v5152\(0) = '1' then
                        \$19506\ := \$18792_wait662_arg\(33 to 64) & \$19505\(32 to 47);
                        \$19589_copy_root_in_ram6634353_id\ := "000000110000";
                        \$19589_copy_root_in_ram6634353_arg\ := X"0" & X"3e8" & \$18792_wait662_arg\(65 to 80) & \$19506\(32 to 47) & \$19493\(96 to 111) & \$19493\(112 to 127);
                        state_var5921 := \$19589_COPY_ROOT_IN_RAM6634353\;
                      else
                        \$v5151\ := \$ram_lock\;
                        if \$v5151\(0) = '1' then
                          state_var5921 := Q_WAIT5150;
                        else
                          acquire(\$ram_lock\);
                          \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$18792_wait662_arg\(33 to 63),16), X"000" & X"1")));
                          state_var5921 := PAUSE_GET5149;
                        end if;
                      end if;
                    else
                      \$v5168\ := \$ram_lock\;
                      if \$v5168\(0) = '1' then
                        state_var5921 := Q_WAIT5167;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$18792_wait662_arg\(1 to 31),16), X"000" & X"1")));
                        state_var5921 := PAUSE_GET5166;
                      end if;
                    end if;
                  else
                    result4963 := \$18792_wait662_arg\(1 to 32) & \$18792_wait662_arg\(33 to 64) & \$19493\(80 to 95) & 
                    work.Int.add(\$19493\(80 to 95), \$18792_wait662_arg\(81 to 96)) & \$19493\(96 to 111) & \$19493\(112 to 127);
                    rdy4964 := eclat_true;
                    state_var5921 := IDLE4965;
                  end if;
                end case;
                
                if rdy4964(0) = '1' then
                  
                else
                  result4963 := \$19493\(0 to 31) & \$19493\(32 to 63) & \$19493\(64 to 79) & \$19493\(80 to 95) & \$19493\(96 to 111) & \$19493\(112 to 127);
                end if;
                \$19493\ := result4963 & rdy4964;
                \$19492\ := \$19493\;
                \$v4962\ := ""&\$19492\(128);
                if \$v4962\(0) = '1' then
                  \$18792_wait662_result\ := \$19492\(0 to 31) & \$19492\(32 to 63) & \$19492\(64 to 79);
                  \$19485\ := \$18792_wait662_result\;
                  \$19486\ := work.Print.print_string(clk,of_string("size:"));
                  \$19487\ := work.Int.print(clk,eclat_if(work.Int.eq(
                                                          \$18793_make_block579_arg\(88 to 103), X"000" & X"0") & X"000" & X"1" & \$18793_make_block579_arg\(88 to 103)));
                  \$19488\ := work.Print.print_newline(clk,eclat_unit);
                  \$v5174\ := \$ram_lock\;
                  if \$v5174\(0) = '1' then
                    state_var5920 := Q_WAIT5173;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19485\(64 to 79)));
                    \$ram_write\ <= work.Int.lor(work.Int.lsl(eclat_resize(\$18793_make_block579_arg\(80 to 87),31), X"000000" & X"18"), 
                                                 work.Int.lsl(eclat_resize(
                                                              eclat_if(
                                                              work.Int.eq(
                                                              \$18793_make_block579_arg\(88 to 103), X"000" & X"0") & X"000" & X"1" & \$18793_make_block579_arg\(88 to 103)),31), X"0000000" & X"2")) & eclat_true; \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5172;
                  end if;
                else
                  \$18792_wait662_arg\ := eclat_unit & \$18792_wait662_arg\(1 to 32) & \$18792_wait662_arg\(33 to 64) & \$18792_wait662_arg\(65 to 80) & \$18792_wait662_arg\(81 to 96);
                  state_var5920 := \$18792_WAIT662\;
                end if;
              when \$18793_MAKE_BLOCK579\ =>
                \$19481\ := work.Print.print_string(clk,of_string("GC-ALLOC:(size="));
                \$19482\ := work.Int.print(clk,work.Int.add(eclat_if(
                                                            work.Int.eq(
                                                            \$18793_make_block579_arg\(88 to 103), X"000" & X"0") & X"000" & X"1" & \$18793_make_block579_arg\(88 to 103)), X"000" & X"1"));
                \$19483\ := work.Print.print_string(clk,of_string(")"));
                \$19484\ := work.Print.print_newline(clk,eclat_unit);
                \$18792_wait662_id\ := "000000110011";
                \$18792_wait662_arg\ := eclat_unit & \$18793_make_block579_arg\(16 to 47) & \$18793_make_block579_arg\(48 to 79) & \$18793_make_block579_arg\(0 to 15) & 
                work.Int.add(eclat_if(work.Int.eq(\$18793_make_block579_arg\(88 to 103), X"000" & X"0") & X"000" & X"1" & \$18793_make_block579_arg\(88 to 103)), X"000" & X"1");
                state_var5920 := \$18792_WAIT662\;
              when \$18794_APPLY638\ =>
                \$19456\ := work.Print.print_string(clk,of_string("ENV:"));
                \$19457\ := work.Int.print(clk,\$18794_apply638_arg\(110 to 140));
                \$19458\ := work.Print.print_string(clk,of_string("<"));
                \$v5212\ := ""&\$18794_apply638_arg\(141);
                if \$v5212\(0) = '1' then
                  \$19459\ := work.Print.print_string(clk,of_string("int"));
                  \$19460\ := work.Print.print_string(clk,of_string(">"));
                  \$19461\ := work.Print.print_newline(clk,eclat_unit);
                  \$v5211\ := ""&\$18794_apply638_arg\(0);
                  if \$v5211\(0) = '1' then
                    \$v5210\ := \$ram_lock\;
                    if \$v5210\(0) = '1' then
                      state_var5920 := Q_WAIT5209;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(
                                                        \$18794_apply638_arg\(92 to 107), X"000" & X"1")));
                      state_var5920 := PAUSE_GET5208;
                    end if;
                  else
                    \$19462\ := "000"& X"000000" & X"1" & eclat_true & \$18794_apply638_arg\(92 to 107);
                    \$v5207\ := ""&\$18794_apply638_arg\(1);
                    if \$v5207\(0) = '1' then
                      \$v5206\ := \$ram_lock\;
                      if \$v5206\(0) = '1' then
                        state_var5920 := Q_WAIT5205;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(
                                                          \$19462\(32 to 47), X"000" & X"1")));
                        state_var5920 := PAUSE_GET5204;
                      end if;
                    else
                      \$19463\ := "000"& X"000000" & X"1" & eclat_true & \$19462\(32 to 47);
                      \$v5203\ := ""&\$18794_apply638_arg\(2);
                      if \$v5203\(0) = '1' then
                        \$v5202\ := \$ram_lock\;
                        if \$v5202\(0) = '1' then
                          state_var5920 := Q_WAIT5201;
                        else
                          acquire(\$ram_lock\);
                          \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(
                                                            \$19463\(32 to 47), X"000" & X"1")));
                          state_var5920 := PAUSE_GET5200;
                        end if;
                      else
                        \$19464\ := "000"& X"000000" & X"1" & eclat_true & \$19463\(32 to 47);
                        \$v5199\ := ""&\$18794_apply638_arg\(11);
                        if \$v5199\(0) = '1' then
                          \$19465_sp\ := work.Int.add(work.Int.sub(\$19464\(32 to 47), \$18794_apply638_arg\(12 to 27)), \$18794_apply638_arg\(28 to 43));
                          \$v5189\ := ""&\$18794_apply638_arg\(2);
                          if \$v5189\(0) = '1' then
                            \$v5188\ := \$ram_lock\;
                            if \$v5188\(0) = '1' then
                              state_var5920 := Q_WAIT5187;
                            else
                              acquire(\$ram_lock\);
                              \$ram_ptr_write\ <= to_integer(unsigned(\$19465_sp\));
                              \$ram_write\ <= \$19464\(0 to 31); \$ram_write_request\ <= '1';
                              state_var5920 := PAUSE_SET5186;
                            end if;
                          else
                            \$19466_sp\ := \$19465_sp\;
                            \$v5185\ := ""&\$18794_apply638_arg\(1);
                            if \$v5185\(0) = '1' then
                              \$v5184\ := \$ram_lock\;
                              if \$v5184\(0) = '1' then
                                state_var5920 := Q_WAIT5183;
                              else
                                acquire(\$ram_lock\);
                                \$ram_ptr_write\ <= to_integer(unsigned(\$19466_sp\));
                                \$ram_write\ <= \$19463\(0 to 31); \$ram_write_request\ <= '1';
                                state_var5920 := PAUSE_SET5182;
                              end if;
                            else
                              \$19467_sp\ := \$19466_sp\;
                              \$v5181\ := ""&\$18794_apply638_arg\(0);
                              if \$v5181\(0) = '1' then
                                \$v5180\ := \$ram_lock\;
                                if \$v5180\(0) = '1' then
                                  state_var5920 := Q_WAIT5179;
                                else
                                  acquire(\$ram_lock\);
                                  \$ram_ptr_write\ <= to_integer(unsigned(\$19467_sp\));
                                  \$ram_write\ <= \$19462\(0 to 31); \$ram_write_request\ <= '1';
                                  state_var5920 := PAUSE_SET5178;
                                end if;
                              else
                                \$19468_sp\ := \$19467_sp\;
                                \$v5177\ := \$ram_lock\;
                                if \$v5177\(0) = '1' then
                                  state_var5920 := Q_WAIT5176;
                                else
                                  acquire(\$ram_lock\);
                                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                                    work.Int.add(
                                                                    eclat_resize(\$18794_apply638_arg\(60 to 90),16), X"000" & X"0"), X"000" & X"1")));
                                  state_var5920 := PAUSE_GET5175;
                                end if;
                              end if;
                            end if;
                          end if;
                        else
                          \$v5198\ := \$ram_lock\;
                          if \$v5198\(0) = '1' then
                            state_var5920 := Q_WAIT5197;
                          else
                            acquire(\$ram_lock\);
                            \$ram_ptr_write\ <= to_integer(unsigned(\$19464\(32 to 47)));
                            \$ram_write\ <= eclat_resize(\$18794_apply638_arg\(142 to 149),31) & eclat_true; \$ram_write_request\ <= '1';
                            state_var5920 := PAUSE_SET5196;
                          end if;
                        end if;
                      end if;
                    end if;
                  end if;
                else
                  \$19459\ := work.Print.print_string(clk,of_string("ptr"));
                  \$19460\ := work.Print.print_string(clk,of_string(">"));
                  \$19461\ := work.Print.print_newline(clk,eclat_unit);
                  \$v5211\ := ""&\$18794_apply638_arg\(0);
                  if \$v5211\(0) = '1' then
                    \$v5210\ := \$ram_lock\;
                    if \$v5210\(0) = '1' then
                      state_var5920 := Q_WAIT5209;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(
                                                        \$18794_apply638_arg\(92 to 107), X"000" & X"1")));
                      state_var5920 := PAUSE_GET5208;
                    end if;
                  else
                    \$19462\ := "000"& X"000000" & X"1" & eclat_true & \$18794_apply638_arg\(92 to 107);
                    \$v5207\ := ""&\$18794_apply638_arg\(1);
                    if \$v5207\(0) = '1' then
                      \$v5206\ := \$ram_lock\;
                      if \$v5206\(0) = '1' then
                        state_var5920 := Q_WAIT5205;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(
                                                          \$19462\(32 to 47), X"000" & X"1")));
                        state_var5920 := PAUSE_GET5204;
                      end if;
                    else
                      \$19463\ := "000"& X"000000" & X"1" & eclat_true & \$19462\(32 to 47);
                      \$v5203\ := ""&\$18794_apply638_arg\(2);
                      if \$v5203\(0) = '1' then
                        \$v5202\ := \$ram_lock\;
                        if \$v5202\(0) = '1' then
                          state_var5920 := Q_WAIT5201;
                        else
                          acquire(\$ram_lock\);
                          \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(
                                                            \$19463\(32 to 47), X"000" & X"1")));
                          state_var5920 := PAUSE_GET5200;
                        end if;
                      else
                        \$19464\ := "000"& X"000000" & X"1" & eclat_true & \$19463\(32 to 47);
                        \$v5199\ := ""&\$18794_apply638_arg\(11);
                        if \$v5199\(0) = '1' then
                          \$19465_sp\ := work.Int.add(work.Int.sub(\$19464\(32 to 47), \$18794_apply638_arg\(12 to 27)), \$18794_apply638_arg\(28 to 43));
                          \$v5189\ := ""&\$18794_apply638_arg\(2);
                          if \$v5189\(0) = '1' then
                            \$v5188\ := \$ram_lock\;
                            if \$v5188\(0) = '1' then
                              state_var5920 := Q_WAIT5187;
                            else
                              acquire(\$ram_lock\);
                              \$ram_ptr_write\ <= to_integer(unsigned(\$19465_sp\));
                              \$ram_write\ <= \$19464\(0 to 31); \$ram_write_request\ <= '1';
                              state_var5920 := PAUSE_SET5186;
                            end if;
                          else
                            \$19466_sp\ := \$19465_sp\;
                            \$v5185\ := ""&\$18794_apply638_arg\(1);
                            if \$v5185\(0) = '1' then
                              \$v5184\ := \$ram_lock\;
                              if \$v5184\(0) = '1' then
                                state_var5920 := Q_WAIT5183;
                              else
                                acquire(\$ram_lock\);
                                \$ram_ptr_write\ <= to_integer(unsigned(\$19466_sp\));
                                \$ram_write\ <= \$19463\(0 to 31); \$ram_write_request\ <= '1';
                                state_var5920 := PAUSE_SET5182;
                              end if;
                            else
                              \$19467_sp\ := \$19466_sp\;
                              \$v5181\ := ""&\$18794_apply638_arg\(0);
                              if \$v5181\(0) = '1' then
                                \$v5180\ := \$ram_lock\;
                                if \$v5180\(0) = '1' then
                                  state_var5920 := Q_WAIT5179;
                                else
                                  acquire(\$ram_lock\);
                                  \$ram_ptr_write\ <= to_integer(unsigned(\$19467_sp\));
                                  \$ram_write\ <= \$19462\(0 to 31); \$ram_write_request\ <= '1';
                                  state_var5920 := PAUSE_SET5178;
                                end if;
                              else
                                \$19468_sp\ := \$19467_sp\;
                                \$v5177\ := \$ram_lock\;
                                if \$v5177\(0) = '1' then
                                  state_var5920 := Q_WAIT5176;
                                else
                                  acquire(\$ram_lock\);
                                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                                    work.Int.add(
                                                                    eclat_resize(\$18794_apply638_arg\(60 to 90),16), X"000" & X"0"), X"000" & X"1")));
                                  state_var5920 := PAUSE_GET5175;
                                end if;
                              end if;
                            end if;
                          end if;
                        else
                          \$v5198\ := \$ram_lock\;
                          if \$v5198\(0) = '1' then
                            state_var5920 := Q_WAIT5197;
                          else
                            acquire(\$ram_lock\);
                            \$ram_ptr_write\ <= to_integer(unsigned(\$19464\(32 to 47)));
                            \$ram_write\ <= eclat_resize(\$18794_apply638_arg\(142 to 149),31) & eclat_true; \$ram_write_request\ <= '1';
                            state_var5920 := PAUSE_SET5196;
                          end if;
                        end if;
                      end if;
                    end if;
                  end if;
                end if;
              when \$18795_OFFSETCLOSURE_N639\ =>
                \$18795_offsetclosure_n639_result\ := \$18795_offsetclosure_n639_arg\(0 to 15) & eclat_resize(
                work.Int.add(eclat_resize(\$18795_offsetclosure_n639_arg\(106 to 136),16), \$18795_offsetclosure_n639_arg\(32 to 47)),31) & eclat_false & \$18795_offsetclosure_n639_arg\(16 to 31) & \$18795_offsetclosure_n639_arg\(48 to 103) & \$18795_offsetclosure_n639_arg\(104 to 105);
                result4928 := \$18795_offsetclosure_n639_result\;
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when \$18796_MAKE_BLOCK_N646\ =>
                \$18793_make_block579_id\ := "000000110100";
                \$18793_make_block579_arg\ := \$18796_make_block_n646_arg\(16 to 31) & \$18796_make_block_n646_arg\(82 to 113) & \$18796_make_block_n646_arg\(116 to 147) & eclat_resize(\$18796_make_block_n646_arg\(35 to 65),8) & \$18796_make_block_n646_arg\(66 to 81);
                state_var5920 := \$18793_MAKE_BLOCK579\;
              when \$18797_BRANCH_IF648\ =>
                \$v5234\ := eclat_if(""&\$18797_branch_if648_arg\(0) & 
                            work.Bool.lnot(work.Int.neq(\$18797_branch_if648_arg\(17 to 47), "000"& X"000000" & X"0")) & 
                            work.Int.neq(\$18797_branch_if648_arg\(17 to 47), "000"& X"000000" & X"0"));
                if \$v5234\(0) = '1' then
                  \$v5233\ := \$code_lock\;
                  if \$v5233\(0) = '1' then
                    state_var5920 := Q_WAIT5232;
                  else
                    acquire(\$code_lock\);
                    \$code_ptr\ <= to_integer(unsigned(work.Int.add(\$18797_branch_if648_arg\(1 to 16), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5231;
                  end if;
                else
                  \$18797_branch_if648_result\ := work.Int.add(\$18797_branch_if648_arg\(1 to 16), X"000" & X"2") & \$18797_branch_if648_arg\(17 to 48) & \$18797_branch_if648_arg\(49 to 64) & \$18797_branch_if648_arg\(65 to 120) & \$18797_branch_if648_arg\(121 to 122);
                  result4928 := \$18797_branch_if648_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                end if;
              when \$18798_W652\ =>
                \$v5241\ := work.Int.gt(\$18798_w652_arg\(0 to 15), \$18798_w652_arg\(32 to 47));
                if \$v5241\(0) = '1' then
                  \$18798_w652_result\ := eclat_unit;
                  \$19341\ := \$18798_w652_result\;
                  \$v5828\ := \$ram_lock\;
                  if \$v5828\(0) = '1' then
                    state_var5920 := Q_WAIT5827;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$18788\(16 to 46),16), X"000" & X"0"), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5826;
                  end if;
                else
                  \$v5240\ := \$ram_lock\;
                  if \$v5240\(0) = '1' then
                    state_var5920 := Q_WAIT5239;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18798_w652_arg\(16 to 31), \$18798_w652_arg\(0 to 15))));
                    state_var5920 := PAUSE_GET5238;
                  end if;
                end if;
              when \$18799_W1656\ =>
                \$v5251\ := work.Int.ge(\$18799_w1656_arg\(0 to 15), \$18799_w1656_arg\(32 to 47));
                if \$v5251\(0) = '1' then
                  \$18799_w1656_result\ := eclat_unit;
                  \$19413\ := \$18799_w1656_result\;
                  \$v5880\ := \$ram_lock\;
                  if \$v5880\(0) = '1' then
                    state_var5920 := Q_WAIT5879;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19412_sp\));
                    \$ram_write\ <= \$19410\(64 to 95); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5878;
                  end if;
                else
                  \$v5250\ := \$ram_lock\;
                  if \$v5250\(0) = '1' then
                    state_var5920 := Q_WAIT5249;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            work.Int.add(
                                                            eclat_resize(\$18799_w1656_arg\(48 to 78),16), 
                                                            work.Int.sub(
                                                            work.Int.mul(
                                                            X"000" & X"2", \$18799_w1656_arg\(0 to 15)), X"000" & X"1")), X"000" & X"1")));
                    \$ram_write\ <= work.Int.lor(work.Int.lsl(eclat_resize("11111001",31), X"000000" & X"18"), 
                                                 work.Int.lsl(eclat_resize(
                                                              work.Int.mul(
                                                              X"000" & X"2", \$18799_w1656_arg\(0 to 15)),31), X"0000000" & X"2")) & eclat_true; \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5248;
                  end if;
                end if;
              when \$18856_LOOP_PUSH6494360\ =>
                \$v5369\ := work.Int.ge(\$18856_loop_push6494360_arg\(16 to 23), 
                                        work.Int.sub(\$18856_loop_push6494360_arg\(56 to 63), "00000010"));
                if \$v5369\(0) = '1' then
                  \$18856_loop_push6494360_result\ := \$18856_loop_push6494360_arg\(0 to 15);
                  \$18854_sp\ := \$18856_loop_push6494360_result\;
                  \$v5362\ := \$ram_lock\;
                  if \$v5362\(0) = '1' then
                    state_var5920 := Q_WAIT5361;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$18788\(64 to 94),16), X"000" & X"1"), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5360;
                  end if;
                else
                  \$v5368\ := \$ram_lock\;
                  if \$v5368\(0) = '1' then
                    state_var5920 := Q_WAIT5367;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$18856_loop_push6494360_arg\(24 to 54),16), eclat_resize(
                                                                   work.Int.add(
                                                                   \$18856_loop_push6494360_arg\(16 to 23), "00000010"),16)), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5366;
                  end if;
                end if;
              when \$18901_BINOP_INT6434361\ =>
                \$v5490\ := \$ram_lock\;
                if \$v5490\(0) = '1' then
                  state_var5920 := Q_WAIT5489;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18901_binop_int6434361_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5488;
                end if;
              when \$18907_MODULO6684356\ =>
                \$v5482\ := work.Int.lt(\$18907_modulo6684356_arg\(0 to 30), \$18907_modulo6684356_arg\(31 to 61));
                if \$v5482\(0) = '1' then
                  \$18907_modulo6684356_result\ := \$18907_modulo6684356_arg\(0 to 30);
                  \$18906_r\ := \$18907_modulo6684356_result\;
                  \$18905_res\ := eclat_if(work.Int.lt(\$18901_binop_int6434361_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$18906_r\) & \$18906_r\);
                  \$18901_binop_int6434361_result\ := work.Int.add(\$18901_binop_int6434361_arg\(32 to 47), X"000" & X"1") & \$18905_res\ & eclat_true & 
                  work.Int.sub(\$18901_binop_int6434361_arg\(80 to 95), X"000" & X"1") & \$18901_binop_int6434361_arg\(96 to 151) & \$18901_binop_int6434361_arg\(152 to 153);
                  result4928 := \$18901_binop_int6434361_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$18910_modulo6684349_id\ := "000001000011";
                  \$18910_modulo6684349_arg\ := work.Int.sub(\$18907_modulo6684356_arg\(0 to 30), \$18907_modulo6684356_arg\(31 to 61)) & \$18907_modulo6684356_arg\(31 to 61);
                  state_var5920 := \$18910_MODULO6684349\;
                end if;
              when \$18910_MODULO6684349\ =>
                \$v5481\ := work.Int.lt(\$18910_modulo6684349_arg\(0 to 30), \$18910_modulo6684349_arg\(31 to 61));
                if \$v5481\(0) = '1' then
                  \$18910_modulo6684349_result\ := \$18910_modulo6684349_arg\(0 to 30);
                  \$18907_modulo6684356_result\ := \$18910_modulo6684349_result\;
                  \$18906_r\ := \$18907_modulo6684356_result\;
                  \$18905_res\ := eclat_if(work.Int.lt(\$18901_binop_int6434361_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$18906_r\) & \$18906_r\);
                  \$18901_binop_int6434361_result\ := work.Int.add(\$18901_binop_int6434361_arg\(32 to 47), X"000" & X"1") & \$18905_res\ & eclat_true & 
                  work.Int.sub(\$18901_binop_int6434361_arg\(80 to 95), X"000" & X"1") & \$18901_binop_int6434361_arg\(96 to 151) & \$18901_binop_int6434361_arg\(152 to 153);
                  result4928 := \$18901_binop_int6434361_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$18910_modulo6684349_arg\ := work.Int.sub(\$18910_modulo6684349_arg\(0 to 30), \$18910_modulo6684349_arg\(31 to 61)) & \$18910_modulo6684349_arg\(31 to 61);
                  state_var5920 := \$18910_MODULO6684349\;
                end if;
              when \$18914_MODULO6684357\ =>
                \$v5485\ := work.Int.lt(\$18914_modulo6684357_arg\(0 to 30), \$18914_modulo6684357_arg\(31 to 61));
                if \$v5485\(0) = '1' then
                  \$18914_modulo6684357_result\ := \$18914_modulo6684357_arg\(0 to 30);
                  \$18913_r\ := \$18914_modulo6684357_result\;
                  \$18905_res\ := eclat_if(work.Int.lt(\$18901_binop_int6434361_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$18913_r\) & \$18913_r\);
                  \$18901_binop_int6434361_result\ := work.Int.add(\$18901_binop_int6434361_arg\(32 to 47), X"000" & X"1") & \$18905_res\ & eclat_true & 
                  work.Int.sub(\$18901_binop_int6434361_arg\(80 to 95), X"000" & X"1") & \$18901_binop_int6434361_arg\(96 to 151) & \$18901_binop_int6434361_arg\(152 to 153);
                  result4928 := \$18901_binop_int6434361_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$18917_modulo6684349_id\ := "000001000101";
                  \$18917_modulo6684349_arg\ := work.Int.sub(\$18914_modulo6684357_arg\(0 to 30), \$18914_modulo6684357_arg\(31 to 61)) & \$18914_modulo6684357_arg\(31 to 61);
                  state_var5920 := \$18917_MODULO6684349\;
                end if;
              when \$18917_MODULO6684349\ =>
                \$v5484\ := work.Int.lt(\$18917_modulo6684349_arg\(0 to 30), \$18917_modulo6684349_arg\(31 to 61));
                if \$v5484\(0) = '1' then
                  \$18917_modulo6684349_result\ := \$18917_modulo6684349_arg\(0 to 30);
                  \$18914_modulo6684357_result\ := \$18917_modulo6684349_result\;
                  \$18913_r\ := \$18914_modulo6684357_result\;
                  \$18905_res\ := eclat_if(work.Int.lt(\$18901_binop_int6434361_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$18913_r\) & \$18913_r\);
                  \$18901_binop_int6434361_result\ := work.Int.add(\$18901_binop_int6434361_arg\(32 to 47), X"000" & X"1") & \$18905_res\ & eclat_true & 
                  work.Int.sub(\$18901_binop_int6434361_arg\(80 to 95), X"000" & X"1") & \$18901_binop_int6434361_arg\(96 to 151) & \$18901_binop_int6434361_arg\(152 to 153);
                  result4928 := \$18901_binop_int6434361_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$18917_modulo6684349_arg\ := work.Int.sub(\$18917_modulo6684349_arg\(0 to 30), \$18917_modulo6684349_arg\(31 to 61)) & \$18917_modulo6684349_arg\(31 to 61);
                  state_var5920 := \$18917_MODULO6684349\;
                end if;
              when \$18920_BINOP_INT6434362\ =>
                \$v5500\ := \$ram_lock\;
                if \$v5500\(0) = '1' then
                  state_var5920 := Q_WAIT5499;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18920_binop_int6434362_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5498;
                end if;
              when \$18926_MODULO6684356\ =>
                \$v5492\ := work.Int.lt(\$18926_modulo6684356_arg\(0 to 30), \$18926_modulo6684356_arg\(31 to 61));
                if \$v5492\(0) = '1' then
                  \$18926_modulo6684356_result\ := \$18926_modulo6684356_arg\(0 to 30);
                  \$18925_r\ := \$18926_modulo6684356_result\;
                  \$18924_res\ := eclat_if(work.Int.lt(\$18920_binop_int6434362_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$18925_r\) & \$18925_r\);
                  \$18920_binop_int6434362_result\ := work.Int.add(\$18920_binop_int6434362_arg\(32 to 47), X"000" & X"1") & \$18924_res\ & eclat_true & 
                  work.Int.sub(\$18920_binop_int6434362_arg\(80 to 95), X"000" & X"1") & \$18920_binop_int6434362_arg\(96 to 151) & \$18920_binop_int6434362_arg\(152 to 153);
                  result4928 := \$18920_binop_int6434362_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$18929_modulo6684349_id\ := "000001001000";
                  \$18929_modulo6684349_arg\ := work.Int.sub(\$18926_modulo6684356_arg\(0 to 30), \$18926_modulo6684356_arg\(31 to 61)) & \$18926_modulo6684356_arg\(31 to 61);
                  state_var5920 := \$18929_MODULO6684349\;
                end if;
              when \$18929_MODULO6684349\ =>
                \$v5491\ := work.Int.lt(\$18929_modulo6684349_arg\(0 to 30), \$18929_modulo6684349_arg\(31 to 61));
                if \$v5491\(0) = '1' then
                  \$18929_modulo6684349_result\ := \$18929_modulo6684349_arg\(0 to 30);
                  \$18926_modulo6684356_result\ := \$18929_modulo6684349_result\;
                  \$18925_r\ := \$18926_modulo6684356_result\;
                  \$18924_res\ := eclat_if(work.Int.lt(\$18920_binop_int6434362_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$18925_r\) & \$18925_r\);
                  \$18920_binop_int6434362_result\ := work.Int.add(\$18920_binop_int6434362_arg\(32 to 47), X"000" & X"1") & \$18924_res\ & eclat_true & 
                  work.Int.sub(\$18920_binop_int6434362_arg\(80 to 95), X"000" & X"1") & \$18920_binop_int6434362_arg\(96 to 151) & \$18920_binop_int6434362_arg\(152 to 153);
                  result4928 := \$18920_binop_int6434362_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$18929_modulo6684349_arg\ := work.Int.sub(\$18929_modulo6684349_arg\(0 to 30), \$18929_modulo6684349_arg\(31 to 61)) & \$18929_modulo6684349_arg\(31 to 61);
                  state_var5920 := \$18929_MODULO6684349\;
                end if;
              when \$18933_MODULO6684357\ =>
                \$v5495\ := work.Int.lt(\$18933_modulo6684357_arg\(0 to 30), \$18933_modulo6684357_arg\(31 to 61));
                if \$v5495\(0) = '1' then
                  \$18933_modulo6684357_result\ := \$18933_modulo6684357_arg\(0 to 30);
                  \$18932_r\ := \$18933_modulo6684357_result\;
                  \$18924_res\ := eclat_if(work.Int.lt(\$18920_binop_int6434362_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$18932_r\) & \$18932_r\);
                  \$18920_binop_int6434362_result\ := work.Int.add(\$18920_binop_int6434362_arg\(32 to 47), X"000" & X"1") & \$18924_res\ & eclat_true & 
                  work.Int.sub(\$18920_binop_int6434362_arg\(80 to 95), X"000" & X"1") & \$18920_binop_int6434362_arg\(96 to 151) & \$18920_binop_int6434362_arg\(152 to 153);
                  result4928 := \$18920_binop_int6434362_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$18936_modulo6684349_id\ := "000001001010";
                  \$18936_modulo6684349_arg\ := work.Int.sub(\$18933_modulo6684357_arg\(0 to 30), \$18933_modulo6684357_arg\(31 to 61)) & \$18933_modulo6684357_arg\(31 to 61);
                  state_var5920 := \$18936_MODULO6684349\;
                end if;
              when \$18936_MODULO6684349\ =>
                \$v5494\ := work.Int.lt(\$18936_modulo6684349_arg\(0 to 30), \$18936_modulo6684349_arg\(31 to 61));
                if \$v5494\(0) = '1' then
                  \$18936_modulo6684349_result\ := \$18936_modulo6684349_arg\(0 to 30);
                  \$18933_modulo6684357_result\ := \$18936_modulo6684349_result\;
                  \$18932_r\ := \$18933_modulo6684357_result\;
                  \$18924_res\ := eclat_if(work.Int.lt(\$18920_binop_int6434362_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$18932_r\) & \$18932_r\);
                  \$18920_binop_int6434362_result\ := work.Int.add(\$18920_binop_int6434362_arg\(32 to 47), X"000" & X"1") & \$18924_res\ & eclat_true & 
                  work.Int.sub(\$18920_binop_int6434362_arg\(80 to 95), X"000" & X"1") & \$18920_binop_int6434362_arg\(96 to 151) & \$18920_binop_int6434362_arg\(152 to 153);
                  result4928 := \$18920_binop_int6434362_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$18936_modulo6684349_arg\ := work.Int.sub(\$18936_modulo6684349_arg\(0 to 30), \$18936_modulo6684349_arg\(31 to 61)) & \$18936_modulo6684349_arg\(31 to 61);
                  state_var5920 := \$18936_MODULO6684349\;
                end if;
              when \$18939_BINOP_INT6434363\ =>
                \$v5510\ := \$ram_lock\;
                if \$v5510\(0) = '1' then
                  state_var5920 := Q_WAIT5509;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18939_binop_int6434363_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5508;
                end if;
              when \$18945_MODULO6684356\ =>
                \$v5502\ := work.Int.lt(\$18945_modulo6684356_arg\(0 to 30), \$18945_modulo6684356_arg\(31 to 61));
                if \$v5502\(0) = '1' then
                  \$18945_modulo6684356_result\ := \$18945_modulo6684356_arg\(0 to 30);
                  \$18944_r\ := \$18945_modulo6684356_result\;
                  \$18943_res\ := eclat_if(work.Int.lt(\$18939_binop_int6434363_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$18944_r\) & \$18944_r\);
                  \$18939_binop_int6434363_result\ := work.Int.add(\$18939_binop_int6434363_arg\(32 to 47), X"000" & X"1") & \$18943_res\ & eclat_true & 
                  work.Int.sub(\$18939_binop_int6434363_arg\(80 to 95), X"000" & X"1") & \$18939_binop_int6434363_arg\(96 to 151) & \$18939_binop_int6434363_arg\(152 to 153);
                  result4928 := \$18939_binop_int6434363_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$18948_modulo6684349_id\ := "000001001101";
                  \$18948_modulo6684349_arg\ := work.Int.sub(\$18945_modulo6684356_arg\(0 to 30), \$18945_modulo6684356_arg\(31 to 61)) & \$18945_modulo6684356_arg\(31 to 61);
                  state_var5920 := \$18948_MODULO6684349\;
                end if;
              when \$18948_MODULO6684349\ =>
                \$v5501\ := work.Int.lt(\$18948_modulo6684349_arg\(0 to 30), \$18948_modulo6684349_arg\(31 to 61));
                if \$v5501\(0) = '1' then
                  \$18948_modulo6684349_result\ := \$18948_modulo6684349_arg\(0 to 30);
                  \$18945_modulo6684356_result\ := \$18948_modulo6684349_result\;
                  \$18944_r\ := \$18945_modulo6684356_result\;
                  \$18943_res\ := eclat_if(work.Int.lt(\$18939_binop_int6434363_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$18944_r\) & \$18944_r\);
                  \$18939_binop_int6434363_result\ := work.Int.add(\$18939_binop_int6434363_arg\(32 to 47), X"000" & X"1") & \$18943_res\ & eclat_true & 
                  work.Int.sub(\$18939_binop_int6434363_arg\(80 to 95), X"000" & X"1") & \$18939_binop_int6434363_arg\(96 to 151) & \$18939_binop_int6434363_arg\(152 to 153);
                  result4928 := \$18939_binop_int6434363_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$18948_modulo6684349_arg\ := work.Int.sub(\$18948_modulo6684349_arg\(0 to 30), \$18948_modulo6684349_arg\(31 to 61)) & \$18948_modulo6684349_arg\(31 to 61);
                  state_var5920 := \$18948_MODULO6684349\;
                end if;
              when \$18952_MODULO6684357\ =>
                \$v5505\ := work.Int.lt(\$18952_modulo6684357_arg\(0 to 30), \$18952_modulo6684357_arg\(31 to 61));
                if \$v5505\(0) = '1' then
                  \$18952_modulo6684357_result\ := \$18952_modulo6684357_arg\(0 to 30);
                  \$18951_r\ := \$18952_modulo6684357_result\;
                  \$18943_res\ := eclat_if(work.Int.lt(\$18939_binop_int6434363_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$18951_r\) & \$18951_r\);
                  \$18939_binop_int6434363_result\ := work.Int.add(\$18939_binop_int6434363_arg\(32 to 47), X"000" & X"1") & \$18943_res\ & eclat_true & 
                  work.Int.sub(\$18939_binop_int6434363_arg\(80 to 95), X"000" & X"1") & \$18939_binop_int6434363_arg\(96 to 151) & \$18939_binop_int6434363_arg\(152 to 153);
                  result4928 := \$18939_binop_int6434363_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$18955_modulo6684349_id\ := "000001001111";
                  \$18955_modulo6684349_arg\ := work.Int.sub(\$18952_modulo6684357_arg\(0 to 30), \$18952_modulo6684357_arg\(31 to 61)) & \$18952_modulo6684357_arg\(31 to 61);
                  state_var5920 := \$18955_MODULO6684349\;
                end if;
              when \$18955_MODULO6684349\ =>
                \$v5504\ := work.Int.lt(\$18955_modulo6684349_arg\(0 to 30), \$18955_modulo6684349_arg\(31 to 61));
                if \$v5504\(0) = '1' then
                  \$18955_modulo6684349_result\ := \$18955_modulo6684349_arg\(0 to 30);
                  \$18952_modulo6684357_result\ := \$18955_modulo6684349_result\;
                  \$18951_r\ := \$18952_modulo6684357_result\;
                  \$18943_res\ := eclat_if(work.Int.lt(\$18939_binop_int6434363_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$18951_r\) & \$18951_r\);
                  \$18939_binop_int6434363_result\ := work.Int.add(\$18939_binop_int6434363_arg\(32 to 47), X"000" & X"1") & \$18943_res\ & eclat_true & 
                  work.Int.sub(\$18939_binop_int6434363_arg\(80 to 95), X"000" & X"1") & \$18939_binop_int6434363_arg\(96 to 151) & \$18939_binop_int6434363_arg\(152 to 153);
                  result4928 := \$18939_binop_int6434363_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$18955_modulo6684349_arg\ := work.Int.sub(\$18955_modulo6684349_arg\(0 to 30), \$18955_modulo6684349_arg\(31 to 61)) & \$18955_modulo6684349_arg\(31 to 61);
                  state_var5920 := \$18955_MODULO6684349\;
                end if;
              when \$18958_BINOP_INT6434364\ =>
                \$v5520\ := \$ram_lock\;
                if \$v5520\(0) = '1' then
                  state_var5920 := Q_WAIT5519;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18958_binop_int6434364_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5518;
                end if;
              when \$18964_MODULO6684356\ =>
                \$v5512\ := work.Int.lt(\$18964_modulo6684356_arg\(0 to 30), \$18964_modulo6684356_arg\(31 to 61));
                if \$v5512\(0) = '1' then
                  \$18964_modulo6684356_result\ := \$18964_modulo6684356_arg\(0 to 30);
                  \$18963_r\ := \$18964_modulo6684356_result\;
                  \$18962_res\ := eclat_if(work.Int.lt(\$18958_binop_int6434364_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$18963_r\) & \$18963_r\);
                  \$18958_binop_int6434364_result\ := work.Int.add(\$18958_binop_int6434364_arg\(32 to 47), X"000" & X"1") & \$18962_res\ & eclat_true & 
                  work.Int.sub(\$18958_binop_int6434364_arg\(80 to 95), X"000" & X"1") & \$18958_binop_int6434364_arg\(96 to 151) & \$18958_binop_int6434364_arg\(152 to 153);
                  result4928 := \$18958_binop_int6434364_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$18967_modulo6684349_id\ := "000001010010";
                  \$18967_modulo6684349_arg\ := work.Int.sub(\$18964_modulo6684356_arg\(0 to 30), \$18964_modulo6684356_arg\(31 to 61)) & \$18964_modulo6684356_arg\(31 to 61);
                  state_var5920 := \$18967_MODULO6684349\;
                end if;
              when \$18967_MODULO6684349\ =>
                \$v5511\ := work.Int.lt(\$18967_modulo6684349_arg\(0 to 30), \$18967_modulo6684349_arg\(31 to 61));
                if \$v5511\(0) = '1' then
                  \$18967_modulo6684349_result\ := \$18967_modulo6684349_arg\(0 to 30);
                  \$18964_modulo6684356_result\ := \$18967_modulo6684349_result\;
                  \$18963_r\ := \$18964_modulo6684356_result\;
                  \$18962_res\ := eclat_if(work.Int.lt(\$18958_binop_int6434364_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$18963_r\) & \$18963_r\);
                  \$18958_binop_int6434364_result\ := work.Int.add(\$18958_binop_int6434364_arg\(32 to 47), X"000" & X"1") & \$18962_res\ & eclat_true & 
                  work.Int.sub(\$18958_binop_int6434364_arg\(80 to 95), X"000" & X"1") & \$18958_binop_int6434364_arg\(96 to 151) & \$18958_binop_int6434364_arg\(152 to 153);
                  result4928 := \$18958_binop_int6434364_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$18967_modulo6684349_arg\ := work.Int.sub(\$18967_modulo6684349_arg\(0 to 30), \$18967_modulo6684349_arg\(31 to 61)) & \$18967_modulo6684349_arg\(31 to 61);
                  state_var5920 := \$18967_MODULO6684349\;
                end if;
              when \$18971_MODULO6684357\ =>
                \$v5515\ := work.Int.lt(\$18971_modulo6684357_arg\(0 to 30), \$18971_modulo6684357_arg\(31 to 61));
                if \$v5515\(0) = '1' then
                  \$18971_modulo6684357_result\ := \$18971_modulo6684357_arg\(0 to 30);
                  \$18970_r\ := \$18971_modulo6684357_result\;
                  \$18962_res\ := eclat_if(work.Int.lt(\$18958_binop_int6434364_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$18970_r\) & \$18970_r\);
                  \$18958_binop_int6434364_result\ := work.Int.add(\$18958_binop_int6434364_arg\(32 to 47), X"000" & X"1") & \$18962_res\ & eclat_true & 
                  work.Int.sub(\$18958_binop_int6434364_arg\(80 to 95), X"000" & X"1") & \$18958_binop_int6434364_arg\(96 to 151) & \$18958_binop_int6434364_arg\(152 to 153);
                  result4928 := \$18958_binop_int6434364_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$18974_modulo6684349_id\ := "000001010100";
                  \$18974_modulo6684349_arg\ := work.Int.sub(\$18971_modulo6684357_arg\(0 to 30), \$18971_modulo6684357_arg\(31 to 61)) & \$18971_modulo6684357_arg\(31 to 61);
                  state_var5920 := \$18974_MODULO6684349\;
                end if;
              when \$18974_MODULO6684349\ =>
                \$v5514\ := work.Int.lt(\$18974_modulo6684349_arg\(0 to 30), \$18974_modulo6684349_arg\(31 to 61));
                if \$v5514\(0) = '1' then
                  \$18974_modulo6684349_result\ := \$18974_modulo6684349_arg\(0 to 30);
                  \$18971_modulo6684357_result\ := \$18974_modulo6684349_result\;
                  \$18970_r\ := \$18971_modulo6684357_result\;
                  \$18962_res\ := eclat_if(work.Int.lt(\$18958_binop_int6434364_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$18970_r\) & \$18970_r\);
                  \$18958_binop_int6434364_result\ := work.Int.add(\$18958_binop_int6434364_arg\(32 to 47), X"000" & X"1") & \$18962_res\ & eclat_true & 
                  work.Int.sub(\$18958_binop_int6434364_arg\(80 to 95), X"000" & X"1") & \$18958_binop_int6434364_arg\(96 to 151) & \$18958_binop_int6434364_arg\(152 to 153);
                  result4928 := \$18958_binop_int6434364_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$18974_modulo6684349_arg\ := work.Int.sub(\$18974_modulo6684349_arg\(0 to 30), \$18974_modulo6684349_arg\(31 to 61)) & \$18974_modulo6684349_arg\(31 to 61);
                  state_var5920 := \$18974_MODULO6684349\;
                end if;
              when \$18977_BINOP_INT6434365\ =>
                \$v5530\ := \$ram_lock\;
                if \$v5530\(0) = '1' then
                  state_var5920 := Q_WAIT5529;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18977_binop_int6434365_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5528;
                end if;
              when \$18983_MODULO6684356\ =>
                \$v5522\ := work.Int.lt(\$18983_modulo6684356_arg\(0 to 30), \$18983_modulo6684356_arg\(31 to 61));
                if \$v5522\(0) = '1' then
                  \$18983_modulo6684356_result\ := \$18983_modulo6684356_arg\(0 to 30);
                  \$18982_r\ := \$18983_modulo6684356_result\;
                  \$18981_res\ := eclat_if(work.Int.lt(\$18977_binop_int6434365_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$18982_r\) & \$18982_r\);
                  \$18977_binop_int6434365_result\ := work.Int.add(\$18977_binop_int6434365_arg\(32 to 47), X"000" & X"1") & \$18981_res\ & eclat_true & 
                  work.Int.sub(\$18977_binop_int6434365_arg\(80 to 95), X"000" & X"1") & \$18977_binop_int6434365_arg\(96 to 151) & \$18977_binop_int6434365_arg\(152 to 153);
                  result4928 := \$18977_binop_int6434365_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$18986_modulo6684349_id\ := "000001010111";
                  \$18986_modulo6684349_arg\ := work.Int.sub(\$18983_modulo6684356_arg\(0 to 30), \$18983_modulo6684356_arg\(31 to 61)) & \$18983_modulo6684356_arg\(31 to 61);
                  state_var5920 := \$18986_MODULO6684349\;
                end if;
              when \$18986_MODULO6684349\ =>
                \$v5521\ := work.Int.lt(\$18986_modulo6684349_arg\(0 to 30), \$18986_modulo6684349_arg\(31 to 61));
                if \$v5521\(0) = '1' then
                  \$18986_modulo6684349_result\ := \$18986_modulo6684349_arg\(0 to 30);
                  \$18983_modulo6684356_result\ := \$18986_modulo6684349_result\;
                  \$18982_r\ := \$18983_modulo6684356_result\;
                  \$18981_res\ := eclat_if(work.Int.lt(\$18977_binop_int6434365_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$18982_r\) & \$18982_r\);
                  \$18977_binop_int6434365_result\ := work.Int.add(\$18977_binop_int6434365_arg\(32 to 47), X"000" & X"1") & \$18981_res\ & eclat_true & 
                  work.Int.sub(\$18977_binop_int6434365_arg\(80 to 95), X"000" & X"1") & \$18977_binop_int6434365_arg\(96 to 151) & \$18977_binop_int6434365_arg\(152 to 153);
                  result4928 := \$18977_binop_int6434365_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$18986_modulo6684349_arg\ := work.Int.sub(\$18986_modulo6684349_arg\(0 to 30), \$18986_modulo6684349_arg\(31 to 61)) & \$18986_modulo6684349_arg\(31 to 61);
                  state_var5920 := \$18986_MODULO6684349\;
                end if;
              when \$18990_MODULO6684357\ =>
                \$v5525\ := work.Int.lt(\$18990_modulo6684357_arg\(0 to 30), \$18990_modulo6684357_arg\(31 to 61));
                if \$v5525\(0) = '1' then
                  \$18990_modulo6684357_result\ := \$18990_modulo6684357_arg\(0 to 30);
                  \$18989_r\ := \$18990_modulo6684357_result\;
                  \$18981_res\ := eclat_if(work.Int.lt(\$18977_binop_int6434365_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$18989_r\) & \$18989_r\);
                  \$18977_binop_int6434365_result\ := work.Int.add(\$18977_binop_int6434365_arg\(32 to 47), X"000" & X"1") & \$18981_res\ & eclat_true & 
                  work.Int.sub(\$18977_binop_int6434365_arg\(80 to 95), X"000" & X"1") & \$18977_binop_int6434365_arg\(96 to 151) & \$18977_binop_int6434365_arg\(152 to 153);
                  result4928 := \$18977_binop_int6434365_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$18993_modulo6684349_id\ := "000001011001";
                  \$18993_modulo6684349_arg\ := work.Int.sub(\$18990_modulo6684357_arg\(0 to 30), \$18990_modulo6684357_arg\(31 to 61)) & \$18990_modulo6684357_arg\(31 to 61);
                  state_var5920 := \$18993_MODULO6684349\;
                end if;
              when \$18993_MODULO6684349\ =>
                \$v5524\ := work.Int.lt(\$18993_modulo6684349_arg\(0 to 30), \$18993_modulo6684349_arg\(31 to 61));
                if \$v5524\(0) = '1' then
                  \$18993_modulo6684349_result\ := \$18993_modulo6684349_arg\(0 to 30);
                  \$18990_modulo6684357_result\ := \$18993_modulo6684349_result\;
                  \$18989_r\ := \$18990_modulo6684357_result\;
                  \$18981_res\ := eclat_if(work.Int.lt(\$18977_binop_int6434365_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$18989_r\) & \$18989_r\);
                  \$18977_binop_int6434365_result\ := work.Int.add(\$18977_binop_int6434365_arg\(32 to 47), X"000" & X"1") & \$18981_res\ & eclat_true & 
                  work.Int.sub(\$18977_binop_int6434365_arg\(80 to 95), X"000" & X"1") & \$18977_binop_int6434365_arg\(96 to 151) & \$18977_binop_int6434365_arg\(152 to 153);
                  result4928 := \$18977_binop_int6434365_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$18993_modulo6684349_arg\ := work.Int.sub(\$18993_modulo6684349_arg\(0 to 30), \$18993_modulo6684349_arg\(31 to 61)) & \$18993_modulo6684349_arg\(31 to 61);
                  state_var5920 := \$18993_MODULO6684349\;
                end if;
              when \$18996_BINOP_INT6434366\ =>
                \$v5540\ := \$ram_lock\;
                if \$v5540\(0) = '1' then
                  state_var5920 := Q_WAIT5539;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18996_binop_int6434366_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5538;
                end if;
              when \$19002_MODULO6684356\ =>
                \$v5532\ := work.Int.lt(\$19002_modulo6684356_arg\(0 to 30), \$19002_modulo6684356_arg\(31 to 61));
                if \$v5532\(0) = '1' then
                  \$19002_modulo6684356_result\ := \$19002_modulo6684356_arg\(0 to 30);
                  \$19001_r\ := \$19002_modulo6684356_result\;
                  \$19000_res\ := eclat_if(work.Int.lt(\$18996_binop_int6434366_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19001_r\) & \$19001_r\);
                  \$18996_binop_int6434366_result\ := work.Int.add(\$18996_binop_int6434366_arg\(32 to 47), X"000" & X"1") & \$19000_res\ & eclat_true & 
                  work.Int.sub(\$18996_binop_int6434366_arg\(80 to 95), X"000" & X"1") & \$18996_binop_int6434366_arg\(96 to 151) & \$18996_binop_int6434366_arg\(152 to 153);
                  result4928 := \$18996_binop_int6434366_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19005_modulo6684349_id\ := "000001011100";
                  \$19005_modulo6684349_arg\ := work.Int.sub(\$19002_modulo6684356_arg\(0 to 30), \$19002_modulo6684356_arg\(31 to 61)) & \$19002_modulo6684356_arg\(31 to 61);
                  state_var5920 := \$19005_MODULO6684349\;
                end if;
              when \$19005_MODULO6684349\ =>
                \$v5531\ := work.Int.lt(\$19005_modulo6684349_arg\(0 to 30), \$19005_modulo6684349_arg\(31 to 61));
                if \$v5531\(0) = '1' then
                  \$19005_modulo6684349_result\ := \$19005_modulo6684349_arg\(0 to 30);
                  \$19002_modulo6684356_result\ := \$19005_modulo6684349_result\;
                  \$19001_r\ := \$19002_modulo6684356_result\;
                  \$19000_res\ := eclat_if(work.Int.lt(\$18996_binop_int6434366_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19001_r\) & \$19001_r\);
                  \$18996_binop_int6434366_result\ := work.Int.add(\$18996_binop_int6434366_arg\(32 to 47), X"000" & X"1") & \$19000_res\ & eclat_true & 
                  work.Int.sub(\$18996_binop_int6434366_arg\(80 to 95), X"000" & X"1") & \$18996_binop_int6434366_arg\(96 to 151) & \$18996_binop_int6434366_arg\(152 to 153);
                  result4928 := \$18996_binop_int6434366_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19005_modulo6684349_arg\ := work.Int.sub(\$19005_modulo6684349_arg\(0 to 30), \$19005_modulo6684349_arg\(31 to 61)) & \$19005_modulo6684349_arg\(31 to 61);
                  state_var5920 := \$19005_MODULO6684349\;
                end if;
              when \$19009_MODULO6684357\ =>
                \$v5535\ := work.Int.lt(\$19009_modulo6684357_arg\(0 to 30), \$19009_modulo6684357_arg\(31 to 61));
                if \$v5535\(0) = '1' then
                  \$19009_modulo6684357_result\ := \$19009_modulo6684357_arg\(0 to 30);
                  \$19008_r\ := \$19009_modulo6684357_result\;
                  \$19000_res\ := eclat_if(work.Int.lt(\$18996_binop_int6434366_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19008_r\) & \$19008_r\);
                  \$18996_binop_int6434366_result\ := work.Int.add(\$18996_binop_int6434366_arg\(32 to 47), X"000" & X"1") & \$19000_res\ & eclat_true & 
                  work.Int.sub(\$18996_binop_int6434366_arg\(80 to 95), X"000" & X"1") & \$18996_binop_int6434366_arg\(96 to 151) & \$18996_binop_int6434366_arg\(152 to 153);
                  result4928 := \$18996_binop_int6434366_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19012_modulo6684349_id\ := "000001011110";
                  \$19012_modulo6684349_arg\ := work.Int.sub(\$19009_modulo6684357_arg\(0 to 30), \$19009_modulo6684357_arg\(31 to 61)) & \$19009_modulo6684357_arg\(31 to 61);
                  state_var5920 := \$19012_MODULO6684349\;
                end if;
              when \$19012_MODULO6684349\ =>
                \$v5534\ := work.Int.lt(\$19012_modulo6684349_arg\(0 to 30), \$19012_modulo6684349_arg\(31 to 61));
                if \$v5534\(0) = '1' then
                  \$19012_modulo6684349_result\ := \$19012_modulo6684349_arg\(0 to 30);
                  \$19009_modulo6684357_result\ := \$19012_modulo6684349_result\;
                  \$19008_r\ := \$19009_modulo6684357_result\;
                  \$19000_res\ := eclat_if(work.Int.lt(\$18996_binop_int6434366_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19008_r\) & \$19008_r\);
                  \$18996_binop_int6434366_result\ := work.Int.add(\$18996_binop_int6434366_arg\(32 to 47), X"000" & X"1") & \$19000_res\ & eclat_true & 
                  work.Int.sub(\$18996_binop_int6434366_arg\(80 to 95), X"000" & X"1") & \$18996_binop_int6434366_arg\(96 to 151) & \$18996_binop_int6434366_arg\(152 to 153);
                  result4928 := \$18996_binop_int6434366_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19012_modulo6684349_arg\ := work.Int.sub(\$19012_modulo6684349_arg\(0 to 30), \$19012_modulo6684349_arg\(31 to 61)) & \$19012_modulo6684349_arg\(31 to 61);
                  state_var5920 := \$19012_MODULO6684349\;
                end if;
              when \$19015_BINOP_INT6434367\ =>
                \$v5550\ := \$ram_lock\;
                if \$v5550\(0) = '1' then
                  state_var5920 := Q_WAIT5549;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19015_binop_int6434367_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5548;
                end if;
              when \$19021_MODULO6684356\ =>
                \$v5542\ := work.Int.lt(\$19021_modulo6684356_arg\(0 to 30), \$19021_modulo6684356_arg\(31 to 61));
                if \$v5542\(0) = '1' then
                  \$19021_modulo6684356_result\ := \$19021_modulo6684356_arg\(0 to 30);
                  \$19020_r\ := \$19021_modulo6684356_result\;
                  \$19019_res\ := eclat_if(work.Int.lt(\$19015_binop_int6434367_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19020_r\) & \$19020_r\);
                  \$19015_binop_int6434367_result\ := work.Int.add(\$19015_binop_int6434367_arg\(32 to 47), X"000" & X"1") & \$19019_res\ & eclat_true & 
                  work.Int.sub(\$19015_binop_int6434367_arg\(80 to 95), X"000" & X"1") & \$19015_binop_int6434367_arg\(96 to 151) & \$19015_binop_int6434367_arg\(152 to 153);
                  result4928 := \$19015_binop_int6434367_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19024_modulo6684349_id\ := "000001100001";
                  \$19024_modulo6684349_arg\ := work.Int.sub(\$19021_modulo6684356_arg\(0 to 30), \$19021_modulo6684356_arg\(31 to 61)) & \$19021_modulo6684356_arg\(31 to 61);
                  state_var5920 := \$19024_MODULO6684349\;
                end if;
              when \$19024_MODULO6684349\ =>
                \$v5541\ := work.Int.lt(\$19024_modulo6684349_arg\(0 to 30), \$19024_modulo6684349_arg\(31 to 61));
                if \$v5541\(0) = '1' then
                  \$19024_modulo6684349_result\ := \$19024_modulo6684349_arg\(0 to 30);
                  \$19021_modulo6684356_result\ := \$19024_modulo6684349_result\;
                  \$19020_r\ := \$19021_modulo6684356_result\;
                  \$19019_res\ := eclat_if(work.Int.lt(\$19015_binop_int6434367_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19020_r\) & \$19020_r\);
                  \$19015_binop_int6434367_result\ := work.Int.add(\$19015_binop_int6434367_arg\(32 to 47), X"000" & X"1") & \$19019_res\ & eclat_true & 
                  work.Int.sub(\$19015_binop_int6434367_arg\(80 to 95), X"000" & X"1") & \$19015_binop_int6434367_arg\(96 to 151) & \$19015_binop_int6434367_arg\(152 to 153);
                  result4928 := \$19015_binop_int6434367_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19024_modulo6684349_arg\ := work.Int.sub(\$19024_modulo6684349_arg\(0 to 30), \$19024_modulo6684349_arg\(31 to 61)) & \$19024_modulo6684349_arg\(31 to 61);
                  state_var5920 := \$19024_MODULO6684349\;
                end if;
              when \$19028_MODULO6684357\ =>
                \$v5545\ := work.Int.lt(\$19028_modulo6684357_arg\(0 to 30), \$19028_modulo6684357_arg\(31 to 61));
                if \$v5545\(0) = '1' then
                  \$19028_modulo6684357_result\ := \$19028_modulo6684357_arg\(0 to 30);
                  \$19027_r\ := \$19028_modulo6684357_result\;
                  \$19019_res\ := eclat_if(work.Int.lt(\$19015_binop_int6434367_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19027_r\) & \$19027_r\);
                  \$19015_binop_int6434367_result\ := work.Int.add(\$19015_binop_int6434367_arg\(32 to 47), X"000" & X"1") & \$19019_res\ & eclat_true & 
                  work.Int.sub(\$19015_binop_int6434367_arg\(80 to 95), X"000" & X"1") & \$19015_binop_int6434367_arg\(96 to 151) & \$19015_binop_int6434367_arg\(152 to 153);
                  result4928 := \$19015_binop_int6434367_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19031_modulo6684349_id\ := "000001100011";
                  \$19031_modulo6684349_arg\ := work.Int.sub(\$19028_modulo6684357_arg\(0 to 30), \$19028_modulo6684357_arg\(31 to 61)) & \$19028_modulo6684357_arg\(31 to 61);
                  state_var5920 := \$19031_MODULO6684349\;
                end if;
              when \$19031_MODULO6684349\ =>
                \$v5544\ := work.Int.lt(\$19031_modulo6684349_arg\(0 to 30), \$19031_modulo6684349_arg\(31 to 61));
                if \$v5544\(0) = '1' then
                  \$19031_modulo6684349_result\ := \$19031_modulo6684349_arg\(0 to 30);
                  \$19028_modulo6684357_result\ := \$19031_modulo6684349_result\;
                  \$19027_r\ := \$19028_modulo6684357_result\;
                  \$19019_res\ := eclat_if(work.Int.lt(\$19015_binop_int6434367_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19027_r\) & \$19027_r\);
                  \$19015_binop_int6434367_result\ := work.Int.add(\$19015_binop_int6434367_arg\(32 to 47), X"000" & X"1") & \$19019_res\ & eclat_true & 
                  work.Int.sub(\$19015_binop_int6434367_arg\(80 to 95), X"000" & X"1") & \$19015_binop_int6434367_arg\(96 to 151) & \$19015_binop_int6434367_arg\(152 to 153);
                  result4928 := \$19015_binop_int6434367_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19031_modulo6684349_arg\ := work.Int.sub(\$19031_modulo6684349_arg\(0 to 30), \$19031_modulo6684349_arg\(31 to 61)) & \$19031_modulo6684349_arg\(31 to 61);
                  state_var5920 := \$19031_MODULO6684349\;
                end if;
              when \$19034_BINOP_INT6434368\ =>
                \$v5560\ := \$ram_lock\;
                if \$v5560\(0) = '1' then
                  state_var5920 := Q_WAIT5559;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19034_binop_int6434368_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5558;
                end if;
              when \$19040_MODULO6684356\ =>
                \$v5552\ := work.Int.lt(\$19040_modulo6684356_arg\(0 to 30), \$19040_modulo6684356_arg\(31 to 61));
                if \$v5552\(0) = '1' then
                  \$19040_modulo6684356_result\ := \$19040_modulo6684356_arg\(0 to 30);
                  \$19039_r\ := \$19040_modulo6684356_result\;
                  \$19038_res\ := eclat_if(work.Int.lt(\$19034_binop_int6434368_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19039_r\) & \$19039_r\);
                  \$19034_binop_int6434368_result\ := work.Int.add(\$19034_binop_int6434368_arg\(32 to 47), X"000" & X"1") & \$19038_res\ & eclat_true & 
                  work.Int.sub(\$19034_binop_int6434368_arg\(80 to 95), X"000" & X"1") & \$19034_binop_int6434368_arg\(96 to 151) & \$19034_binop_int6434368_arg\(152 to 153);
                  result4928 := \$19034_binop_int6434368_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19043_modulo6684349_id\ := "000001100110";
                  \$19043_modulo6684349_arg\ := work.Int.sub(\$19040_modulo6684356_arg\(0 to 30), \$19040_modulo6684356_arg\(31 to 61)) & \$19040_modulo6684356_arg\(31 to 61);
                  state_var5920 := \$19043_MODULO6684349\;
                end if;
              when \$19043_MODULO6684349\ =>
                \$v5551\ := work.Int.lt(\$19043_modulo6684349_arg\(0 to 30), \$19043_modulo6684349_arg\(31 to 61));
                if \$v5551\(0) = '1' then
                  \$19043_modulo6684349_result\ := \$19043_modulo6684349_arg\(0 to 30);
                  \$19040_modulo6684356_result\ := \$19043_modulo6684349_result\;
                  \$19039_r\ := \$19040_modulo6684356_result\;
                  \$19038_res\ := eclat_if(work.Int.lt(\$19034_binop_int6434368_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19039_r\) & \$19039_r\);
                  \$19034_binop_int6434368_result\ := work.Int.add(\$19034_binop_int6434368_arg\(32 to 47), X"000" & X"1") & \$19038_res\ & eclat_true & 
                  work.Int.sub(\$19034_binop_int6434368_arg\(80 to 95), X"000" & X"1") & \$19034_binop_int6434368_arg\(96 to 151) & \$19034_binop_int6434368_arg\(152 to 153);
                  result4928 := \$19034_binop_int6434368_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19043_modulo6684349_arg\ := work.Int.sub(\$19043_modulo6684349_arg\(0 to 30), \$19043_modulo6684349_arg\(31 to 61)) & \$19043_modulo6684349_arg\(31 to 61);
                  state_var5920 := \$19043_MODULO6684349\;
                end if;
              when \$19047_MODULO6684357\ =>
                \$v5555\ := work.Int.lt(\$19047_modulo6684357_arg\(0 to 30), \$19047_modulo6684357_arg\(31 to 61));
                if \$v5555\(0) = '1' then
                  \$19047_modulo6684357_result\ := \$19047_modulo6684357_arg\(0 to 30);
                  \$19046_r\ := \$19047_modulo6684357_result\;
                  \$19038_res\ := eclat_if(work.Int.lt(\$19034_binop_int6434368_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19046_r\) & \$19046_r\);
                  \$19034_binop_int6434368_result\ := work.Int.add(\$19034_binop_int6434368_arg\(32 to 47), X"000" & X"1") & \$19038_res\ & eclat_true & 
                  work.Int.sub(\$19034_binop_int6434368_arg\(80 to 95), X"000" & X"1") & \$19034_binop_int6434368_arg\(96 to 151) & \$19034_binop_int6434368_arg\(152 to 153);
                  result4928 := \$19034_binop_int6434368_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19050_modulo6684349_id\ := "000001101000";
                  \$19050_modulo6684349_arg\ := work.Int.sub(\$19047_modulo6684357_arg\(0 to 30), \$19047_modulo6684357_arg\(31 to 61)) & \$19047_modulo6684357_arg\(31 to 61);
                  state_var5920 := \$19050_MODULO6684349\;
                end if;
              when \$19050_MODULO6684349\ =>
                \$v5554\ := work.Int.lt(\$19050_modulo6684349_arg\(0 to 30), \$19050_modulo6684349_arg\(31 to 61));
                if \$v5554\(0) = '1' then
                  \$19050_modulo6684349_result\ := \$19050_modulo6684349_arg\(0 to 30);
                  \$19047_modulo6684357_result\ := \$19050_modulo6684349_result\;
                  \$19046_r\ := \$19047_modulo6684357_result\;
                  \$19038_res\ := eclat_if(work.Int.lt(\$19034_binop_int6434368_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19046_r\) & \$19046_r\);
                  \$19034_binop_int6434368_result\ := work.Int.add(\$19034_binop_int6434368_arg\(32 to 47), X"000" & X"1") & \$19038_res\ & eclat_true & 
                  work.Int.sub(\$19034_binop_int6434368_arg\(80 to 95), X"000" & X"1") & \$19034_binop_int6434368_arg\(96 to 151) & \$19034_binop_int6434368_arg\(152 to 153);
                  result4928 := \$19034_binop_int6434368_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19050_modulo6684349_arg\ := work.Int.sub(\$19050_modulo6684349_arg\(0 to 30), \$19050_modulo6684349_arg\(31 to 61)) & \$19050_modulo6684349_arg\(31 to 61);
                  state_var5920 := \$19050_MODULO6684349\;
                end if;
              when \$19053_BINOP_INT6434369\ =>
                \$v5570\ := \$ram_lock\;
                if \$v5570\(0) = '1' then
                  state_var5920 := Q_WAIT5569;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19053_binop_int6434369_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5568;
                end if;
              when \$19059_MODULO6684356\ =>
                \$v5562\ := work.Int.lt(\$19059_modulo6684356_arg\(0 to 30), \$19059_modulo6684356_arg\(31 to 61));
                if \$v5562\(0) = '1' then
                  \$19059_modulo6684356_result\ := \$19059_modulo6684356_arg\(0 to 30);
                  \$19058_r\ := \$19059_modulo6684356_result\;
                  \$19057_res\ := eclat_if(work.Int.lt(\$19053_binop_int6434369_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19058_r\) & \$19058_r\);
                  \$19053_binop_int6434369_result\ := work.Int.add(\$19053_binop_int6434369_arg\(32 to 47), X"000" & X"1") & \$19057_res\ & eclat_true & 
                  work.Int.sub(\$19053_binop_int6434369_arg\(80 to 95), X"000" & X"1") & \$19053_binop_int6434369_arg\(96 to 151) & \$19053_binop_int6434369_arg\(152 to 153);
                  result4928 := \$19053_binop_int6434369_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19062_modulo6684349_id\ := "000001101011";
                  \$19062_modulo6684349_arg\ := work.Int.sub(\$19059_modulo6684356_arg\(0 to 30), \$19059_modulo6684356_arg\(31 to 61)) & \$19059_modulo6684356_arg\(31 to 61);
                  state_var5920 := \$19062_MODULO6684349\;
                end if;
              when \$19062_MODULO6684349\ =>
                \$v5561\ := work.Int.lt(\$19062_modulo6684349_arg\(0 to 30), \$19062_modulo6684349_arg\(31 to 61));
                if \$v5561\(0) = '1' then
                  \$19062_modulo6684349_result\ := \$19062_modulo6684349_arg\(0 to 30);
                  \$19059_modulo6684356_result\ := \$19062_modulo6684349_result\;
                  \$19058_r\ := \$19059_modulo6684356_result\;
                  \$19057_res\ := eclat_if(work.Int.lt(\$19053_binop_int6434369_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19058_r\) & \$19058_r\);
                  \$19053_binop_int6434369_result\ := work.Int.add(\$19053_binop_int6434369_arg\(32 to 47), X"000" & X"1") & \$19057_res\ & eclat_true & 
                  work.Int.sub(\$19053_binop_int6434369_arg\(80 to 95), X"000" & X"1") & \$19053_binop_int6434369_arg\(96 to 151) & \$19053_binop_int6434369_arg\(152 to 153);
                  result4928 := \$19053_binop_int6434369_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19062_modulo6684349_arg\ := work.Int.sub(\$19062_modulo6684349_arg\(0 to 30), \$19062_modulo6684349_arg\(31 to 61)) & \$19062_modulo6684349_arg\(31 to 61);
                  state_var5920 := \$19062_MODULO6684349\;
                end if;
              when \$19066_MODULO6684357\ =>
                \$v5565\ := work.Int.lt(\$19066_modulo6684357_arg\(0 to 30), \$19066_modulo6684357_arg\(31 to 61));
                if \$v5565\(0) = '1' then
                  \$19066_modulo6684357_result\ := \$19066_modulo6684357_arg\(0 to 30);
                  \$19065_r\ := \$19066_modulo6684357_result\;
                  \$19057_res\ := eclat_if(work.Int.lt(\$19053_binop_int6434369_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19065_r\) & \$19065_r\);
                  \$19053_binop_int6434369_result\ := work.Int.add(\$19053_binop_int6434369_arg\(32 to 47), X"000" & X"1") & \$19057_res\ & eclat_true & 
                  work.Int.sub(\$19053_binop_int6434369_arg\(80 to 95), X"000" & X"1") & \$19053_binop_int6434369_arg\(96 to 151) & \$19053_binop_int6434369_arg\(152 to 153);
                  result4928 := \$19053_binop_int6434369_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19069_modulo6684349_id\ := "000001101101";
                  \$19069_modulo6684349_arg\ := work.Int.sub(\$19066_modulo6684357_arg\(0 to 30), \$19066_modulo6684357_arg\(31 to 61)) & \$19066_modulo6684357_arg\(31 to 61);
                  state_var5920 := \$19069_MODULO6684349\;
                end if;
              when \$19069_MODULO6684349\ =>
                \$v5564\ := work.Int.lt(\$19069_modulo6684349_arg\(0 to 30), \$19069_modulo6684349_arg\(31 to 61));
                if \$v5564\(0) = '1' then
                  \$19069_modulo6684349_result\ := \$19069_modulo6684349_arg\(0 to 30);
                  \$19066_modulo6684357_result\ := \$19069_modulo6684349_result\;
                  \$19065_r\ := \$19066_modulo6684357_result\;
                  \$19057_res\ := eclat_if(work.Int.lt(\$19053_binop_int6434369_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19065_r\) & \$19065_r\);
                  \$19053_binop_int6434369_result\ := work.Int.add(\$19053_binop_int6434369_arg\(32 to 47), X"000" & X"1") & \$19057_res\ & eclat_true & 
                  work.Int.sub(\$19053_binop_int6434369_arg\(80 to 95), X"000" & X"1") & \$19053_binop_int6434369_arg\(96 to 151) & \$19053_binop_int6434369_arg\(152 to 153);
                  result4928 := \$19053_binop_int6434369_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19069_modulo6684349_arg\ := work.Int.sub(\$19069_modulo6684349_arg\(0 to 30), \$19069_modulo6684349_arg\(31 to 61)) & \$19069_modulo6684349_arg\(31 to 61);
                  state_var5920 := \$19069_MODULO6684349\;
                end if;
              when \$19072_BINOP_INT6434370\ =>
                \$v5580\ := \$ram_lock\;
                if \$v5580\(0) = '1' then
                  state_var5920 := Q_WAIT5579;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19072_binop_int6434370_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5578;
                end if;
              when \$19078_MODULO6684356\ =>
                \$v5572\ := work.Int.lt(\$19078_modulo6684356_arg\(0 to 30), \$19078_modulo6684356_arg\(31 to 61));
                if \$v5572\(0) = '1' then
                  \$19078_modulo6684356_result\ := \$19078_modulo6684356_arg\(0 to 30);
                  \$19077_r\ := \$19078_modulo6684356_result\;
                  \$19076_res\ := eclat_if(work.Int.lt(\$19072_binop_int6434370_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19077_r\) & \$19077_r\);
                  \$19072_binop_int6434370_result\ := work.Int.add(\$19072_binop_int6434370_arg\(32 to 47), X"000" & X"1") & \$19076_res\ & eclat_true & 
                  work.Int.sub(\$19072_binop_int6434370_arg\(80 to 95), X"000" & X"1") & \$19072_binop_int6434370_arg\(96 to 151) & \$19072_binop_int6434370_arg\(152 to 153);
                  result4928 := \$19072_binop_int6434370_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19081_modulo6684349_id\ := "000001110000";
                  \$19081_modulo6684349_arg\ := work.Int.sub(\$19078_modulo6684356_arg\(0 to 30), \$19078_modulo6684356_arg\(31 to 61)) & \$19078_modulo6684356_arg\(31 to 61);
                  state_var5920 := \$19081_MODULO6684349\;
                end if;
              when \$19081_MODULO6684349\ =>
                \$v5571\ := work.Int.lt(\$19081_modulo6684349_arg\(0 to 30), \$19081_modulo6684349_arg\(31 to 61));
                if \$v5571\(0) = '1' then
                  \$19081_modulo6684349_result\ := \$19081_modulo6684349_arg\(0 to 30);
                  \$19078_modulo6684356_result\ := \$19081_modulo6684349_result\;
                  \$19077_r\ := \$19078_modulo6684356_result\;
                  \$19076_res\ := eclat_if(work.Int.lt(\$19072_binop_int6434370_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19077_r\) & \$19077_r\);
                  \$19072_binop_int6434370_result\ := work.Int.add(\$19072_binop_int6434370_arg\(32 to 47), X"000" & X"1") & \$19076_res\ & eclat_true & 
                  work.Int.sub(\$19072_binop_int6434370_arg\(80 to 95), X"000" & X"1") & \$19072_binop_int6434370_arg\(96 to 151) & \$19072_binop_int6434370_arg\(152 to 153);
                  result4928 := \$19072_binop_int6434370_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19081_modulo6684349_arg\ := work.Int.sub(\$19081_modulo6684349_arg\(0 to 30), \$19081_modulo6684349_arg\(31 to 61)) & \$19081_modulo6684349_arg\(31 to 61);
                  state_var5920 := \$19081_MODULO6684349\;
                end if;
              when \$19085_MODULO6684357\ =>
                \$v5575\ := work.Int.lt(\$19085_modulo6684357_arg\(0 to 30), \$19085_modulo6684357_arg\(31 to 61));
                if \$v5575\(0) = '1' then
                  \$19085_modulo6684357_result\ := \$19085_modulo6684357_arg\(0 to 30);
                  \$19084_r\ := \$19085_modulo6684357_result\;
                  \$19076_res\ := eclat_if(work.Int.lt(\$19072_binop_int6434370_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19084_r\) & \$19084_r\);
                  \$19072_binop_int6434370_result\ := work.Int.add(\$19072_binop_int6434370_arg\(32 to 47), X"000" & X"1") & \$19076_res\ & eclat_true & 
                  work.Int.sub(\$19072_binop_int6434370_arg\(80 to 95), X"000" & X"1") & \$19072_binop_int6434370_arg\(96 to 151) & \$19072_binop_int6434370_arg\(152 to 153);
                  result4928 := \$19072_binop_int6434370_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19088_modulo6684349_id\ := "000001110010";
                  \$19088_modulo6684349_arg\ := work.Int.sub(\$19085_modulo6684357_arg\(0 to 30), \$19085_modulo6684357_arg\(31 to 61)) & \$19085_modulo6684357_arg\(31 to 61);
                  state_var5920 := \$19088_MODULO6684349\;
                end if;
              when \$19088_MODULO6684349\ =>
                \$v5574\ := work.Int.lt(\$19088_modulo6684349_arg\(0 to 30), \$19088_modulo6684349_arg\(31 to 61));
                if \$v5574\(0) = '1' then
                  \$19088_modulo6684349_result\ := \$19088_modulo6684349_arg\(0 to 30);
                  \$19085_modulo6684357_result\ := \$19088_modulo6684349_result\;
                  \$19084_r\ := \$19085_modulo6684357_result\;
                  \$19076_res\ := eclat_if(work.Int.lt(\$19072_binop_int6434370_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19084_r\) & \$19084_r\);
                  \$19072_binop_int6434370_result\ := work.Int.add(\$19072_binop_int6434370_arg\(32 to 47), X"000" & X"1") & \$19076_res\ & eclat_true & 
                  work.Int.sub(\$19072_binop_int6434370_arg\(80 to 95), X"000" & X"1") & \$19072_binop_int6434370_arg\(96 to 151) & \$19072_binop_int6434370_arg\(152 to 153);
                  result4928 := \$19072_binop_int6434370_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19088_modulo6684349_arg\ := work.Int.sub(\$19088_modulo6684349_arg\(0 to 30), \$19088_modulo6684349_arg\(31 to 61)) & \$19088_modulo6684349_arg\(31 to 61);
                  state_var5920 := \$19088_MODULO6684349\;
                end if;
              when \$19091_BINOP_INT6434371\ =>
                \$v5590\ := \$ram_lock\;
                if \$v5590\(0) = '1' then
                  state_var5920 := Q_WAIT5589;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19091_binop_int6434371_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5588;
                end if;
              when \$19097_MODULO6684356\ =>
                \$v5582\ := work.Int.lt(\$19097_modulo6684356_arg\(0 to 30), \$19097_modulo6684356_arg\(31 to 61));
                if \$v5582\(0) = '1' then
                  \$19097_modulo6684356_result\ := \$19097_modulo6684356_arg\(0 to 30);
                  \$19096_r\ := \$19097_modulo6684356_result\;
                  \$19095_res\ := eclat_if(work.Int.lt(\$19091_binop_int6434371_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19096_r\) & \$19096_r\);
                  \$19091_binop_int6434371_result\ := work.Int.add(\$19091_binop_int6434371_arg\(32 to 47), X"000" & X"1") & \$19095_res\ & eclat_true & 
                  work.Int.sub(\$19091_binop_int6434371_arg\(80 to 95), X"000" & X"1") & \$19091_binop_int6434371_arg\(96 to 151) & \$19091_binop_int6434371_arg\(152 to 153);
                  result4928 := \$19091_binop_int6434371_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19100_modulo6684349_id\ := "000001110101";
                  \$19100_modulo6684349_arg\ := work.Int.sub(\$19097_modulo6684356_arg\(0 to 30), \$19097_modulo6684356_arg\(31 to 61)) & \$19097_modulo6684356_arg\(31 to 61);
                  state_var5920 := \$19100_MODULO6684349\;
                end if;
              when \$19100_MODULO6684349\ =>
                \$v5581\ := work.Int.lt(\$19100_modulo6684349_arg\(0 to 30), \$19100_modulo6684349_arg\(31 to 61));
                if \$v5581\(0) = '1' then
                  \$19100_modulo6684349_result\ := \$19100_modulo6684349_arg\(0 to 30);
                  \$19097_modulo6684356_result\ := \$19100_modulo6684349_result\;
                  \$19096_r\ := \$19097_modulo6684356_result\;
                  \$19095_res\ := eclat_if(work.Int.lt(\$19091_binop_int6434371_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19096_r\) & \$19096_r\);
                  \$19091_binop_int6434371_result\ := work.Int.add(\$19091_binop_int6434371_arg\(32 to 47), X"000" & X"1") & \$19095_res\ & eclat_true & 
                  work.Int.sub(\$19091_binop_int6434371_arg\(80 to 95), X"000" & X"1") & \$19091_binop_int6434371_arg\(96 to 151) & \$19091_binop_int6434371_arg\(152 to 153);
                  result4928 := \$19091_binop_int6434371_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19100_modulo6684349_arg\ := work.Int.sub(\$19100_modulo6684349_arg\(0 to 30), \$19100_modulo6684349_arg\(31 to 61)) & \$19100_modulo6684349_arg\(31 to 61);
                  state_var5920 := \$19100_MODULO6684349\;
                end if;
              when \$19104_MODULO6684357\ =>
                \$v5585\ := work.Int.lt(\$19104_modulo6684357_arg\(0 to 30), \$19104_modulo6684357_arg\(31 to 61));
                if \$v5585\(0) = '1' then
                  \$19104_modulo6684357_result\ := \$19104_modulo6684357_arg\(0 to 30);
                  \$19103_r\ := \$19104_modulo6684357_result\;
                  \$19095_res\ := eclat_if(work.Int.lt(\$19091_binop_int6434371_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19103_r\) & \$19103_r\);
                  \$19091_binop_int6434371_result\ := work.Int.add(\$19091_binop_int6434371_arg\(32 to 47), X"000" & X"1") & \$19095_res\ & eclat_true & 
                  work.Int.sub(\$19091_binop_int6434371_arg\(80 to 95), X"000" & X"1") & \$19091_binop_int6434371_arg\(96 to 151) & \$19091_binop_int6434371_arg\(152 to 153);
                  result4928 := \$19091_binop_int6434371_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19107_modulo6684349_id\ := "000001110111";
                  \$19107_modulo6684349_arg\ := work.Int.sub(\$19104_modulo6684357_arg\(0 to 30), \$19104_modulo6684357_arg\(31 to 61)) & \$19104_modulo6684357_arg\(31 to 61);
                  state_var5920 := \$19107_MODULO6684349\;
                end if;
              when \$19107_MODULO6684349\ =>
                \$v5584\ := work.Int.lt(\$19107_modulo6684349_arg\(0 to 30), \$19107_modulo6684349_arg\(31 to 61));
                if \$v5584\(0) = '1' then
                  \$19107_modulo6684349_result\ := \$19107_modulo6684349_arg\(0 to 30);
                  \$19104_modulo6684357_result\ := \$19107_modulo6684349_result\;
                  \$19103_r\ := \$19104_modulo6684357_result\;
                  \$19095_res\ := eclat_if(work.Int.lt(\$19091_binop_int6434371_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19103_r\) & \$19103_r\);
                  \$19091_binop_int6434371_result\ := work.Int.add(\$19091_binop_int6434371_arg\(32 to 47), X"000" & X"1") & \$19095_res\ & eclat_true & 
                  work.Int.sub(\$19091_binop_int6434371_arg\(80 to 95), X"000" & X"1") & \$19091_binop_int6434371_arg\(96 to 151) & \$19091_binop_int6434371_arg\(152 to 153);
                  result4928 := \$19091_binop_int6434371_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19107_modulo6684349_arg\ := work.Int.sub(\$19107_modulo6684349_arg\(0 to 30), \$19107_modulo6684349_arg\(31 to 61)) & \$19107_modulo6684349_arg\(31 to 61);
                  state_var5920 := \$19107_MODULO6684349\;
                end if;
              when \$19113_FOREVER6704372\ =>
                \$19113_forever6704372_arg\ := eclat_unit;
                state_var5920 := \$19113_FOREVER6704372\;
              when \$19116_BINOP_INT6434373\ =>
                \$v5600\ := \$ram_lock\;
                if \$v5600\(0) = '1' then
                  state_var5920 := Q_WAIT5599;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19116_binop_int6434373_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5598;
                end if;
              when \$19122_MODULO6684356\ =>
                \$v5592\ := work.Int.lt(\$19122_modulo6684356_arg\(0 to 30), \$19122_modulo6684356_arg\(31 to 61));
                if \$v5592\(0) = '1' then
                  \$19122_modulo6684356_result\ := \$19122_modulo6684356_arg\(0 to 30);
                  \$19121_r\ := \$19122_modulo6684356_result\;
                  \$19120_res\ := eclat_if(work.Int.lt(\$19116_binop_int6434373_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19121_r\) & \$19121_r\);
                  \$19116_binop_int6434373_result\ := work.Int.add(\$19116_binop_int6434373_arg\(32 to 47), X"000" & X"1") & \$19120_res\ & eclat_true & 
                  work.Int.sub(\$19116_binop_int6434373_arg\(80 to 95), X"000" & X"1") & \$19116_binop_int6434373_arg\(96 to 151) & \$19116_binop_int6434373_arg\(152 to 153);
                  result4928 := \$19116_binop_int6434373_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19125_modulo6684349_id\ := "000001111011";
                  \$19125_modulo6684349_arg\ := work.Int.sub(\$19122_modulo6684356_arg\(0 to 30), \$19122_modulo6684356_arg\(31 to 61)) & \$19122_modulo6684356_arg\(31 to 61);
                  state_var5920 := \$19125_MODULO6684349\;
                end if;
              when \$19125_MODULO6684349\ =>
                \$v5591\ := work.Int.lt(\$19125_modulo6684349_arg\(0 to 30), \$19125_modulo6684349_arg\(31 to 61));
                if \$v5591\(0) = '1' then
                  \$19125_modulo6684349_result\ := \$19125_modulo6684349_arg\(0 to 30);
                  \$19122_modulo6684356_result\ := \$19125_modulo6684349_result\;
                  \$19121_r\ := \$19122_modulo6684356_result\;
                  \$19120_res\ := eclat_if(work.Int.lt(\$19116_binop_int6434373_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19121_r\) & \$19121_r\);
                  \$19116_binop_int6434373_result\ := work.Int.add(\$19116_binop_int6434373_arg\(32 to 47), X"000" & X"1") & \$19120_res\ & eclat_true & 
                  work.Int.sub(\$19116_binop_int6434373_arg\(80 to 95), X"000" & X"1") & \$19116_binop_int6434373_arg\(96 to 151) & \$19116_binop_int6434373_arg\(152 to 153);
                  result4928 := \$19116_binop_int6434373_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19125_modulo6684349_arg\ := work.Int.sub(\$19125_modulo6684349_arg\(0 to 30), \$19125_modulo6684349_arg\(31 to 61)) & \$19125_modulo6684349_arg\(31 to 61);
                  state_var5920 := \$19125_MODULO6684349\;
                end if;
              when \$19129_MODULO6684357\ =>
                \$v5595\ := work.Int.lt(\$19129_modulo6684357_arg\(0 to 30), \$19129_modulo6684357_arg\(31 to 61));
                if \$v5595\(0) = '1' then
                  \$19129_modulo6684357_result\ := \$19129_modulo6684357_arg\(0 to 30);
                  \$19128_r\ := \$19129_modulo6684357_result\;
                  \$19120_res\ := eclat_if(work.Int.lt(\$19116_binop_int6434373_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19128_r\) & \$19128_r\);
                  \$19116_binop_int6434373_result\ := work.Int.add(\$19116_binop_int6434373_arg\(32 to 47), X"000" & X"1") & \$19120_res\ & eclat_true & 
                  work.Int.sub(\$19116_binop_int6434373_arg\(80 to 95), X"000" & X"1") & \$19116_binop_int6434373_arg\(96 to 151) & \$19116_binop_int6434373_arg\(152 to 153);
                  result4928 := \$19116_binop_int6434373_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19132_modulo6684349_id\ := "000001111101";
                  \$19132_modulo6684349_arg\ := work.Int.sub(\$19129_modulo6684357_arg\(0 to 30), \$19129_modulo6684357_arg\(31 to 61)) & \$19129_modulo6684357_arg\(31 to 61);
                  state_var5920 := \$19132_MODULO6684349\;
                end if;
              when \$19132_MODULO6684349\ =>
                \$v5594\ := work.Int.lt(\$19132_modulo6684349_arg\(0 to 30), \$19132_modulo6684349_arg\(31 to 61));
                if \$v5594\(0) = '1' then
                  \$19132_modulo6684349_result\ := \$19132_modulo6684349_arg\(0 to 30);
                  \$19129_modulo6684357_result\ := \$19132_modulo6684349_result\;
                  \$19128_r\ := \$19129_modulo6684357_result\;
                  \$19120_res\ := eclat_if(work.Int.lt(\$19116_binop_int6434373_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19128_r\) & \$19128_r\);
                  \$19116_binop_int6434373_result\ := work.Int.add(\$19116_binop_int6434373_arg\(32 to 47), X"000" & X"1") & \$19120_res\ & eclat_true & 
                  work.Int.sub(\$19116_binop_int6434373_arg\(80 to 95), X"000" & X"1") & \$19116_binop_int6434373_arg\(96 to 151) & \$19116_binop_int6434373_arg\(152 to 153);
                  result4928 := \$19116_binop_int6434373_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19132_modulo6684349_arg\ := work.Int.sub(\$19132_modulo6684349_arg\(0 to 30), \$19132_modulo6684349_arg\(31 to 61)) & \$19132_modulo6684349_arg\(31 to 61);
                  state_var5920 := \$19132_MODULO6684349\;
                end if;
              when \$19135_BINOP_INT6434374\ =>
                \$v5610\ := \$ram_lock\;
                if \$v5610\(0) = '1' then
                  state_var5920 := Q_WAIT5609;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19135_binop_int6434374_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5608;
                end if;
              when \$19141_MODULO6684356\ =>
                \$v5602\ := work.Int.lt(\$19141_modulo6684356_arg\(0 to 30), \$19141_modulo6684356_arg\(31 to 61));
                if \$v5602\(0) = '1' then
                  \$19141_modulo6684356_result\ := \$19141_modulo6684356_arg\(0 to 30);
                  \$19140_r\ := \$19141_modulo6684356_result\;
                  \$19139_res\ := eclat_if(work.Int.lt(\$19135_binop_int6434374_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19140_r\) & \$19140_r\);
                  \$19135_binop_int6434374_result\ := work.Int.add(\$19135_binop_int6434374_arg\(32 to 47), X"000" & X"1") & \$19139_res\ & eclat_true & 
                  work.Int.sub(\$19135_binop_int6434374_arg\(80 to 95), X"000" & X"1") & \$19135_binop_int6434374_arg\(96 to 151) & \$19135_binop_int6434374_arg\(152 to 153);
                  result4928 := \$19135_binop_int6434374_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19144_modulo6684349_id\ := "000010000000";
                  \$19144_modulo6684349_arg\ := work.Int.sub(\$19141_modulo6684356_arg\(0 to 30), \$19141_modulo6684356_arg\(31 to 61)) & \$19141_modulo6684356_arg\(31 to 61);
                  state_var5920 := \$19144_MODULO6684349\;
                end if;
              when \$19144_MODULO6684349\ =>
                \$v5601\ := work.Int.lt(\$19144_modulo6684349_arg\(0 to 30), \$19144_modulo6684349_arg\(31 to 61));
                if \$v5601\(0) = '1' then
                  \$19144_modulo6684349_result\ := \$19144_modulo6684349_arg\(0 to 30);
                  \$19141_modulo6684356_result\ := \$19144_modulo6684349_result\;
                  \$19140_r\ := \$19141_modulo6684356_result\;
                  \$19139_res\ := eclat_if(work.Int.lt(\$19135_binop_int6434374_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19140_r\) & \$19140_r\);
                  \$19135_binop_int6434374_result\ := work.Int.add(\$19135_binop_int6434374_arg\(32 to 47), X"000" & X"1") & \$19139_res\ & eclat_true & 
                  work.Int.sub(\$19135_binop_int6434374_arg\(80 to 95), X"000" & X"1") & \$19135_binop_int6434374_arg\(96 to 151) & \$19135_binop_int6434374_arg\(152 to 153);
                  result4928 := \$19135_binop_int6434374_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19144_modulo6684349_arg\ := work.Int.sub(\$19144_modulo6684349_arg\(0 to 30), \$19144_modulo6684349_arg\(31 to 61)) & \$19144_modulo6684349_arg\(31 to 61);
                  state_var5920 := \$19144_MODULO6684349\;
                end if;
              when \$19148_MODULO6684357\ =>
                \$v5605\ := work.Int.lt(\$19148_modulo6684357_arg\(0 to 30), \$19148_modulo6684357_arg\(31 to 61));
                if \$v5605\(0) = '1' then
                  \$19148_modulo6684357_result\ := \$19148_modulo6684357_arg\(0 to 30);
                  \$19147_r\ := \$19148_modulo6684357_result\;
                  \$19139_res\ := eclat_if(work.Int.lt(\$19135_binop_int6434374_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19147_r\) & \$19147_r\);
                  \$19135_binop_int6434374_result\ := work.Int.add(\$19135_binop_int6434374_arg\(32 to 47), X"000" & X"1") & \$19139_res\ & eclat_true & 
                  work.Int.sub(\$19135_binop_int6434374_arg\(80 to 95), X"000" & X"1") & \$19135_binop_int6434374_arg\(96 to 151) & \$19135_binop_int6434374_arg\(152 to 153);
                  result4928 := \$19135_binop_int6434374_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19151_modulo6684349_id\ := "000010000010";
                  \$19151_modulo6684349_arg\ := work.Int.sub(\$19148_modulo6684357_arg\(0 to 30), \$19148_modulo6684357_arg\(31 to 61)) & \$19148_modulo6684357_arg\(31 to 61);
                  state_var5920 := \$19151_MODULO6684349\;
                end if;
              when \$19151_MODULO6684349\ =>
                \$v5604\ := work.Int.lt(\$19151_modulo6684349_arg\(0 to 30), \$19151_modulo6684349_arg\(31 to 61));
                if \$v5604\(0) = '1' then
                  \$19151_modulo6684349_result\ := \$19151_modulo6684349_arg\(0 to 30);
                  \$19148_modulo6684357_result\ := \$19151_modulo6684349_result\;
                  \$19147_r\ := \$19148_modulo6684357_result\;
                  \$19139_res\ := eclat_if(work.Int.lt(\$19135_binop_int6434374_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$19147_r\) & \$19147_r\);
                  \$19135_binop_int6434374_result\ := work.Int.add(\$19135_binop_int6434374_arg\(32 to 47), X"000" & X"1") & \$19139_res\ & eclat_true & 
                  work.Int.sub(\$19135_binop_int6434374_arg\(80 to 95), X"000" & X"1") & \$19135_binop_int6434374_arg\(96 to 151) & \$19135_binop_int6434374_arg\(152 to 153);
                  result4928 := \$19135_binop_int6434374_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$19151_modulo6684349_arg\ := work.Int.sub(\$19151_modulo6684349_arg\(0 to 30), \$19151_modulo6684349_arg\(31 to 61)) & \$19151_modulo6684349_arg\(31 to 61);
                  state_var5920 := \$19151_MODULO6684349\;
                end if;
              when \$19157_FOREVER6704375\ =>
                \$19157_forever6704375_arg\ := eclat_unit;
                state_var5920 := \$19157_FOREVER6704375\;
              when \$19163_FOREVER6704376\ =>
                \$19163_forever6704376_arg\ := eclat_unit;
                state_var5920 := \$19163_FOREVER6704376\;
              when \$19166_BINOP_COMPARE6454377\ =>
                \$v5614\ := \$ram_lock\;
                if \$v5614\(0) = '1' then
                  state_var5920 := Q_WAIT5613;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19166_binop_compare6454377_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5612;
                end if;
              when \$19171_COMPARE6444358\ =>
                \$v5611\ := \$19171_compare6444358_arg\(0 to 31);
                case \$v5611\ is
                when X"0000000" & X"0" =>
                  \$19171_compare6444358_result\ := work.Int.eq(\$19171_compare6444358_arg\(32 to 62), \$19171_compare6444358_arg\(63 to 93));
                when X"0000000" & X"1" =>
                  \$19171_compare6444358_result\ := work.Bool.lnot(work.Int.eq(
                                                                   \$19171_compare6444358_arg\(32 to 62), \$19171_compare6444358_arg\(63 to 93)));
                when X"0000000" & X"2" =>
                  \$19171_compare6444358_result\ := work.Int.lt(\$19171_compare6444358_arg\(32 to 62), \$19171_compare6444358_arg\(63 to 93));
                when X"0000000" & X"3" =>
                  \$19171_compare6444358_result\ := eclat_if(work.Int.lt(
                                                             \$19171_compare6444358_arg\(32 to 62), \$19171_compare6444358_arg\(63 to 93)) & eclat_true & 
                                                    work.Int.eq(\$19171_compare6444358_arg\(32 to 62), \$19171_compare6444358_arg\(63 to 93)));
                when X"0000000" & X"4" =>
                  \$19171_compare6444358_result\ := work.Bool.lnot(eclat_if(
                                                                   work.Int.lt(
                                                                   \$19171_compare6444358_arg\(32 to 62), \$19171_compare6444358_arg\(63 to 93)) & eclat_true & 
                                                                   work.Int.eq(
                                                                   \$19171_compare6444358_arg\(32 to 62), \$19171_compare6444358_arg\(63 to 93))));
                when X"0000000" & X"5" =>
                  \$19171_compare6444358_result\ := work.Bool.lnot(work.Int.lt(
                                                                   \$19171_compare6444358_arg\(32 to 62), \$19171_compare6444358_arg\(63 to 93)));
                when others =>
                  \$19171_compare6444358_result\ := eclat_false;
                end case;
                \$19170_res\ := \$19171_compare6444358_result\;
                \$19166_binop_compare6454377_result\ := work.Int.add(
                                                        \$19166_binop_compare6454377_arg\(32 to 47), X"000" & X"1") & 
                eclat_if(\$19170_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & 
                work.Int.sub(\$19166_binop_compare6454377_arg\(80 to 95), X"000" & X"1") & \$19166_binop_compare6454377_arg\(96 to 151) & \$19166_binop_compare6454377_arg\(152 to 153);
                result4928 := \$19166_binop_compare6454377_result\;
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when \$19174_BINOP_COMPARE6454378\ =>
                \$v5618\ := \$ram_lock\;
                if \$v5618\(0) = '1' then
                  state_var5920 := Q_WAIT5617;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19174_binop_compare6454378_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5616;
                end if;
              when \$19179_COMPARE6444358\ =>
                \$v5615\ := \$19179_compare6444358_arg\(0 to 31);
                case \$v5615\ is
                when X"0000000" & X"0" =>
                  \$19179_compare6444358_result\ := work.Int.eq(\$19179_compare6444358_arg\(32 to 62), \$19179_compare6444358_arg\(63 to 93));
                when X"0000000" & X"1" =>
                  \$19179_compare6444358_result\ := work.Bool.lnot(work.Int.eq(
                                                                   \$19179_compare6444358_arg\(32 to 62), \$19179_compare6444358_arg\(63 to 93)));
                when X"0000000" & X"2" =>
                  \$19179_compare6444358_result\ := work.Int.lt(\$19179_compare6444358_arg\(32 to 62), \$19179_compare6444358_arg\(63 to 93));
                when X"0000000" & X"3" =>
                  \$19179_compare6444358_result\ := eclat_if(work.Int.lt(
                                                             \$19179_compare6444358_arg\(32 to 62), \$19179_compare6444358_arg\(63 to 93)) & eclat_true & 
                                                    work.Int.eq(\$19179_compare6444358_arg\(32 to 62), \$19179_compare6444358_arg\(63 to 93)));
                when X"0000000" & X"4" =>
                  \$19179_compare6444358_result\ := work.Bool.lnot(eclat_if(
                                                                   work.Int.lt(
                                                                   \$19179_compare6444358_arg\(32 to 62), \$19179_compare6444358_arg\(63 to 93)) & eclat_true & 
                                                                   work.Int.eq(
                                                                   \$19179_compare6444358_arg\(32 to 62), \$19179_compare6444358_arg\(63 to 93))));
                when X"0000000" & X"5" =>
                  \$19179_compare6444358_result\ := work.Bool.lnot(work.Int.lt(
                                                                   \$19179_compare6444358_arg\(32 to 62), \$19179_compare6444358_arg\(63 to 93)));
                when others =>
                  \$19179_compare6444358_result\ := eclat_false;
                end case;
                \$19178_res\ := \$19179_compare6444358_result\;
                \$19174_binop_compare6454378_result\ := work.Int.add(
                                                        \$19174_binop_compare6454378_arg\(32 to 47), X"000" & X"1") & 
                eclat_if(\$19178_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & 
                work.Int.sub(\$19174_binop_compare6454378_arg\(80 to 95), X"000" & X"1") & \$19174_binop_compare6454378_arg\(96 to 151) & \$19174_binop_compare6454378_arg\(152 to 153);
                result4928 := \$19174_binop_compare6454378_result\;
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when \$19182_BINOP_COMPARE6454379\ =>
                \$v5622\ := \$ram_lock\;
                if \$v5622\(0) = '1' then
                  state_var5920 := Q_WAIT5621;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19182_binop_compare6454379_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5620;
                end if;
              when \$19187_COMPARE6444358\ =>
                \$v5619\ := \$19187_compare6444358_arg\(0 to 31);
                case \$v5619\ is
                when X"0000000" & X"0" =>
                  \$19187_compare6444358_result\ := work.Int.eq(\$19187_compare6444358_arg\(32 to 62), \$19187_compare6444358_arg\(63 to 93));
                when X"0000000" & X"1" =>
                  \$19187_compare6444358_result\ := work.Bool.lnot(work.Int.eq(
                                                                   \$19187_compare6444358_arg\(32 to 62), \$19187_compare6444358_arg\(63 to 93)));
                when X"0000000" & X"2" =>
                  \$19187_compare6444358_result\ := work.Int.lt(\$19187_compare6444358_arg\(32 to 62), \$19187_compare6444358_arg\(63 to 93));
                when X"0000000" & X"3" =>
                  \$19187_compare6444358_result\ := eclat_if(work.Int.lt(
                                                             \$19187_compare6444358_arg\(32 to 62), \$19187_compare6444358_arg\(63 to 93)) & eclat_true & 
                                                    work.Int.eq(\$19187_compare6444358_arg\(32 to 62), \$19187_compare6444358_arg\(63 to 93)));
                when X"0000000" & X"4" =>
                  \$19187_compare6444358_result\ := work.Bool.lnot(eclat_if(
                                                                   work.Int.lt(
                                                                   \$19187_compare6444358_arg\(32 to 62), \$19187_compare6444358_arg\(63 to 93)) & eclat_true & 
                                                                   work.Int.eq(
                                                                   \$19187_compare6444358_arg\(32 to 62), \$19187_compare6444358_arg\(63 to 93))));
                when X"0000000" & X"5" =>
                  \$19187_compare6444358_result\ := work.Bool.lnot(work.Int.lt(
                                                                   \$19187_compare6444358_arg\(32 to 62), \$19187_compare6444358_arg\(63 to 93)));
                when others =>
                  \$19187_compare6444358_result\ := eclat_false;
                end case;
                \$19186_res\ := \$19187_compare6444358_result\;
                \$19182_binop_compare6454379_result\ := work.Int.add(
                                                        \$19182_binop_compare6454379_arg\(32 to 47), X"000" & X"1") & 
                eclat_if(\$19186_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & 
                work.Int.sub(\$19182_binop_compare6454379_arg\(80 to 95), X"000" & X"1") & \$19182_binop_compare6454379_arg\(96 to 151) & \$19182_binop_compare6454379_arg\(152 to 153);
                result4928 := \$19182_binop_compare6454379_result\;
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when \$19190_BINOP_COMPARE6454380\ =>
                \$v5626\ := \$ram_lock\;
                if \$v5626\(0) = '1' then
                  state_var5920 := Q_WAIT5625;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19190_binop_compare6454380_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5624;
                end if;
              when \$19195_COMPARE6444358\ =>
                \$v5623\ := \$19195_compare6444358_arg\(0 to 31);
                case \$v5623\ is
                when X"0000000" & X"0" =>
                  \$19195_compare6444358_result\ := work.Int.eq(\$19195_compare6444358_arg\(32 to 62), \$19195_compare6444358_arg\(63 to 93));
                when X"0000000" & X"1" =>
                  \$19195_compare6444358_result\ := work.Bool.lnot(work.Int.eq(
                                                                   \$19195_compare6444358_arg\(32 to 62), \$19195_compare6444358_arg\(63 to 93)));
                when X"0000000" & X"2" =>
                  \$19195_compare6444358_result\ := work.Int.lt(\$19195_compare6444358_arg\(32 to 62), \$19195_compare6444358_arg\(63 to 93));
                when X"0000000" & X"3" =>
                  \$19195_compare6444358_result\ := eclat_if(work.Int.lt(
                                                             \$19195_compare6444358_arg\(32 to 62), \$19195_compare6444358_arg\(63 to 93)) & eclat_true & 
                                                    work.Int.eq(\$19195_compare6444358_arg\(32 to 62), \$19195_compare6444358_arg\(63 to 93)));
                when X"0000000" & X"4" =>
                  \$19195_compare6444358_result\ := work.Bool.lnot(eclat_if(
                                                                   work.Int.lt(
                                                                   \$19195_compare6444358_arg\(32 to 62), \$19195_compare6444358_arg\(63 to 93)) & eclat_true & 
                                                                   work.Int.eq(
                                                                   \$19195_compare6444358_arg\(32 to 62), \$19195_compare6444358_arg\(63 to 93))));
                when X"0000000" & X"5" =>
                  \$19195_compare6444358_result\ := work.Bool.lnot(work.Int.lt(
                                                                   \$19195_compare6444358_arg\(32 to 62), \$19195_compare6444358_arg\(63 to 93)));
                when others =>
                  \$19195_compare6444358_result\ := eclat_false;
                end case;
                \$19194_res\ := \$19195_compare6444358_result\;
                \$19190_binop_compare6454380_result\ := work.Int.add(
                                                        \$19190_binop_compare6454380_arg\(32 to 47), X"000" & X"1") & 
                eclat_if(\$19194_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & 
                work.Int.sub(\$19190_binop_compare6454380_arg\(80 to 95), X"000" & X"1") & \$19190_binop_compare6454380_arg\(96 to 151) & \$19190_binop_compare6454380_arg\(152 to 153);
                result4928 := \$19190_binop_compare6454380_result\;
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when \$19198_BINOP_COMPARE6454381\ =>
                \$v5630\ := \$ram_lock\;
                if \$v5630\(0) = '1' then
                  state_var5920 := Q_WAIT5629;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19198_binop_compare6454381_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5628;
                end if;
              when \$19203_COMPARE6444358\ =>
                \$v5627\ := \$19203_compare6444358_arg\(0 to 31);
                case \$v5627\ is
                when X"0000000" & X"0" =>
                  \$19203_compare6444358_result\ := work.Int.eq(\$19203_compare6444358_arg\(32 to 62), \$19203_compare6444358_arg\(63 to 93));
                when X"0000000" & X"1" =>
                  \$19203_compare6444358_result\ := work.Bool.lnot(work.Int.eq(
                                                                   \$19203_compare6444358_arg\(32 to 62), \$19203_compare6444358_arg\(63 to 93)));
                when X"0000000" & X"2" =>
                  \$19203_compare6444358_result\ := work.Int.lt(\$19203_compare6444358_arg\(32 to 62), \$19203_compare6444358_arg\(63 to 93));
                when X"0000000" & X"3" =>
                  \$19203_compare6444358_result\ := eclat_if(work.Int.lt(
                                                             \$19203_compare6444358_arg\(32 to 62), \$19203_compare6444358_arg\(63 to 93)) & eclat_true & 
                                                    work.Int.eq(\$19203_compare6444358_arg\(32 to 62), \$19203_compare6444358_arg\(63 to 93)));
                when X"0000000" & X"4" =>
                  \$19203_compare6444358_result\ := work.Bool.lnot(eclat_if(
                                                                   work.Int.lt(
                                                                   \$19203_compare6444358_arg\(32 to 62), \$19203_compare6444358_arg\(63 to 93)) & eclat_true & 
                                                                   work.Int.eq(
                                                                   \$19203_compare6444358_arg\(32 to 62), \$19203_compare6444358_arg\(63 to 93))));
                when X"0000000" & X"5" =>
                  \$19203_compare6444358_result\ := work.Bool.lnot(work.Int.lt(
                                                                   \$19203_compare6444358_arg\(32 to 62), \$19203_compare6444358_arg\(63 to 93)));
                when others =>
                  \$19203_compare6444358_result\ := eclat_false;
                end case;
                \$19202_res\ := \$19203_compare6444358_result\;
                \$19198_binop_compare6454381_result\ := work.Int.add(
                                                        \$19198_binop_compare6454381_arg\(32 to 47), X"000" & X"1") & 
                eclat_if(\$19202_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & 
                work.Int.sub(\$19198_binop_compare6454381_arg\(80 to 95), X"000" & X"1") & \$19198_binop_compare6454381_arg\(96 to 151) & \$19198_binop_compare6454381_arg\(152 to 153);
                result4928 := \$19198_binop_compare6454381_result\;
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when \$19206_BINOP_COMPARE6454382\ =>
                \$v5634\ := \$ram_lock\;
                if \$v5634\(0) = '1' then
                  state_var5920 := Q_WAIT5633;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19206_binop_compare6454382_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5632;
                end if;
              when \$19211_COMPARE6444358\ =>
                \$v5631\ := \$19211_compare6444358_arg\(0 to 31);
                case \$v5631\ is
                when X"0000000" & X"0" =>
                  \$19211_compare6444358_result\ := work.Int.eq(\$19211_compare6444358_arg\(32 to 62), \$19211_compare6444358_arg\(63 to 93));
                when X"0000000" & X"1" =>
                  \$19211_compare6444358_result\ := work.Bool.lnot(work.Int.eq(
                                                                   \$19211_compare6444358_arg\(32 to 62), \$19211_compare6444358_arg\(63 to 93)));
                when X"0000000" & X"2" =>
                  \$19211_compare6444358_result\ := work.Int.lt(\$19211_compare6444358_arg\(32 to 62), \$19211_compare6444358_arg\(63 to 93));
                when X"0000000" & X"3" =>
                  \$19211_compare6444358_result\ := eclat_if(work.Int.lt(
                                                             \$19211_compare6444358_arg\(32 to 62), \$19211_compare6444358_arg\(63 to 93)) & eclat_true & 
                                                    work.Int.eq(\$19211_compare6444358_arg\(32 to 62), \$19211_compare6444358_arg\(63 to 93)));
                when X"0000000" & X"4" =>
                  \$19211_compare6444358_result\ := work.Bool.lnot(eclat_if(
                                                                   work.Int.lt(
                                                                   \$19211_compare6444358_arg\(32 to 62), \$19211_compare6444358_arg\(63 to 93)) & eclat_true & 
                                                                   work.Int.eq(
                                                                   \$19211_compare6444358_arg\(32 to 62), \$19211_compare6444358_arg\(63 to 93))));
                when X"0000000" & X"5" =>
                  \$19211_compare6444358_result\ := work.Bool.lnot(work.Int.lt(
                                                                   \$19211_compare6444358_arg\(32 to 62), \$19211_compare6444358_arg\(63 to 93)));
                when others =>
                  \$19211_compare6444358_result\ := eclat_false;
                end case;
                \$19210_res\ := \$19211_compare6444358_result\;
                \$19206_binop_compare6454382_result\ := work.Int.add(
                                                        \$19206_binop_compare6454382_arg\(32 to 47), X"000" & X"1") & 
                eclat_if(\$19210_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & 
                work.Int.sub(\$19206_binop_compare6454382_arg\(80 to 95), X"000" & X"1") & \$19206_binop_compare6454382_arg\(96 to 151) & \$19206_binop_compare6454382_arg\(152 to 153);
                result4928 := \$19206_binop_compare6454382_result\;
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when \$19238_W6514383\ =>
                \$v5696\ := work.Int.gt(\$19238_w6514383_arg\(0 to 7), \$19238_w6514383_arg\(24 to 31));
                if \$v5696\(0) = '1' then
                  \$19238_w6514383_result\ := \$19238_w6514383_arg\(8 to 23);
                  \$19234_sp\ := \$19238_w6514383_result\;
                  \$v5689\ := \$ram_lock\;
                  if \$v5689\(0) = '1' then
                    state_var5920 := Q_WAIT5688;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19234_sp\, X"000" & X"1")));
                    state_var5920 := PAUSE_GET5687;
                  end if;
                else
                  \$v5695\ := \$ram_lock\;
                  if \$v5695\(0) = '1' then
                    state_var5920 := Q_WAIT5694;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19238_w6514383_arg\(8 to 23), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5693;
                  end if;
                end if;
              when \$19252_FOREVER6704384\ =>
                \$19252_forever6704384_arg\ := eclat_unit;
                state_var5920 := \$19252_FOREVER6704384\;
              when \$19262_FOREVER6704385\ =>
                \$19262_forever6704385_arg\ := eclat_unit;
                state_var5920 := \$19262_FOREVER6704385\;
              when \$19320_FOREVER6704386\ =>
                \$19320_forever6704386_arg\ := eclat_unit;
                state_var5920 := \$19320_FOREVER6704386\;
              when \$19326_COMPBRANCH6504387\ =>
                \$19330_compare6444359_id\ := "000010100010";
                \$19330_compare6444359_arg\ := \$19326_compbranch6504387_arg\(0 to 31) & \$19326_compbranch6504387_arg\(32 to 62) & \$19326_compbranch6504387_arg\(110 to 140);
                state_var5920 := \$19330_COMPARE6444359\;
              when \$19330_COMPARE6444359\ =>
                \$v5824\ := \$19330_compare6444359_arg\(0 to 31);
                case \$v5824\ is
                when X"0000000" & X"0" =>
                  \$19330_compare6444359_result\ := work.Int.eq(\$19330_compare6444359_arg\(32 to 62), \$19330_compare6444359_arg\(63 to 93));
                when X"0000000" & X"1" =>
                  \$19330_compare6444359_result\ := work.Bool.lnot(work.Int.eq(
                                                                   \$19330_compare6444359_arg\(32 to 62), \$19330_compare6444359_arg\(63 to 93)));
                when X"0000000" & X"2" =>
                  \$19330_compare6444359_result\ := work.Int.lt(\$19330_compare6444359_arg\(32 to 62), \$19330_compare6444359_arg\(63 to 93));
                when X"0000000" & X"3" =>
                  \$19330_compare6444359_result\ := eclat_if(work.Int.lt(
                                                             \$19330_compare6444359_arg\(32 to 62), \$19330_compare6444359_arg\(63 to 93)) & eclat_true & 
                                                    work.Int.eq(\$19330_compare6444359_arg\(32 to 62), \$19330_compare6444359_arg\(63 to 93)));
                when X"0000000" & X"4" =>
                  \$19330_compare6444359_result\ := work.Bool.lnot(eclat_if(
                                                                   work.Int.lt(
                                                                   \$19330_compare6444359_arg\(32 to 62), \$19330_compare6444359_arg\(63 to 93)) & eclat_true & 
                                                                   work.Int.eq(
                                                                   \$19330_compare6444359_arg\(32 to 62), \$19330_compare6444359_arg\(63 to 93))));
                when X"0000000" & X"5" =>
                  \$19330_compare6444359_result\ := work.Bool.lnot(work.Int.lt(
                                                                   \$19330_compare6444359_arg\(32 to 62), \$19330_compare6444359_arg\(63 to 93)));
                when others =>
                  \$19330_compare6444359_result\ := eclat_false;
                end case;
                \$19329_b\ := \$19330_compare6444359_result\;
                \$19326_compbranch6504387_result\ := eclat_if(\$19329_b\ & 
                                                     work.Int.add(work.Int.add(
                                                                  \$19326_compbranch6504387_arg\(94 to 109), X"000" & X"2"), eclat_resize(\$19326_compbranch6504387_arg\(63 to 93),16)) & \$19326_compbranch6504387_arg\(110 to 141) & \$19326_compbranch6504387_arg\(142 to 157) & \$19326_compbranch6504387_arg\(158 to 213) & \$19326_compbranch6504387_arg\(214 to 215) & 
                                                     work.Int.add(\$19326_compbranch6504387_arg\(94 to 109), X"000" & X"3") & \$19326_compbranch6504387_arg\(110 to 141) & \$19326_compbranch6504387_arg\(142 to 157) & \$19326_compbranch6504387_arg\(158 to 213) & \$19326_compbranch6504387_arg\(214 to 215));
                result4928 := \$19326_compbranch6504387_result\;
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when \$19333_COMPBRANCH6504388\ =>
                \$19337_compare6444359_id\ := "000010100100";
                \$19337_compare6444359_arg\ := \$19333_compbranch6504388_arg\(0 to 31) & \$19333_compbranch6504388_arg\(32 to 62) & \$19333_compbranch6504388_arg\(110 to 140);
                state_var5920 := \$19337_COMPARE6444359\;
              when \$19337_COMPARE6444359\ =>
                \$v5825\ := \$19337_compare6444359_arg\(0 to 31);
                case \$v5825\ is
                when X"0000000" & X"0" =>
                  \$19337_compare6444359_result\ := work.Int.eq(\$19337_compare6444359_arg\(32 to 62), \$19337_compare6444359_arg\(63 to 93));
                when X"0000000" & X"1" =>
                  \$19337_compare6444359_result\ := work.Bool.lnot(work.Int.eq(
                                                                   \$19337_compare6444359_arg\(32 to 62), \$19337_compare6444359_arg\(63 to 93)));
                when X"0000000" & X"2" =>
                  \$19337_compare6444359_result\ := work.Int.lt(\$19337_compare6444359_arg\(32 to 62), \$19337_compare6444359_arg\(63 to 93));
                when X"0000000" & X"3" =>
                  \$19337_compare6444359_result\ := eclat_if(work.Int.lt(
                                                             \$19337_compare6444359_arg\(32 to 62), \$19337_compare6444359_arg\(63 to 93)) & eclat_true & 
                                                    work.Int.eq(\$19337_compare6444359_arg\(32 to 62), \$19337_compare6444359_arg\(63 to 93)));
                when X"0000000" & X"4" =>
                  \$19337_compare6444359_result\ := work.Bool.lnot(eclat_if(
                                                                   work.Int.lt(
                                                                   \$19337_compare6444359_arg\(32 to 62), \$19337_compare6444359_arg\(63 to 93)) & eclat_true & 
                                                                   work.Int.eq(
                                                                   \$19337_compare6444359_arg\(32 to 62), \$19337_compare6444359_arg\(63 to 93))));
                when X"0000000" & X"5" =>
                  \$19337_compare6444359_result\ := work.Bool.lnot(work.Int.lt(
                                                                   \$19337_compare6444359_arg\(32 to 62), \$19337_compare6444359_arg\(63 to 93)));
                when others =>
                  \$19337_compare6444359_result\ := eclat_false;
                end case;
                \$19336_b\ := \$19337_compare6444359_result\;
                \$19333_compbranch6504388_result\ := eclat_if(\$19336_b\ & 
                                                     work.Int.add(work.Int.add(
                                                                  \$19333_compbranch6504388_arg\(94 to 109), X"000" & X"2"), eclat_resize(\$19333_compbranch6504388_arg\(63 to 93),16)) & \$19333_compbranch6504388_arg\(110 to 141) & \$19333_compbranch6504388_arg\(142 to 157) & \$19333_compbranch6504388_arg\(158 to 213) & \$19333_compbranch6504388_arg\(214 to 215) & 
                                                     work.Int.add(\$19333_compbranch6504388_arg\(94 to 109), X"000" & X"3") & \$19333_compbranch6504388_arg\(110 to 141) & \$19333_compbranch6504388_arg\(142 to 157) & \$19333_compbranch6504388_arg\(158 to 213) & \$19333_compbranch6504388_arg\(214 to 215));
                result4928 := \$19333_compbranch6504388_result\;
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when \$19347_FILL6534389\ =>
                \$v5835\ := work.Int.gt(\$19347_fill6534389_arg\(0 to 15), \$19347_fill6534389_arg\(32 to 47));
                if \$v5835\(0) = '1' then
                  \$19347_fill6534389_result\ := \$19347_fill6534389_arg\(16 to 31);
                  \$19346_sp\ := \$19347_fill6534389_result\;
                  result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"3") & \$19344\(64 to 95) & \$19346_sp\ & \$19344\(32 to 63) & \$18788\(96 to 103) & \$18788\(104 to 119) & \$18788\(120 to 121);
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$v5834\ := \$ram_lock\;
                  if \$v5834\(0) = '1' then
                    state_var5920 := Q_WAIT5833;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19347_fill6534389_arg\(16 to 31), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5832;
                  end if;
                end if;
              when \$19361_FILL6544390\ =>
                \$v5864\ := work.Int.ge(\$19361_fill6544390_arg\(0 to 15), \$19361_fill6544390_arg\(32 to 47));
                if \$v5864\(0) = '1' then
                  \$19361_fill6544390_result\ := \$19361_fill6544390_arg\(16 to 31);
                  \$19360_sp\ := \$19361_fill6544390_result\;
                  result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"3") & \$19358\(64 to 95) & \$19360_sp\ & \$19358\(32 to 63) & \$18788\(96 to 103) & \$18788\(104 to 119) & \$18788\(120 to 121);
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$v5863\ := \$ram_lock\;
                  if \$v5863\(0) = '1' then
                    state_var5920 := Q_WAIT5862;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19361_fill6544390_arg\(16 to 31), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5861;
                  end if;
                end if;
              when \$19366_COMPBRANCH6504391\ =>
                \$19370_compare6444359_id\ := "000010101011";
                \$19370_compare6444359_arg\ := \$19366_compbranch6504391_arg\(0 to 31) & \$19366_compbranch6504391_arg\(32 to 62) & \$19366_compbranch6504391_arg\(110 to 140);
                state_var5920 := \$19370_COMPARE6444359\;
              when \$19370_COMPARE6444359\ =>
                \$v5868\ := \$19370_compare6444359_arg\(0 to 31);
                case \$v5868\ is
                when X"0000000" & X"0" =>
                  \$19370_compare6444359_result\ := work.Int.eq(\$19370_compare6444359_arg\(32 to 62), \$19370_compare6444359_arg\(63 to 93));
                when X"0000000" & X"1" =>
                  \$19370_compare6444359_result\ := work.Bool.lnot(work.Int.eq(
                                                                   \$19370_compare6444359_arg\(32 to 62), \$19370_compare6444359_arg\(63 to 93)));
                when X"0000000" & X"2" =>
                  \$19370_compare6444359_result\ := work.Int.lt(\$19370_compare6444359_arg\(32 to 62), \$19370_compare6444359_arg\(63 to 93));
                when X"0000000" & X"3" =>
                  \$19370_compare6444359_result\ := eclat_if(work.Int.lt(
                                                             \$19370_compare6444359_arg\(32 to 62), \$19370_compare6444359_arg\(63 to 93)) & eclat_true & 
                                                    work.Int.eq(\$19370_compare6444359_arg\(32 to 62), \$19370_compare6444359_arg\(63 to 93)));
                when X"0000000" & X"4" =>
                  \$19370_compare6444359_result\ := work.Bool.lnot(eclat_if(
                                                                   work.Int.lt(
                                                                   \$19370_compare6444359_arg\(32 to 62), \$19370_compare6444359_arg\(63 to 93)) & eclat_true & 
                                                                   work.Int.eq(
                                                                   \$19370_compare6444359_arg\(32 to 62), \$19370_compare6444359_arg\(63 to 93))));
                when X"0000000" & X"5" =>
                  \$19370_compare6444359_result\ := work.Bool.lnot(work.Int.lt(
                                                                   \$19370_compare6444359_arg\(32 to 62), \$19370_compare6444359_arg\(63 to 93)));
                when others =>
                  \$19370_compare6444359_result\ := eclat_false;
                end case;
                \$19369_b\ := \$19370_compare6444359_result\;
                \$19366_compbranch6504391_result\ := eclat_if(\$19369_b\ & 
                                                     work.Int.add(work.Int.add(
                                                                  \$19366_compbranch6504391_arg\(94 to 109), X"000" & X"2"), eclat_resize(\$19366_compbranch6504391_arg\(63 to 93),16)) & \$19366_compbranch6504391_arg\(110 to 141) & \$19366_compbranch6504391_arg\(142 to 157) & \$19366_compbranch6504391_arg\(158 to 213) & \$19366_compbranch6504391_arg\(214 to 215) & 
                                                     work.Int.add(\$19366_compbranch6504391_arg\(94 to 109), X"000" & X"3") & \$19366_compbranch6504391_arg\(110 to 141) & \$19366_compbranch6504391_arg\(142 to 157) & \$19366_compbranch6504391_arg\(158 to 213) & \$19366_compbranch6504391_arg\(214 to 215));
                result4928 := \$19366_compbranch6504391_result\;
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when \$19373_COMPBRANCH6504392\ =>
                \$19377_compare6444359_id\ := "000010101101";
                \$19377_compare6444359_arg\ := \$19373_compbranch6504392_arg\(0 to 31) & \$19373_compbranch6504392_arg\(32 to 62) & \$19373_compbranch6504392_arg\(110 to 140);
                state_var5920 := \$19377_COMPARE6444359\;
              when \$19377_COMPARE6444359\ =>
                \$v5869\ := \$19377_compare6444359_arg\(0 to 31);
                case \$v5869\ is
                when X"0000000" & X"0" =>
                  \$19377_compare6444359_result\ := work.Int.eq(\$19377_compare6444359_arg\(32 to 62), \$19377_compare6444359_arg\(63 to 93));
                when X"0000000" & X"1" =>
                  \$19377_compare6444359_result\ := work.Bool.lnot(work.Int.eq(
                                                                   \$19377_compare6444359_arg\(32 to 62), \$19377_compare6444359_arg\(63 to 93)));
                when X"0000000" & X"2" =>
                  \$19377_compare6444359_result\ := work.Int.lt(\$19377_compare6444359_arg\(32 to 62), \$19377_compare6444359_arg\(63 to 93));
                when X"0000000" & X"3" =>
                  \$19377_compare6444359_result\ := eclat_if(work.Int.lt(
                                                             \$19377_compare6444359_arg\(32 to 62), \$19377_compare6444359_arg\(63 to 93)) & eclat_true & 
                                                    work.Int.eq(\$19377_compare6444359_arg\(32 to 62), \$19377_compare6444359_arg\(63 to 93)));
                when X"0000000" & X"4" =>
                  \$19377_compare6444359_result\ := work.Bool.lnot(eclat_if(
                                                                   work.Int.lt(
                                                                   \$19377_compare6444359_arg\(32 to 62), \$19377_compare6444359_arg\(63 to 93)) & eclat_true & 
                                                                   work.Int.eq(
                                                                   \$19377_compare6444359_arg\(32 to 62), \$19377_compare6444359_arg\(63 to 93))));
                when X"0000000" & X"5" =>
                  \$19377_compare6444359_result\ := work.Bool.lnot(work.Int.lt(
                                                                   \$19377_compare6444359_arg\(32 to 62), \$19377_compare6444359_arg\(63 to 93)));
                when others =>
                  \$19377_compare6444359_result\ := eclat_false;
                end case;
                \$19376_b\ := \$19377_compare6444359_result\;
                \$19373_compbranch6504392_result\ := eclat_if(\$19376_b\ & 
                                                     work.Int.add(work.Int.add(
                                                                  \$19373_compbranch6504392_arg\(94 to 109), X"000" & X"2"), eclat_resize(\$19373_compbranch6504392_arg\(63 to 93),16)) & \$19373_compbranch6504392_arg\(110 to 141) & \$19373_compbranch6504392_arg\(142 to 157) & \$19373_compbranch6504392_arg\(158 to 213) & \$19373_compbranch6504392_arg\(214 to 215) & 
                                                     work.Int.add(\$19373_compbranch6504392_arg\(94 to 109), X"000" & X"3") & \$19373_compbranch6504392_arg\(110 to 141) & \$19373_compbranch6504392_arg\(142 to 157) & \$19373_compbranch6504392_arg\(158 to 213) & \$19373_compbranch6504392_arg\(214 to 215));
                result4928 := \$19373_compbranch6504392_result\;
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when \$19380_COMPBRANCH6504393\ =>
                \$19384_compare6444359_id\ := "000010101111";
                \$19384_compare6444359_arg\ := \$19380_compbranch6504393_arg\(0 to 31) & \$19380_compbranch6504393_arg\(32 to 62) & \$19380_compbranch6504393_arg\(110 to 140);
                state_var5920 := \$19384_COMPARE6444359\;
              when \$19384_COMPARE6444359\ =>
                \$v5870\ := \$19384_compare6444359_arg\(0 to 31);
                case \$v5870\ is
                when X"0000000" & X"0" =>
                  \$19384_compare6444359_result\ := work.Int.eq(\$19384_compare6444359_arg\(32 to 62), \$19384_compare6444359_arg\(63 to 93));
                when X"0000000" & X"1" =>
                  \$19384_compare6444359_result\ := work.Bool.lnot(work.Int.eq(
                                                                   \$19384_compare6444359_arg\(32 to 62), \$19384_compare6444359_arg\(63 to 93)));
                when X"0000000" & X"2" =>
                  \$19384_compare6444359_result\ := work.Int.lt(\$19384_compare6444359_arg\(32 to 62), \$19384_compare6444359_arg\(63 to 93));
                when X"0000000" & X"3" =>
                  \$19384_compare6444359_result\ := eclat_if(work.Int.lt(
                                                             \$19384_compare6444359_arg\(32 to 62), \$19384_compare6444359_arg\(63 to 93)) & eclat_true & 
                                                    work.Int.eq(\$19384_compare6444359_arg\(32 to 62), \$19384_compare6444359_arg\(63 to 93)));
                when X"0000000" & X"4" =>
                  \$19384_compare6444359_result\ := work.Bool.lnot(eclat_if(
                                                                   work.Int.lt(
                                                                   \$19384_compare6444359_arg\(32 to 62), \$19384_compare6444359_arg\(63 to 93)) & eclat_true & 
                                                                   work.Int.eq(
                                                                   \$19384_compare6444359_arg\(32 to 62), \$19384_compare6444359_arg\(63 to 93))));
                when X"0000000" & X"5" =>
                  \$19384_compare6444359_result\ := work.Bool.lnot(work.Int.lt(
                                                                   \$19384_compare6444359_arg\(32 to 62), \$19384_compare6444359_arg\(63 to 93)));
                when others =>
                  \$19384_compare6444359_result\ := eclat_false;
                end case;
                \$19383_b\ := \$19384_compare6444359_result\;
                \$19380_compbranch6504393_result\ := eclat_if(\$19383_b\ & 
                                                     work.Int.add(work.Int.add(
                                                                  \$19380_compbranch6504393_arg\(94 to 109), X"000" & X"2"), eclat_resize(\$19380_compbranch6504393_arg\(63 to 93),16)) & \$19380_compbranch6504393_arg\(110 to 141) & \$19380_compbranch6504393_arg\(142 to 157) & \$19380_compbranch6504393_arg\(158 to 213) & \$19380_compbranch6504393_arg\(214 to 215) & 
                                                     work.Int.add(\$19380_compbranch6504393_arg\(94 to 109), X"000" & X"3") & \$19380_compbranch6504393_arg\(110 to 141) & \$19380_compbranch6504393_arg\(142 to 157) & \$19380_compbranch6504393_arg\(158 to 213) & \$19380_compbranch6504393_arg\(214 to 215));
                result4928 := \$19380_compbranch6504393_result\;
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when \$19387_COMPBRANCH6504394\ =>
                \$19391_compare6444359_id\ := "000010110001";
                \$19391_compare6444359_arg\ := \$19387_compbranch6504394_arg\(0 to 31) & \$19387_compbranch6504394_arg\(32 to 62) & \$19387_compbranch6504394_arg\(110 to 140);
                state_var5920 := \$19391_COMPARE6444359\;
              when \$19391_COMPARE6444359\ =>
                \$v5871\ := \$19391_compare6444359_arg\(0 to 31);
                case \$v5871\ is
                when X"0000000" & X"0" =>
                  \$19391_compare6444359_result\ := work.Int.eq(\$19391_compare6444359_arg\(32 to 62), \$19391_compare6444359_arg\(63 to 93));
                when X"0000000" & X"1" =>
                  \$19391_compare6444359_result\ := work.Bool.lnot(work.Int.eq(
                                                                   \$19391_compare6444359_arg\(32 to 62), \$19391_compare6444359_arg\(63 to 93)));
                when X"0000000" & X"2" =>
                  \$19391_compare6444359_result\ := work.Int.lt(\$19391_compare6444359_arg\(32 to 62), \$19391_compare6444359_arg\(63 to 93));
                when X"0000000" & X"3" =>
                  \$19391_compare6444359_result\ := eclat_if(work.Int.lt(
                                                             \$19391_compare6444359_arg\(32 to 62), \$19391_compare6444359_arg\(63 to 93)) & eclat_true & 
                                                    work.Int.eq(\$19391_compare6444359_arg\(32 to 62), \$19391_compare6444359_arg\(63 to 93)));
                when X"0000000" & X"4" =>
                  \$19391_compare6444359_result\ := work.Bool.lnot(eclat_if(
                                                                   work.Int.lt(
                                                                   \$19391_compare6444359_arg\(32 to 62), \$19391_compare6444359_arg\(63 to 93)) & eclat_true & 
                                                                   work.Int.eq(
                                                                   \$19391_compare6444359_arg\(32 to 62), \$19391_compare6444359_arg\(63 to 93))));
                when X"0000000" & X"5" =>
                  \$19391_compare6444359_result\ := work.Bool.lnot(work.Int.lt(
                                                                   \$19391_compare6444359_arg\(32 to 62), \$19391_compare6444359_arg\(63 to 93)));
                when others =>
                  \$19391_compare6444359_result\ := eclat_false;
                end case;
                \$19390_b\ := \$19391_compare6444359_result\;
                \$19387_compbranch6504394_result\ := eclat_if(\$19390_b\ & 
                                                     work.Int.add(work.Int.add(
                                                                  \$19387_compbranch6504394_arg\(94 to 109), X"000" & X"2"), eclat_resize(\$19387_compbranch6504394_arg\(63 to 93),16)) & \$19387_compbranch6504394_arg\(110 to 141) & \$19387_compbranch6504394_arg\(142 to 157) & \$19387_compbranch6504394_arg\(158 to 213) & \$19387_compbranch6504394_arg\(214 to 215) & 
                                                     work.Int.add(\$19387_compbranch6504394_arg\(94 to 109), X"000" & X"3") & \$19387_compbranch6504394_arg\(110 to 141) & \$19387_compbranch6504394_arg\(142 to 157) & \$19387_compbranch6504394_arg\(158 to 213) & \$19387_compbranch6504394_arg\(214 to 215));
                result4928 := \$19387_compbranch6504394_result\;
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when \$19394_COMPBRANCH6504395\ =>
                \$19398_compare6444359_id\ := "000010110011";
                \$19398_compare6444359_arg\ := \$19394_compbranch6504395_arg\(0 to 31) & \$19394_compbranch6504395_arg\(32 to 62) & \$19394_compbranch6504395_arg\(110 to 140);
                state_var5920 := \$19398_COMPARE6444359\;
              when \$19398_COMPARE6444359\ =>
                \$v5872\ := \$19398_compare6444359_arg\(0 to 31);
                case \$v5872\ is
                when X"0000000" & X"0" =>
                  \$19398_compare6444359_result\ := work.Int.eq(\$19398_compare6444359_arg\(32 to 62), \$19398_compare6444359_arg\(63 to 93));
                when X"0000000" & X"1" =>
                  \$19398_compare6444359_result\ := work.Bool.lnot(work.Int.eq(
                                                                   \$19398_compare6444359_arg\(32 to 62), \$19398_compare6444359_arg\(63 to 93)));
                when X"0000000" & X"2" =>
                  \$19398_compare6444359_result\ := work.Int.lt(\$19398_compare6444359_arg\(32 to 62), \$19398_compare6444359_arg\(63 to 93));
                when X"0000000" & X"3" =>
                  \$19398_compare6444359_result\ := eclat_if(work.Int.lt(
                                                             \$19398_compare6444359_arg\(32 to 62), \$19398_compare6444359_arg\(63 to 93)) & eclat_true & 
                                                    work.Int.eq(\$19398_compare6444359_arg\(32 to 62), \$19398_compare6444359_arg\(63 to 93)));
                when X"0000000" & X"4" =>
                  \$19398_compare6444359_result\ := work.Bool.lnot(eclat_if(
                                                                   work.Int.lt(
                                                                   \$19398_compare6444359_arg\(32 to 62), \$19398_compare6444359_arg\(63 to 93)) & eclat_true & 
                                                                   work.Int.eq(
                                                                   \$19398_compare6444359_arg\(32 to 62), \$19398_compare6444359_arg\(63 to 93))));
                when X"0000000" & X"5" =>
                  \$19398_compare6444359_result\ := work.Bool.lnot(work.Int.lt(
                                                                   \$19398_compare6444359_arg\(32 to 62), \$19398_compare6444359_arg\(63 to 93)));
                when others =>
                  \$19398_compare6444359_result\ := eclat_false;
                end case;
                \$19397_b\ := \$19398_compare6444359_result\;
                \$19394_compbranch6504395_result\ := eclat_if(\$19397_b\ & 
                                                     work.Int.add(work.Int.add(
                                                                  \$19394_compbranch6504395_arg\(94 to 109), X"000" & X"2"), eclat_resize(\$19394_compbranch6504395_arg\(63 to 93),16)) & \$19394_compbranch6504395_arg\(110 to 141) & \$19394_compbranch6504395_arg\(142 to 157) & \$19394_compbranch6504395_arg\(158 to 213) & \$19394_compbranch6504395_arg\(214 to 215) & 
                                                     work.Int.add(\$19394_compbranch6504395_arg\(94 to 109), X"000" & X"3") & \$19394_compbranch6504395_arg\(110 to 141) & \$19394_compbranch6504395_arg\(142 to 157) & \$19394_compbranch6504395_arg\(158 to 213) & \$19394_compbranch6504395_arg\(214 to 215));
                result4928 := \$19394_compbranch6504395_result\;
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when \$19401_COMPBRANCH6504396\ =>
                \$19405_compare6444359_id\ := "000010110101";
                \$19405_compare6444359_arg\ := \$19401_compbranch6504396_arg\(0 to 31) & \$19401_compbranch6504396_arg\(32 to 62) & \$19401_compbranch6504396_arg\(110 to 140);
                state_var5920 := \$19405_COMPARE6444359\;
              when \$19405_COMPARE6444359\ =>
                \$v5873\ := \$19405_compare6444359_arg\(0 to 31);
                case \$v5873\ is
                when X"0000000" & X"0" =>
                  \$19405_compare6444359_result\ := work.Int.eq(\$19405_compare6444359_arg\(32 to 62), \$19405_compare6444359_arg\(63 to 93));
                when X"0000000" & X"1" =>
                  \$19405_compare6444359_result\ := work.Bool.lnot(work.Int.eq(
                                                                   \$19405_compare6444359_arg\(32 to 62), \$19405_compare6444359_arg\(63 to 93)));
                when X"0000000" & X"2" =>
                  \$19405_compare6444359_result\ := work.Int.lt(\$19405_compare6444359_arg\(32 to 62), \$19405_compare6444359_arg\(63 to 93));
                when X"0000000" & X"3" =>
                  \$19405_compare6444359_result\ := eclat_if(work.Int.lt(
                                                             \$19405_compare6444359_arg\(32 to 62), \$19405_compare6444359_arg\(63 to 93)) & eclat_true & 
                                                    work.Int.eq(\$19405_compare6444359_arg\(32 to 62), \$19405_compare6444359_arg\(63 to 93)));
                when X"0000000" & X"4" =>
                  \$19405_compare6444359_result\ := work.Bool.lnot(eclat_if(
                                                                   work.Int.lt(
                                                                   \$19405_compare6444359_arg\(32 to 62), \$19405_compare6444359_arg\(63 to 93)) & eclat_true & 
                                                                   work.Int.eq(
                                                                   \$19405_compare6444359_arg\(32 to 62), \$19405_compare6444359_arg\(63 to 93))));
                when X"0000000" & X"5" =>
                  \$19405_compare6444359_result\ := work.Bool.lnot(work.Int.lt(
                                                                   \$19405_compare6444359_arg\(32 to 62), \$19405_compare6444359_arg\(63 to 93)));
                when others =>
                  \$19405_compare6444359_result\ := eclat_false;
                end case;
                \$19404_b\ := \$19405_compare6444359_result\;
                \$19401_compbranch6504396_result\ := eclat_if(\$19404_b\ & 
                                                     work.Int.add(work.Int.add(
                                                                  \$19401_compbranch6504396_arg\(94 to 109), X"000" & X"2"), eclat_resize(\$19401_compbranch6504396_arg\(63 to 93),16)) & \$19401_compbranch6504396_arg\(110 to 141) & \$19401_compbranch6504396_arg\(142 to 157) & \$19401_compbranch6504396_arg\(158 to 213) & \$19401_compbranch6504396_arg\(214 to 215) & 
                                                     work.Int.add(\$19401_compbranch6504396_arg\(94 to 109), X"000" & X"3") & \$19401_compbranch6504396_arg\(110 to 141) & \$19401_compbranch6504396_arg\(142 to 157) & \$19401_compbranch6504396_arg\(158 to 213) & \$19401_compbranch6504396_arg\(214 to 215));
                result4928 := \$19401_compbranch6504396_result\;
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when \$19416_W36574398\ =>
                \$v5877\ := work.Int.ge(\$19416_w36574398_arg\(0 to 15), \$19416_w36574398_arg\(32 to 47));
                if \$v5877\(0) = '1' then
                  \$19416_w36574398_result\ := \$19416_w36574398_arg\(16 to 31);
                  \$19415_sp\ := \$19416_w36574398_result\;
                  result4928 := work.Int.add(work.Int.add(\$18788\(0 to 15), X"000" & X"3"), eclat_resize(\$19215_argument1\,16)) & \$19410\(64 to 95) & \$19415_sp\ & \$19410\(32 to 63) & \$18788\(96 to 103) & \$18788\(104 to 119) & \$18788\(120 to 121);
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                else
                  \$v5876\ := \$ram_lock\;
                  if \$v5876\(0) = '1' then
                    state_var5920 := Q_WAIT5875;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19416_w36574398_arg\(16 to 31)));
                    \$ram_write\ <= eclat_resize(work.Int.add(eclat_resize(\$19416_w36574398_arg\(48 to 78),16), 
                                                              work.Int.mul(
                                                              X"000" & X"2", \$19416_w36574398_arg\(0 to 15))),31) & eclat_true; \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5874;
                  end if;
                end if;
              when \$19420_W06554397\ =>
                \$v5887\ := work.Int.ge(\$19420_w06554397_arg\(0 to 15), \$19420_w06554397_arg\(48 to 63));
                if \$v5887\(0) = '1' then
                  \$19420_w06554397_result\ := \$19420_w06554397_arg\(16 to 31);
                  \$19412_sp\ := \$19420_w06554397_result\;
                  \$18799_w1656_id\ := "000010111000";
                  \$18799_w1656_arg\ := X"000" & X"1" & \$18788\(0 to 15) & eclat_resize(\$19215_argument1\,16) & \$19410\(64 to 95);
                  state_var5920 := \$18799_W1656\;
                else
                  \$v5886\ := \$ram_lock\;
                  if \$v5886\(0) = '1' then
                    state_var5920 := Q_WAIT5885;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19420_w06554397_arg\(16 to 31), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5884;
                  end if;
                end if;
              when PAUSE_GET4934 =>
                \$19761\ := \$ram_value\;
                release(\$ram_lock\);
                \$v4933\ := \$ram_lock\;
                if \$v4933\(0) = '1' then
                  state_var5920 := Q_WAIT4932;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$18790_loop666_arg\(16 to 31), \$18790_loop666_arg\(0 to 15))));
                  \$ram_write\ <= \$19761\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET4931;
                end if;
              when PAUSE_GET4950 =>
                \$19745_hd\ := \$ram_value\;
                release(\$ram_lock\);
                \$19746\ := work.Print.print_string(clk,of_string("bloc "));
                \$19747\ := work.Int.print(clk,eclat_resize(\$19741\(0 to 30),16));
                \$19748\ := work.Print.print_string(clk,of_string(" of size "));
                \$19749\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                            work.Int.lsr(
                                                            \$19745_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$19750\ := work.Print.print_string(clk,of_string(" from "));
                \$19751\ := work.Int.print(clk,eclat_resize(\$19741\(0 to 30),16));
                \$19752\ := work.Print.print_string(clk,of_string(" to "));
                \$19753\ := work.Int.print(clk,\$18791_loop665_arg\(16 to 31));
                \$19754\ := work.Print.print_newline(clk,eclat_unit);
                \$v4949\ := \$ram_lock\;
                if \$v4949\(0) = '1' then
                  state_var5920 := Q_WAIT4948;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18791_loop665_arg\(16 to 31)));
                  \$ram_write\ <= \$19745_hd\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET4947;
                end if;
              when PAUSE_GET4954 =>
                \$19744_w\ := \$ram_value\;
                release(\$ram_lock\);
                \$v4953\ := eclat_if(work.Bool.lnot(""&\$19744_w\(31)) & 
                            eclat_if(work.Int.le(\$18791_loop665_arg\(48 to 63), eclat_resize(\$19744_w\(0 to 30),16)) & 
                            work.Int.lt(eclat_resize(\$19744_w\(0 to 30),16), 
                                        work.Int.add(\$18791_loop665_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false);
                if \$v4953\(0) = '1' then
                  \$19742\ := \$19744_w\ & \$18791_loop665_arg\(16 to 31);
                  \$v4940\ := \$ram_lock\;
                  if \$v4940\(0) = '1' then
                    state_var5920 := Q_WAIT4939;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            \$18791_loop665_arg\(64 to 79), \$18791_loop665_arg\(0 to 15))));
                    \$ram_write\ <= \$19742\(0 to 31); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET4938;
                  end if;
                else
                  \$v4952\ := \$ram_lock\;
                  if \$v4952\(0) = '1' then
                    state_var5920 := Q_WAIT4951;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$19741\(0 to 30),16)));
                    state_var5920 := PAUSE_GET4950;
                  end if;
                end if;
              when PAUSE_GET4958 =>
                \$19741\ := \$ram_value\;
                release(\$ram_lock\);
                \$v4957\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$19741\(31)) & 
                                           eclat_if(work.Int.le(\$18791_loop665_arg\(32 to 47), eclat_resize(\$19741\(0 to 30),16)) & 
                                           work.Int.lt(eclat_resize(\$19741\(0 to 30),16), 
                                                       work.Int.add(\$18791_loop665_arg\(32 to 47), X"1770")) & eclat_false) & eclat_false));
                if \$v4957\(0) = '1' then
                  \$19742\ := \$19741\ & \$18791_loop665_arg\(16 to 31);
                  \$v4940\ := \$ram_lock\;
                  if \$v4940\(0) = '1' then
                    state_var5920 := Q_WAIT4939;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            \$18791_loop665_arg\(64 to 79), \$18791_loop665_arg\(0 to 15))));
                    \$ram_write\ <= \$19742\(0 to 31); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET4938;
                  end if;
                else
                  \$v4956\ := \$ram_lock\;
                  if \$v4956\(0) = '1' then
                    state_var5920 := Q_WAIT4955;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19741\(0 to 30),16), X"000" & X"1")));
                    state_var5920 := PAUSE_GET4954;
                  end if;
                end if;
              when PAUSE_GET5175 =>
                \$19469\ := \$ram_value\;
                release(\$ram_lock\);
                \$18794_apply638_result\ := eclat_resize(\$19469\(0 to 30),16) & \$18794_apply638_arg\(60 to 91) & \$19468_sp\ & \$18794_apply638_arg\(60 to 91) & \$18794_apply638_arg\(3 to 10) & \$18794_apply638_arg\(150 to 165) & \$18794_apply638_arg\(108 to 109);
                result4928 := \$18794_apply638_result\;
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5200 =>
                \$19476_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$19464\ := \$19476_v\ & work.Int.sub(\$19463\(32 to 47), X"000" & X"1");
                \$v5199\ := ""&\$18794_apply638_arg\(11);
                if \$v5199\(0) = '1' then
                  \$19465_sp\ := work.Int.add(work.Int.sub(\$19464\(32 to 47), \$18794_apply638_arg\(12 to 27)), \$18794_apply638_arg\(28 to 43));
                  \$v5189\ := ""&\$18794_apply638_arg\(2);
                  if \$v5189\(0) = '1' then
                    \$v5188\ := \$ram_lock\;
                    if \$v5188\(0) = '1' then
                      state_var5920 := Q_WAIT5187;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(\$19465_sp\));
                      \$ram_write\ <= \$19464\(0 to 31); \$ram_write_request\ <= '1';
                      state_var5920 := PAUSE_SET5186;
                    end if;
                  else
                    \$19466_sp\ := \$19465_sp\;
                    \$v5185\ := ""&\$18794_apply638_arg\(1);
                    if \$v5185\(0) = '1' then
                      \$v5184\ := \$ram_lock\;
                      if \$v5184\(0) = '1' then
                        state_var5920 := Q_WAIT5183;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr_write\ <= to_integer(unsigned(\$19466_sp\));
                        \$ram_write\ <= \$19463\(0 to 31); \$ram_write_request\ <= '1';
                        state_var5920 := PAUSE_SET5182;
                      end if;
                    else
                      \$19467_sp\ := \$19466_sp\;
                      \$v5181\ := ""&\$18794_apply638_arg\(0);
                      if \$v5181\(0) = '1' then
                        \$v5180\ := \$ram_lock\;
                        if \$v5180\(0) = '1' then
                          state_var5920 := Q_WAIT5179;
                        else
                          acquire(\$ram_lock\);
                          \$ram_ptr_write\ <= to_integer(unsigned(\$19467_sp\));
                          \$ram_write\ <= \$19462\(0 to 31); \$ram_write_request\ <= '1';
                          state_var5920 := PAUSE_SET5178;
                        end if;
                      else
                        \$19468_sp\ := \$19467_sp\;
                        \$v5177\ := \$ram_lock\;
                        if \$v5177\(0) = '1' then
                          state_var5920 := Q_WAIT5176;
                        else
                          acquire(\$ram_lock\);
                          \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                            work.Int.add(
                                                            eclat_resize(\$18794_apply638_arg\(60 to 90),16), X"000" & X"0"), X"000" & X"1")));
                          state_var5920 := PAUSE_GET5175;
                        end if;
                      end if;
                    end if;
                  end if;
                else
                  \$v5198\ := \$ram_lock\;
                  if \$v5198\(0) = '1' then
                    state_var5920 := Q_WAIT5197;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19464\(32 to 47)));
                    \$ram_write\ <= eclat_resize(\$18794_apply638_arg\(142 to 149),31) & eclat_true; \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5196;
                  end if;
                end if;
              when PAUSE_GET5204 =>
                \$19477_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$19463\ := \$19477_v\ & work.Int.sub(\$19462\(32 to 47), X"000" & X"1");
                \$v5203\ := ""&\$18794_apply638_arg\(2);
                if \$v5203\(0) = '1' then
                  \$v5202\ := \$ram_lock\;
                  if \$v5202\(0) = '1' then
                    state_var5920 := Q_WAIT5201;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19463\(32 to 47), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5200;
                  end if;
                else
                  \$19464\ := "000"& X"000000" & X"1" & eclat_true & \$19463\(32 to 47);
                  \$v5199\ := ""&\$18794_apply638_arg\(11);
                  if \$v5199\(0) = '1' then
                    \$19465_sp\ := work.Int.add(work.Int.sub(\$19464\(32 to 47), \$18794_apply638_arg\(12 to 27)), \$18794_apply638_arg\(28 to 43));
                    \$v5189\ := ""&\$18794_apply638_arg\(2);
                    if \$v5189\(0) = '1' then
                      \$v5188\ := \$ram_lock\;
                      if \$v5188\(0) = '1' then
                        state_var5920 := Q_WAIT5187;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr_write\ <= to_integer(unsigned(\$19465_sp\));
                        \$ram_write\ <= \$19464\(0 to 31); \$ram_write_request\ <= '1';
                        state_var5920 := PAUSE_SET5186;
                      end if;
                    else
                      \$19466_sp\ := \$19465_sp\;
                      \$v5185\ := ""&\$18794_apply638_arg\(1);
                      if \$v5185\(0) = '1' then
                        \$v5184\ := \$ram_lock\;
                        if \$v5184\(0) = '1' then
                          state_var5920 := Q_WAIT5183;
                        else
                          acquire(\$ram_lock\);
                          \$ram_ptr_write\ <= to_integer(unsigned(\$19466_sp\));
                          \$ram_write\ <= \$19463\(0 to 31); \$ram_write_request\ <= '1';
                          state_var5920 := PAUSE_SET5182;
                        end if;
                      else
                        \$19467_sp\ := \$19466_sp\;
                        \$v5181\ := ""&\$18794_apply638_arg\(0);
                        if \$v5181\(0) = '1' then
                          \$v5180\ := \$ram_lock\;
                          if \$v5180\(0) = '1' then
                            state_var5920 := Q_WAIT5179;
                          else
                            acquire(\$ram_lock\);
                            \$ram_ptr_write\ <= to_integer(unsigned(\$19467_sp\));
                            \$ram_write\ <= \$19462\(0 to 31); \$ram_write_request\ <= '1';
                            state_var5920 := PAUSE_SET5178;
                          end if;
                        else
                          \$19468_sp\ := \$19467_sp\;
                          \$v5177\ := \$ram_lock\;
                          if \$v5177\(0) = '1' then
                            state_var5920 := Q_WAIT5176;
                          else
                            acquire(\$ram_lock\);
                            \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                              work.Int.add(
                                                              eclat_resize(\$18794_apply638_arg\(60 to 90),16), X"000" & X"0"), X"000" & X"1")));
                            state_var5920 := PAUSE_GET5175;
                          end if;
                        end if;
                      end if;
                    end if;
                  else
                    \$v5198\ := \$ram_lock\;
                    if \$v5198\(0) = '1' then
                      state_var5920 := Q_WAIT5197;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(\$19464\(32 to 47)));
                      \$ram_write\ <= eclat_resize(\$18794_apply638_arg\(142 to 149),31) & eclat_true; \$ram_write_request\ <= '1';
                      state_var5920 := PAUSE_SET5196;
                    end if;
                  end if;
                end if;
              when PAUSE_GET5208 =>
                \$19478_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$19462\ := \$19478_v\ & work.Int.sub(\$18794_apply638_arg\(92 to 107), X"000" & X"1");
                \$v5207\ := ""&\$18794_apply638_arg\(1);
                if \$v5207\(0) = '1' then
                  \$v5206\ := \$ram_lock\;
                  if \$v5206\(0) = '1' then
                    state_var5920 := Q_WAIT5205;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19462\(32 to 47), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5204;
                  end if;
                else
                  \$19463\ := "000"& X"000000" & X"1" & eclat_true & \$19462\(32 to 47);
                  \$v5203\ := ""&\$18794_apply638_arg\(2);
                  if \$v5203\(0) = '1' then
                    \$v5202\ := \$ram_lock\;
                    if \$v5202\(0) = '1' then
                      state_var5920 := Q_WAIT5201;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(
                                                        \$19463\(32 to 47), X"000" & X"1")));
                      state_var5920 := PAUSE_GET5200;
                    end if;
                  else
                    \$19464\ := "000"& X"000000" & X"1" & eclat_true & \$19463\(32 to 47);
                    \$v5199\ := ""&\$18794_apply638_arg\(11);
                    if \$v5199\(0) = '1' then
                      \$19465_sp\ := work.Int.add(work.Int.sub(\$19464\(32 to 47), \$18794_apply638_arg\(12 to 27)), \$18794_apply638_arg\(28 to 43));
                      \$v5189\ := ""&\$18794_apply638_arg\(2);
                      if \$v5189\(0) = '1' then
                        \$v5188\ := \$ram_lock\;
                        if \$v5188\(0) = '1' then
                          state_var5920 := Q_WAIT5187;
                        else
                          acquire(\$ram_lock\);
                          \$ram_ptr_write\ <= to_integer(unsigned(\$19465_sp\));
                          \$ram_write\ <= \$19464\(0 to 31); \$ram_write_request\ <= '1';
                          state_var5920 := PAUSE_SET5186;
                        end if;
                      else
                        \$19466_sp\ := \$19465_sp\;
                        \$v5185\ := ""&\$18794_apply638_arg\(1);
                        if \$v5185\(0) = '1' then
                          \$v5184\ := \$ram_lock\;
                          if \$v5184\(0) = '1' then
                            state_var5920 := Q_WAIT5183;
                          else
                            acquire(\$ram_lock\);
                            \$ram_ptr_write\ <= to_integer(unsigned(\$19466_sp\));
                            \$ram_write\ <= \$19463\(0 to 31); \$ram_write_request\ <= '1';
                            state_var5920 := PAUSE_SET5182;
                          end if;
                        else
                          \$19467_sp\ := \$19466_sp\;
                          \$v5181\ := ""&\$18794_apply638_arg\(0);
                          if \$v5181\(0) = '1' then
                            \$v5180\ := \$ram_lock\;
                            if \$v5180\(0) = '1' then
                              state_var5920 := Q_WAIT5179;
                            else
                              acquire(\$ram_lock\);
                              \$ram_ptr_write\ <= to_integer(unsigned(\$19467_sp\));
                              \$ram_write\ <= \$19462\(0 to 31); \$ram_write_request\ <= '1';
                              state_var5920 := PAUSE_SET5178;
                            end if;
                          else
                            \$19468_sp\ := \$19467_sp\;
                            \$v5177\ := \$ram_lock\;
                            if \$v5177\(0) = '1' then
                              state_var5920 := Q_WAIT5176;
                            else
                              acquire(\$ram_lock\);
                              \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                                work.Int.add(
                                                                eclat_resize(\$18794_apply638_arg\(60 to 90),16), X"000" & X"0"), X"000" & X"1")));
                              state_var5920 := PAUSE_GET5175;
                            end if;
                          end if;
                        end if;
                      end if;
                    else
                      \$v5198\ := \$ram_lock\;
                      if \$v5198\(0) = '1' then
                        state_var5920 := Q_WAIT5197;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr_write\ <= to_integer(unsigned(\$19464\(32 to 47)));
                        \$ram_write\ <= eclat_resize(\$18794_apply638_arg\(142 to 149),31) & eclat_true; \$ram_write_request\ <= '1';
                        state_var5920 := PAUSE_SET5196;
                      end if;
                    end if;
                  end if;
                end if;
              when PAUSE_GET5216 =>
                \$19448_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5215\ := \$ram_lock\;
                if \$v5215\(0) = '1' then
                  state_var5920 := Q_WAIT5214;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$19444\(64 to 94),16), X"000" & X"2"), X"000" & X"1")));
                  \$ram_write\ <= \$19448_v\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5213;
                end if;
              when PAUSE_GET5223 =>
                \$19450_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5222\ := \$ram_lock\;
                if \$v5222\(0) = '1' then
                  state_var5920 := Q_WAIT5221;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$19444\(64 to 94),16), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= \$19450_v\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5220;
                end if;
              when PAUSE_GET5231 =>
                \$19441_arg\ := \$code_value\;
                release(\$code_lock\);
                \$18797_branch_if648_result\ := work.Int.add(work.Int.add(
                                                             \$18797_branch_if648_arg\(1 to 16), X"000" & X"1"), eclat_resize(\$19441_arg\,16)) & \$18797_branch_if648_arg\(17 to 48) & \$18797_branch_if648_arg\(49 to 64) & \$18797_branch_if648_arg\(65 to 120) & \$18797_branch_if648_arg\(121 to 122);
                result4928 := \$18797_branch_if648_result\;
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5238 =>
                \$19437\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5237\ := \$ram_lock\;
                if \$v5237\(0) = '1' then
                  state_var5920 := Q_WAIT5236;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.sub(
                                                          work.Int.sub(
                                                          work.Int.sub(
                                                          \$18798_w652_arg\(16 to 31), \$18798_w652_arg\(32 to 47)), \$18798_w652_arg\(48 to 63)), \$18798_w652_arg\(0 to 15))));
                  \$ram_write\ <= \$19437\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5235;
                end if;
              when PAUSE_GET5245 =>
                \$19433\ := \$code_value\;
                release(\$code_lock\);
                \$v5244\ := \$ram_lock\;
                if \$v5244\(0) = '1' then
                  state_var5920 := Q_WAIT5243;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$18799_w1656_arg\(48 to 78),16), 
                                                          work.Int.mul(
                                                          X"000" & X"2", \$18799_w1656_arg\(0 to 15))), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(work.Int.add(work.Int.add(
                                                            \$18799_w1656_arg\(16 to 31), X"000" & X"2"), eclat_resize(\$19433\,16)),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5242;
                end if;
              when PAUSE_GET5252 =>
                \$18817_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18817_v\ & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5255 =>
                \$18818_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18818_v\ & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5258 =>
                \$18819_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18819_v\ & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5261 =>
                \$18820_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18820_v\ & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5264 =>
                \$18821_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18821_v\ & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5267 =>
                \$18822_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18822_v\ & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5270 =>
                \$18823_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18823_v\ & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5273 =>
                \$18824_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18824_v\ & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5282 =>
                \$18828_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18828_v\ & 
                work.Int.add(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5288 =>
                \$18830_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18830_v\ & 
                work.Int.add(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5294 =>
                \$18832_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18832_v\ & 
                work.Int.add(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5300 =>
                \$18834_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18834_v\ & 
                work.Int.add(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5306 =>
                \$18836_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18836_v\ & 
                work.Int.add(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5312 =>
                \$18838_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18838_v\ & 
                work.Int.add(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5318 =>
                \$18840_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18840_v\ & 
                work.Int.add(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5324 =>
                \$18841\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18841\ & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5327 =>
                \$18842\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18842\ & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5330 =>
                \$18843\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18843\ & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5333 =>
                \$18844\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18844\ & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5336 =>
                \$18846\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18846\ & 
                work.Int.add(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5342 =>
                \$18848\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18848\ & 
                work.Int.add(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5348 =>
                \$18850\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18850\ & 
                work.Int.add(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5354 =>
                \$18852\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18852\ & 
                work.Int.add(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5360 =>
                \$18855_next_env\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18788\(16 to 47) & \$18854_sp\ & \$18855_next_env\ & 
                work.Int.add(\$18788\(96 to 103), work.Int.sub(eclat_resize(eclat_resize(
                                                               work.Int.lsr(
                                                               eclat_resize(eclat_resize(\$18853_hd\(0 to 30),16),31), X"0000000" & X"2"),16),8), "00000010")) & \$18788\(104 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5366 =>
                \$18859\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5365\ := \$ram_lock\;
                if \$v5365\(0) = '1' then
                  state_var5920 := Q_WAIT5364;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18856_loop_push6494360_arg\(0 to 15)));
                  \$ram_write\ <= \$18859\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5363;
                end if;
              when PAUSE_GET5370 =>
                \$18853_hd\ := \$ram_value\;
                release(\$ram_lock\);
                \$18856_loop_push6494360_id\ := "000000111000";
                \$18856_loop_push6494360_arg\ := \$18788\(48 to 63) & "00000000" & \$18788\(64 to 95) & eclat_resize(eclat_resize(
                work.Int.lsr(eclat_resize(eclat_resize(\$18853_hd\(0 to 30),16),31), X"0000000" & X"2"),16),8);
                state_var5920 := \$18856_LOOP_PUSH6494360\;
              when PAUSE_GET5385 =>
                \$18866_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18866_v\ & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5388 =>
                \$18868_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18868_v\ & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5391 =>
                \$18870_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18870_v\ & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5394 =>
                \$18872_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18872_v\ & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5400 =>
                \$18873_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5399\ := \$ram_lock\;
                if \$v5399\(0) = '1' then
                  state_var5920 := Q_WAIT5398;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$18788\(16 to 46),16), X"000" & X"0"), X"000" & X"1")));
                  \$ram_write\ <= \$18873_v\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5397;
                end if;
              when PAUSE_GET5406 =>
                \$18875_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5405\ := \$ram_lock\;
                if \$v5405\(0) = '1' then
                  state_var5920 := Q_WAIT5404;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$18788\(16 to 46),16), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= \$18875_v\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5403;
                end if;
              when PAUSE_GET5412 =>
                \$18877_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5411\ := \$ram_lock\;
                if \$v5411\(0) = '1' then
                  state_var5920 := Q_WAIT5410;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$18788\(16 to 46),16), X"000" & X"2"), X"000" & X"1")));
                  \$ram_write\ <= \$18877_v\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5409;
                end if;
              when PAUSE_GET5418 =>
                \$18879_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5417\ := \$ram_lock\;
                if \$v5417\(0) = '1' then
                  state_var5920 := Q_WAIT5416;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$18788\(16 to 46),16), X"000" & X"3"), X"000" & X"1")));
                  \$ram_write\ <= \$18879_v\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5415;
                end if;
              when PAUSE_GET5421 =>
                \$18881_hd\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & eclat_resize(eclat_resize(
                work.Int.lsr(eclat_resize(eclat_resize(\$18881_hd\(0 to 30),16),31), X"0000000" & X"2"),16),31) & eclat_true & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5424 =>
                \$18883_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18883_v\ & 
                work.Int.sub(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5427 =>
                \$18882_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5426\ := \$ram_lock\;
                if \$v5426\(0) = '1' then
                  state_var5920 := Q_WAIT5425;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18788\(16 to 46),16), eclat_resize(\$18882_v\(0 to 30),16)), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5424;
                end if;
              when PAUSE_GET5433 =>
                \$18885_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5432\ := \$ram_lock\;
                if \$v5432\(0) = '1' then
                  state_var5920 := Q_WAIT5431;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$18788\(16 to 46),16), eclat_resize(\$18884_v\(0 to 30),16)), X"000" & X"1")));
                  \$ram_write\ <= \$18885_v\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5430;
                end if;
              when PAUSE_GET5436 =>
                \$18884_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5435\ := \$ram_lock\;
                if \$v5435\(0) = '1' then
                  state_var5920 := Q_WAIT5434;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5433;
                end if;
              when PAUSE_GET5439 =>
                \$18888_next_acc\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18888_next_acc\ & 
                work.Int.sub(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5442 =>
                \$18887_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5441\ := \$ram_lock\;
                if \$v5441\(0) = '1' then
                  state_var5920 := Q_WAIT5440;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18788\(16 to 46),16), eclat_resize(\$18887_v\(0 to 30),16)), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5439;
                end if;
              when PAUSE_GET5448 =>
                \$18890_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5447\ := \$ram_lock\;
                if \$v5447\(0) = '1' then
                  state_var5920 := Q_WAIT5446;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$18788\(16 to 46),16), eclat_resize(\$18889_v\(0 to 30),16)), X"000" & X"1")));
                  \$ram_write\ <= \$18890_v\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5445;
                end if;
              when PAUSE_GET5451 =>
                \$18889_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5450\ := \$ram_lock\;
                if \$v5450\(0) = '1' then
                  state_var5920 := Q_WAIT5449;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5448;
                end if;
              when PAUSE_GET5454 =>
                \$18892_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18788\(16 to 47) & 
                work.Int.sub(work.Int.sub(work.Int.sub(\$18788\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"2") & \$18788\(64 to 95) & \$18788\(96 to 103) & eclat_resize(\$18892_v\(0 to 30),16) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5457 =>
                \$18896_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := eclat_resize(\$18893_v\(0 to 30),16) & \$18788\(16 to 47) & 
                work.Int.sub(work.Int.sub(work.Int.sub(work.Int.sub(\$18788\(104 to 119), X"000" & X"1"), X"000" & X"1"), X"000" & X"1"), X"000" & X"1") & \$18895_v\ & eclat_resize(\$18896_v\(0 to 30),8) & eclat_resize(\$18894_v\(0 to 30),16) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5460 =>
                \$18895_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5459\ := \$ram_lock\;
                if \$v5459\(0) = '1' then
                  state_var5920 := Q_WAIT5458;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$18788\(104 to 119), X"000" & X"1"), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5457;
                end if;
              when PAUSE_GET5463 =>
                \$18894_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5462\ := \$ram_lock\;
                if \$v5462\(0) = '1' then
                  state_var5920 := Q_WAIT5461;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$18788\(104 to 119), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5460;
                end if;
              when PAUSE_GET5466 =>
                \$18893_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5465\ := \$ram_lock\;
                if \$v5465\(0) = '1' then
                  state_var5920 := Q_WAIT5464;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$18788\(104 to 119), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5463;
                end if;
              when PAUSE_GET5488 =>
                \$18904_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5487\ := \$18901_binop_int6434361_arg\(0 to 31);
                case \$v5487\ is
                when X"0000000" & X"0" =>
                  \$18905_res\ := work.Int.add(\$18901_binop_int6434361_arg\(48 to 78), \$18904_v\(0 to 30));
                  \$18901_binop_int6434361_result\ := work.Int.add(\$18901_binop_int6434361_arg\(32 to 47), X"000" & X"1") & \$18905_res\ & eclat_true & 
                  work.Int.sub(\$18901_binop_int6434361_arg\(80 to 95), X"000" & X"1") & \$18901_binop_int6434361_arg\(96 to 151) & \$18901_binop_int6434361_arg\(152 to 153);
                  result4928 := \$18901_binop_int6434361_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"1" =>
                  \$18905_res\ := work.Int.sub(\$18901_binop_int6434361_arg\(48 to 78), \$18904_v\(0 to 30));
                  \$18901_binop_int6434361_result\ := work.Int.add(\$18901_binop_int6434361_arg\(32 to 47), X"000" & X"1") & \$18905_res\ & eclat_true & 
                  work.Int.sub(\$18901_binop_int6434361_arg\(80 to 95), X"000" & X"1") & \$18901_binop_int6434361_arg\(96 to 151) & \$18901_binop_int6434361_arg\(152 to 153);
                  result4928 := \$18901_binop_int6434361_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"2" =>
                  \$18905_res\ := work.Int.mul(\$18901_binop_int6434361_arg\(48 to 78), \$18904_v\(0 to 30));
                  \$18901_binop_int6434361_result\ := work.Int.add(\$18901_binop_int6434361_arg\(32 to 47), X"000" & X"1") & \$18905_res\ & eclat_true & 
                  work.Int.sub(\$18901_binop_int6434361_arg\(80 to 95), X"000" & X"1") & \$18901_binop_int6434361_arg\(96 to 151) & \$18901_binop_int6434361_arg\(152 to 153);
                  result4928 := \$18901_binop_int6434361_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"3" =>
                  \$v5483\ := work.Int.eq(\$18904_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v5483\(0) = '1' then
                    \$18905_res\ := "000"& X"000000" & X"0";
                    \$18901_binop_int6434361_result\ := work.Int.add(
                                                        \$18901_binop_int6434361_arg\(32 to 47), X"000" & X"1") & \$18905_res\ & eclat_true & 
                    work.Int.sub(\$18901_binop_int6434361_arg\(80 to 95), X"000" & X"1") & \$18901_binop_int6434361_arg\(96 to 151) & \$18901_binop_int6434361_arg\(152 to 153);
                    result4928 := \$18901_binop_int6434361_result\;
                    rdy4929 := eclat_true;
                    state_var5920 := IDLE4930;
                  else
                    \$18907_modulo6684356_id\ := "000001000100";
                    \$18907_modulo6684356_arg\ := work.Int.absv(\$18901_binop_int6434361_arg\(48 to 78)) & 
                    work.Int.absv(\$18904_v\(0 to 30));
                    state_var5920 := \$18907_MODULO6684356\;
                  end if;
                when X"0000000" & X"4" =>
                  \$v5486\ := work.Int.eq(\$18904_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v5486\(0) = '1' then
                    \$18905_res\ := "000"& X"000000" & X"0";
                    \$18901_binop_int6434361_result\ := work.Int.add(
                                                        \$18901_binop_int6434361_arg\(32 to 47), X"000" & X"1") & \$18905_res\ & eclat_true & 
                    work.Int.sub(\$18901_binop_int6434361_arg\(80 to 95), X"000" & X"1") & \$18901_binop_int6434361_arg\(96 to 151) & \$18901_binop_int6434361_arg\(152 to 153);
                    result4928 := \$18901_binop_int6434361_result\;
                    rdy4929 := eclat_true;
                    state_var5920 := IDLE4930;
                  else
                    \$18914_modulo6684357_id\ := "000001000110";
                    \$18914_modulo6684357_arg\ := work.Int.absv(\$18901_binop_int6434361_arg\(48 to 78)) & 
                    work.Int.absv(\$18904_v\(0 to 30));
                    state_var5920 := \$18914_MODULO6684357\;
                  end if;
                when X"0000000" & X"5" =>
                  \$18905_res\ := work.Int.land(\$18901_binop_int6434361_arg\(48 to 78), \$18904_v\(0 to 30));
                  \$18901_binop_int6434361_result\ := work.Int.add(\$18901_binop_int6434361_arg\(32 to 47), X"000" & X"1") & \$18905_res\ & eclat_true & 
                  work.Int.sub(\$18901_binop_int6434361_arg\(80 to 95), X"000" & X"1") & \$18901_binop_int6434361_arg\(96 to 151) & \$18901_binop_int6434361_arg\(152 to 153);
                  result4928 := \$18901_binop_int6434361_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"6" =>
                  \$18905_res\ := work.Int.lor(\$18901_binop_int6434361_arg\(48 to 78), \$18904_v\(0 to 30));
                  \$18901_binop_int6434361_result\ := work.Int.add(\$18901_binop_int6434361_arg\(32 to 47), X"000" & X"1") & \$18905_res\ & eclat_true & 
                  work.Int.sub(\$18901_binop_int6434361_arg\(80 to 95), X"000" & X"1") & \$18901_binop_int6434361_arg\(96 to 151) & \$18901_binop_int6434361_arg\(152 to 153);
                  result4928 := \$18901_binop_int6434361_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"7" =>
                  \$18905_res\ := work.Int.lxor(\$18901_binop_int6434361_arg\(48 to 78), \$18904_v\(0 to 30));
                  \$18901_binop_int6434361_result\ := work.Int.add(\$18901_binop_int6434361_arg\(32 to 47), X"000" & X"1") & \$18905_res\ & eclat_true & 
                  work.Int.sub(\$18901_binop_int6434361_arg\(80 to 95), X"000" & X"1") & \$18901_binop_int6434361_arg\(96 to 151) & \$18901_binop_int6434361_arg\(152 to 153);
                  result4928 := \$18901_binop_int6434361_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"8" =>
                  \$18905_res\ := work.Int.lsl(\$18901_binop_int6434361_arg\(48 to 78), \$18904_v\(0 to 30));
                  \$18901_binop_int6434361_result\ := work.Int.add(\$18901_binop_int6434361_arg\(32 to 47), X"000" & X"1") & \$18905_res\ & eclat_true & 
                  work.Int.sub(\$18901_binop_int6434361_arg\(80 to 95), X"000" & X"1") & \$18901_binop_int6434361_arg\(96 to 151) & \$18901_binop_int6434361_arg\(152 to 153);
                  result4928 := \$18901_binop_int6434361_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"9" =>
                  \$18905_res\ := work.Int.lsr(\$18901_binop_int6434361_arg\(48 to 78), \$18904_v\(0 to 30));
                  \$18901_binop_int6434361_result\ := work.Int.add(\$18901_binop_int6434361_arg\(32 to 47), X"000" & X"1") & \$18905_res\ & eclat_true & 
                  work.Int.sub(\$18901_binop_int6434361_arg\(80 to 95), X"000" & X"1") & \$18901_binop_int6434361_arg\(96 to 151) & \$18901_binop_int6434361_arg\(152 to 153);
                  result4928 := \$18901_binop_int6434361_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"a" =>
                  \$18905_res\ := work.Int.asr(\$18901_binop_int6434361_arg\(48 to 78), \$18904_v\(0 to 30));
                  \$18901_binop_int6434361_result\ := work.Int.add(\$18901_binop_int6434361_arg\(32 to 47), X"000" & X"1") & \$18905_res\ & eclat_true & 
                  work.Int.sub(\$18901_binop_int6434361_arg\(80 to 95), X"000" & X"1") & \$18901_binop_int6434361_arg\(96 to 151) & \$18901_binop_int6434361_arg\(152 to 153);
                  result4928 := \$18901_binop_int6434361_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"b" =>
                  \$18905_res\ := eclat_if(work.Int.lt(\$18901_binop_int6434361_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$18904_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.gt(\$18901_binop_int6434361_arg\(48 to 78), \$18904_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$18904_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"0" & 
                                  eclat_if(work.Int.lt(\$18901_binop_int6434361_arg\(48 to 78), \$18904_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$18901_binop_int6434361_result\ := work.Int.add(\$18901_binop_int6434361_arg\(32 to 47), X"000" & X"1") & \$18905_res\ & eclat_true & 
                  work.Int.sub(\$18901_binop_int6434361_arg\(80 to 95), X"000" & X"1") & \$18901_binop_int6434361_arg\(96 to 151) & \$18901_binop_int6434361_arg\(152 to 153);
                  result4928 := \$18901_binop_int6434361_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"c" =>
                  \$18905_res\ := eclat_if(work.Int.lt(\$18901_binop_int6434361_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$18904_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.le(\$18901_binop_int6434361_arg\(48 to 78), \$18904_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"1") & 
                                  eclat_if(work.Int.lt(\$18904_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & 
                                  eclat_if(work.Int.ge(\$18901_binop_int6434361_arg\(48 to 78), \$18904_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$18901_binop_int6434361_result\ := work.Int.add(\$18901_binop_int6434361_arg\(32 to 47), X"000" & X"1") & \$18905_res\ & eclat_true & 
                  work.Int.sub(\$18901_binop_int6434361_arg\(80 to 95), X"000" & X"1") & \$18901_binop_int6434361_arg\(96 to 151) & \$18901_binop_int6434361_arg\(152 to 153);
                  result4928 := \$18901_binop_int6434361_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when others =>
                  \$18905_res\ := "000"& X"000000" & X"0";
                  \$18901_binop_int6434361_result\ := work.Int.add(\$18901_binop_int6434361_arg\(32 to 47), X"000" & X"1") & \$18905_res\ & eclat_true & 
                  work.Int.sub(\$18901_binop_int6434361_arg\(80 to 95), X"000" & X"1") & \$18901_binop_int6434361_arg\(96 to 151) & \$18901_binop_int6434361_arg\(152 to 153);
                  result4928 := \$18901_binop_int6434361_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                end case;
              when PAUSE_GET5498 =>
                \$18923_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5497\ := \$18920_binop_int6434362_arg\(0 to 31);
                case \$v5497\ is
                when X"0000000" & X"0" =>
                  \$18924_res\ := work.Int.add(\$18920_binop_int6434362_arg\(48 to 78), \$18923_v\(0 to 30));
                  \$18920_binop_int6434362_result\ := work.Int.add(\$18920_binop_int6434362_arg\(32 to 47), X"000" & X"1") & \$18924_res\ & eclat_true & 
                  work.Int.sub(\$18920_binop_int6434362_arg\(80 to 95), X"000" & X"1") & \$18920_binop_int6434362_arg\(96 to 151) & \$18920_binop_int6434362_arg\(152 to 153);
                  result4928 := \$18920_binop_int6434362_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"1" =>
                  \$18924_res\ := work.Int.sub(\$18920_binop_int6434362_arg\(48 to 78), \$18923_v\(0 to 30));
                  \$18920_binop_int6434362_result\ := work.Int.add(\$18920_binop_int6434362_arg\(32 to 47), X"000" & X"1") & \$18924_res\ & eclat_true & 
                  work.Int.sub(\$18920_binop_int6434362_arg\(80 to 95), X"000" & X"1") & \$18920_binop_int6434362_arg\(96 to 151) & \$18920_binop_int6434362_arg\(152 to 153);
                  result4928 := \$18920_binop_int6434362_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"2" =>
                  \$18924_res\ := work.Int.mul(\$18920_binop_int6434362_arg\(48 to 78), \$18923_v\(0 to 30));
                  \$18920_binop_int6434362_result\ := work.Int.add(\$18920_binop_int6434362_arg\(32 to 47), X"000" & X"1") & \$18924_res\ & eclat_true & 
                  work.Int.sub(\$18920_binop_int6434362_arg\(80 to 95), X"000" & X"1") & \$18920_binop_int6434362_arg\(96 to 151) & \$18920_binop_int6434362_arg\(152 to 153);
                  result4928 := \$18920_binop_int6434362_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"3" =>
                  \$v5493\ := work.Int.eq(\$18923_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v5493\(0) = '1' then
                    \$18924_res\ := "000"& X"000000" & X"0";
                    \$18920_binop_int6434362_result\ := work.Int.add(
                                                        \$18920_binop_int6434362_arg\(32 to 47), X"000" & X"1") & \$18924_res\ & eclat_true & 
                    work.Int.sub(\$18920_binop_int6434362_arg\(80 to 95), X"000" & X"1") & \$18920_binop_int6434362_arg\(96 to 151) & \$18920_binop_int6434362_arg\(152 to 153);
                    result4928 := \$18920_binop_int6434362_result\;
                    rdy4929 := eclat_true;
                    state_var5920 := IDLE4930;
                  else
                    \$18926_modulo6684356_id\ := "000001001001";
                    \$18926_modulo6684356_arg\ := work.Int.absv(\$18920_binop_int6434362_arg\(48 to 78)) & 
                    work.Int.absv(\$18923_v\(0 to 30));
                    state_var5920 := \$18926_MODULO6684356\;
                  end if;
                when X"0000000" & X"4" =>
                  \$v5496\ := work.Int.eq(\$18923_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v5496\(0) = '1' then
                    \$18924_res\ := "000"& X"000000" & X"0";
                    \$18920_binop_int6434362_result\ := work.Int.add(
                                                        \$18920_binop_int6434362_arg\(32 to 47), X"000" & X"1") & \$18924_res\ & eclat_true & 
                    work.Int.sub(\$18920_binop_int6434362_arg\(80 to 95), X"000" & X"1") & \$18920_binop_int6434362_arg\(96 to 151) & \$18920_binop_int6434362_arg\(152 to 153);
                    result4928 := \$18920_binop_int6434362_result\;
                    rdy4929 := eclat_true;
                    state_var5920 := IDLE4930;
                  else
                    \$18933_modulo6684357_id\ := "000001001011";
                    \$18933_modulo6684357_arg\ := work.Int.absv(\$18920_binop_int6434362_arg\(48 to 78)) & 
                    work.Int.absv(\$18923_v\(0 to 30));
                    state_var5920 := \$18933_MODULO6684357\;
                  end if;
                when X"0000000" & X"5" =>
                  \$18924_res\ := work.Int.land(\$18920_binop_int6434362_arg\(48 to 78), \$18923_v\(0 to 30));
                  \$18920_binop_int6434362_result\ := work.Int.add(\$18920_binop_int6434362_arg\(32 to 47), X"000" & X"1") & \$18924_res\ & eclat_true & 
                  work.Int.sub(\$18920_binop_int6434362_arg\(80 to 95), X"000" & X"1") & \$18920_binop_int6434362_arg\(96 to 151) & \$18920_binop_int6434362_arg\(152 to 153);
                  result4928 := \$18920_binop_int6434362_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"6" =>
                  \$18924_res\ := work.Int.lor(\$18920_binop_int6434362_arg\(48 to 78), \$18923_v\(0 to 30));
                  \$18920_binop_int6434362_result\ := work.Int.add(\$18920_binop_int6434362_arg\(32 to 47), X"000" & X"1") & \$18924_res\ & eclat_true & 
                  work.Int.sub(\$18920_binop_int6434362_arg\(80 to 95), X"000" & X"1") & \$18920_binop_int6434362_arg\(96 to 151) & \$18920_binop_int6434362_arg\(152 to 153);
                  result4928 := \$18920_binop_int6434362_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"7" =>
                  \$18924_res\ := work.Int.lxor(\$18920_binop_int6434362_arg\(48 to 78), \$18923_v\(0 to 30));
                  \$18920_binop_int6434362_result\ := work.Int.add(\$18920_binop_int6434362_arg\(32 to 47), X"000" & X"1") & \$18924_res\ & eclat_true & 
                  work.Int.sub(\$18920_binop_int6434362_arg\(80 to 95), X"000" & X"1") & \$18920_binop_int6434362_arg\(96 to 151) & \$18920_binop_int6434362_arg\(152 to 153);
                  result4928 := \$18920_binop_int6434362_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"8" =>
                  \$18924_res\ := work.Int.lsl(\$18920_binop_int6434362_arg\(48 to 78), \$18923_v\(0 to 30));
                  \$18920_binop_int6434362_result\ := work.Int.add(\$18920_binop_int6434362_arg\(32 to 47), X"000" & X"1") & \$18924_res\ & eclat_true & 
                  work.Int.sub(\$18920_binop_int6434362_arg\(80 to 95), X"000" & X"1") & \$18920_binop_int6434362_arg\(96 to 151) & \$18920_binop_int6434362_arg\(152 to 153);
                  result4928 := \$18920_binop_int6434362_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"9" =>
                  \$18924_res\ := work.Int.lsr(\$18920_binop_int6434362_arg\(48 to 78), \$18923_v\(0 to 30));
                  \$18920_binop_int6434362_result\ := work.Int.add(\$18920_binop_int6434362_arg\(32 to 47), X"000" & X"1") & \$18924_res\ & eclat_true & 
                  work.Int.sub(\$18920_binop_int6434362_arg\(80 to 95), X"000" & X"1") & \$18920_binop_int6434362_arg\(96 to 151) & \$18920_binop_int6434362_arg\(152 to 153);
                  result4928 := \$18920_binop_int6434362_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"a" =>
                  \$18924_res\ := work.Int.asr(\$18920_binop_int6434362_arg\(48 to 78), \$18923_v\(0 to 30));
                  \$18920_binop_int6434362_result\ := work.Int.add(\$18920_binop_int6434362_arg\(32 to 47), X"000" & X"1") & \$18924_res\ & eclat_true & 
                  work.Int.sub(\$18920_binop_int6434362_arg\(80 to 95), X"000" & X"1") & \$18920_binop_int6434362_arg\(96 to 151) & \$18920_binop_int6434362_arg\(152 to 153);
                  result4928 := \$18920_binop_int6434362_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"b" =>
                  \$18924_res\ := eclat_if(work.Int.lt(\$18920_binop_int6434362_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$18923_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.gt(\$18920_binop_int6434362_arg\(48 to 78), \$18923_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$18923_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"0" & 
                                  eclat_if(work.Int.lt(\$18920_binop_int6434362_arg\(48 to 78), \$18923_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$18920_binop_int6434362_result\ := work.Int.add(\$18920_binop_int6434362_arg\(32 to 47), X"000" & X"1") & \$18924_res\ & eclat_true & 
                  work.Int.sub(\$18920_binop_int6434362_arg\(80 to 95), X"000" & X"1") & \$18920_binop_int6434362_arg\(96 to 151) & \$18920_binop_int6434362_arg\(152 to 153);
                  result4928 := \$18920_binop_int6434362_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"c" =>
                  \$18924_res\ := eclat_if(work.Int.lt(\$18920_binop_int6434362_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$18923_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.le(\$18920_binop_int6434362_arg\(48 to 78), \$18923_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"1") & 
                                  eclat_if(work.Int.lt(\$18923_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & 
                                  eclat_if(work.Int.ge(\$18920_binop_int6434362_arg\(48 to 78), \$18923_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$18920_binop_int6434362_result\ := work.Int.add(\$18920_binop_int6434362_arg\(32 to 47), X"000" & X"1") & \$18924_res\ & eclat_true & 
                  work.Int.sub(\$18920_binop_int6434362_arg\(80 to 95), X"000" & X"1") & \$18920_binop_int6434362_arg\(96 to 151) & \$18920_binop_int6434362_arg\(152 to 153);
                  result4928 := \$18920_binop_int6434362_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when others =>
                  \$18924_res\ := "000"& X"000000" & X"0";
                  \$18920_binop_int6434362_result\ := work.Int.add(\$18920_binop_int6434362_arg\(32 to 47), X"000" & X"1") & \$18924_res\ & eclat_true & 
                  work.Int.sub(\$18920_binop_int6434362_arg\(80 to 95), X"000" & X"1") & \$18920_binop_int6434362_arg\(96 to 151) & \$18920_binop_int6434362_arg\(152 to 153);
                  result4928 := \$18920_binop_int6434362_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                end case;
              when PAUSE_GET5508 =>
                \$18942_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5507\ := \$18939_binop_int6434363_arg\(0 to 31);
                case \$v5507\ is
                when X"0000000" & X"0" =>
                  \$18943_res\ := work.Int.add(\$18939_binop_int6434363_arg\(48 to 78), \$18942_v\(0 to 30));
                  \$18939_binop_int6434363_result\ := work.Int.add(\$18939_binop_int6434363_arg\(32 to 47), X"000" & X"1") & \$18943_res\ & eclat_true & 
                  work.Int.sub(\$18939_binop_int6434363_arg\(80 to 95), X"000" & X"1") & \$18939_binop_int6434363_arg\(96 to 151) & \$18939_binop_int6434363_arg\(152 to 153);
                  result4928 := \$18939_binop_int6434363_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"1" =>
                  \$18943_res\ := work.Int.sub(\$18939_binop_int6434363_arg\(48 to 78), \$18942_v\(0 to 30));
                  \$18939_binop_int6434363_result\ := work.Int.add(\$18939_binop_int6434363_arg\(32 to 47), X"000" & X"1") & \$18943_res\ & eclat_true & 
                  work.Int.sub(\$18939_binop_int6434363_arg\(80 to 95), X"000" & X"1") & \$18939_binop_int6434363_arg\(96 to 151) & \$18939_binop_int6434363_arg\(152 to 153);
                  result4928 := \$18939_binop_int6434363_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"2" =>
                  \$18943_res\ := work.Int.mul(\$18939_binop_int6434363_arg\(48 to 78), \$18942_v\(0 to 30));
                  \$18939_binop_int6434363_result\ := work.Int.add(\$18939_binop_int6434363_arg\(32 to 47), X"000" & X"1") & \$18943_res\ & eclat_true & 
                  work.Int.sub(\$18939_binop_int6434363_arg\(80 to 95), X"000" & X"1") & \$18939_binop_int6434363_arg\(96 to 151) & \$18939_binop_int6434363_arg\(152 to 153);
                  result4928 := \$18939_binop_int6434363_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"3" =>
                  \$v5503\ := work.Int.eq(\$18942_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v5503\(0) = '1' then
                    \$18943_res\ := "000"& X"000000" & X"0";
                    \$18939_binop_int6434363_result\ := work.Int.add(
                                                        \$18939_binop_int6434363_arg\(32 to 47), X"000" & X"1") & \$18943_res\ & eclat_true & 
                    work.Int.sub(\$18939_binop_int6434363_arg\(80 to 95), X"000" & X"1") & \$18939_binop_int6434363_arg\(96 to 151) & \$18939_binop_int6434363_arg\(152 to 153);
                    result4928 := \$18939_binop_int6434363_result\;
                    rdy4929 := eclat_true;
                    state_var5920 := IDLE4930;
                  else
                    \$18945_modulo6684356_id\ := "000001001110";
                    \$18945_modulo6684356_arg\ := work.Int.absv(\$18939_binop_int6434363_arg\(48 to 78)) & 
                    work.Int.absv(\$18942_v\(0 to 30));
                    state_var5920 := \$18945_MODULO6684356\;
                  end if;
                when X"0000000" & X"4" =>
                  \$v5506\ := work.Int.eq(\$18942_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v5506\(0) = '1' then
                    \$18943_res\ := "000"& X"000000" & X"0";
                    \$18939_binop_int6434363_result\ := work.Int.add(
                                                        \$18939_binop_int6434363_arg\(32 to 47), X"000" & X"1") & \$18943_res\ & eclat_true & 
                    work.Int.sub(\$18939_binop_int6434363_arg\(80 to 95), X"000" & X"1") & \$18939_binop_int6434363_arg\(96 to 151) & \$18939_binop_int6434363_arg\(152 to 153);
                    result4928 := \$18939_binop_int6434363_result\;
                    rdy4929 := eclat_true;
                    state_var5920 := IDLE4930;
                  else
                    \$18952_modulo6684357_id\ := "000001010000";
                    \$18952_modulo6684357_arg\ := work.Int.absv(\$18939_binop_int6434363_arg\(48 to 78)) & 
                    work.Int.absv(\$18942_v\(0 to 30));
                    state_var5920 := \$18952_MODULO6684357\;
                  end if;
                when X"0000000" & X"5" =>
                  \$18943_res\ := work.Int.land(\$18939_binop_int6434363_arg\(48 to 78), \$18942_v\(0 to 30));
                  \$18939_binop_int6434363_result\ := work.Int.add(\$18939_binop_int6434363_arg\(32 to 47), X"000" & X"1") & \$18943_res\ & eclat_true & 
                  work.Int.sub(\$18939_binop_int6434363_arg\(80 to 95), X"000" & X"1") & \$18939_binop_int6434363_arg\(96 to 151) & \$18939_binop_int6434363_arg\(152 to 153);
                  result4928 := \$18939_binop_int6434363_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"6" =>
                  \$18943_res\ := work.Int.lor(\$18939_binop_int6434363_arg\(48 to 78), \$18942_v\(0 to 30));
                  \$18939_binop_int6434363_result\ := work.Int.add(\$18939_binop_int6434363_arg\(32 to 47), X"000" & X"1") & \$18943_res\ & eclat_true & 
                  work.Int.sub(\$18939_binop_int6434363_arg\(80 to 95), X"000" & X"1") & \$18939_binop_int6434363_arg\(96 to 151) & \$18939_binop_int6434363_arg\(152 to 153);
                  result4928 := \$18939_binop_int6434363_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"7" =>
                  \$18943_res\ := work.Int.lxor(\$18939_binop_int6434363_arg\(48 to 78), \$18942_v\(0 to 30));
                  \$18939_binop_int6434363_result\ := work.Int.add(\$18939_binop_int6434363_arg\(32 to 47), X"000" & X"1") & \$18943_res\ & eclat_true & 
                  work.Int.sub(\$18939_binop_int6434363_arg\(80 to 95), X"000" & X"1") & \$18939_binop_int6434363_arg\(96 to 151) & \$18939_binop_int6434363_arg\(152 to 153);
                  result4928 := \$18939_binop_int6434363_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"8" =>
                  \$18943_res\ := work.Int.lsl(\$18939_binop_int6434363_arg\(48 to 78), \$18942_v\(0 to 30));
                  \$18939_binop_int6434363_result\ := work.Int.add(\$18939_binop_int6434363_arg\(32 to 47), X"000" & X"1") & \$18943_res\ & eclat_true & 
                  work.Int.sub(\$18939_binop_int6434363_arg\(80 to 95), X"000" & X"1") & \$18939_binop_int6434363_arg\(96 to 151) & \$18939_binop_int6434363_arg\(152 to 153);
                  result4928 := \$18939_binop_int6434363_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"9" =>
                  \$18943_res\ := work.Int.lsr(\$18939_binop_int6434363_arg\(48 to 78), \$18942_v\(0 to 30));
                  \$18939_binop_int6434363_result\ := work.Int.add(\$18939_binop_int6434363_arg\(32 to 47), X"000" & X"1") & \$18943_res\ & eclat_true & 
                  work.Int.sub(\$18939_binop_int6434363_arg\(80 to 95), X"000" & X"1") & \$18939_binop_int6434363_arg\(96 to 151) & \$18939_binop_int6434363_arg\(152 to 153);
                  result4928 := \$18939_binop_int6434363_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"a" =>
                  \$18943_res\ := work.Int.asr(\$18939_binop_int6434363_arg\(48 to 78), \$18942_v\(0 to 30));
                  \$18939_binop_int6434363_result\ := work.Int.add(\$18939_binop_int6434363_arg\(32 to 47), X"000" & X"1") & \$18943_res\ & eclat_true & 
                  work.Int.sub(\$18939_binop_int6434363_arg\(80 to 95), X"000" & X"1") & \$18939_binop_int6434363_arg\(96 to 151) & \$18939_binop_int6434363_arg\(152 to 153);
                  result4928 := \$18939_binop_int6434363_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"b" =>
                  \$18943_res\ := eclat_if(work.Int.lt(\$18939_binop_int6434363_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$18942_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.gt(\$18939_binop_int6434363_arg\(48 to 78), \$18942_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$18942_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"0" & 
                                  eclat_if(work.Int.lt(\$18939_binop_int6434363_arg\(48 to 78), \$18942_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$18939_binop_int6434363_result\ := work.Int.add(\$18939_binop_int6434363_arg\(32 to 47), X"000" & X"1") & \$18943_res\ & eclat_true & 
                  work.Int.sub(\$18939_binop_int6434363_arg\(80 to 95), X"000" & X"1") & \$18939_binop_int6434363_arg\(96 to 151) & \$18939_binop_int6434363_arg\(152 to 153);
                  result4928 := \$18939_binop_int6434363_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"c" =>
                  \$18943_res\ := eclat_if(work.Int.lt(\$18939_binop_int6434363_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$18942_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.le(\$18939_binop_int6434363_arg\(48 to 78), \$18942_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"1") & 
                                  eclat_if(work.Int.lt(\$18942_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & 
                                  eclat_if(work.Int.ge(\$18939_binop_int6434363_arg\(48 to 78), \$18942_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$18939_binop_int6434363_result\ := work.Int.add(\$18939_binop_int6434363_arg\(32 to 47), X"000" & X"1") & \$18943_res\ & eclat_true & 
                  work.Int.sub(\$18939_binop_int6434363_arg\(80 to 95), X"000" & X"1") & \$18939_binop_int6434363_arg\(96 to 151) & \$18939_binop_int6434363_arg\(152 to 153);
                  result4928 := \$18939_binop_int6434363_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when others =>
                  \$18943_res\ := "000"& X"000000" & X"0";
                  \$18939_binop_int6434363_result\ := work.Int.add(\$18939_binop_int6434363_arg\(32 to 47), X"000" & X"1") & \$18943_res\ & eclat_true & 
                  work.Int.sub(\$18939_binop_int6434363_arg\(80 to 95), X"000" & X"1") & \$18939_binop_int6434363_arg\(96 to 151) & \$18939_binop_int6434363_arg\(152 to 153);
                  result4928 := \$18939_binop_int6434363_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                end case;
              when PAUSE_GET5518 =>
                \$18961_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5517\ := \$18958_binop_int6434364_arg\(0 to 31);
                case \$v5517\ is
                when X"0000000" & X"0" =>
                  \$18962_res\ := work.Int.add(\$18958_binop_int6434364_arg\(48 to 78), \$18961_v\(0 to 30));
                  \$18958_binop_int6434364_result\ := work.Int.add(\$18958_binop_int6434364_arg\(32 to 47), X"000" & X"1") & \$18962_res\ & eclat_true & 
                  work.Int.sub(\$18958_binop_int6434364_arg\(80 to 95), X"000" & X"1") & \$18958_binop_int6434364_arg\(96 to 151) & \$18958_binop_int6434364_arg\(152 to 153);
                  result4928 := \$18958_binop_int6434364_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"1" =>
                  \$18962_res\ := work.Int.sub(\$18958_binop_int6434364_arg\(48 to 78), \$18961_v\(0 to 30));
                  \$18958_binop_int6434364_result\ := work.Int.add(\$18958_binop_int6434364_arg\(32 to 47), X"000" & X"1") & \$18962_res\ & eclat_true & 
                  work.Int.sub(\$18958_binop_int6434364_arg\(80 to 95), X"000" & X"1") & \$18958_binop_int6434364_arg\(96 to 151) & \$18958_binop_int6434364_arg\(152 to 153);
                  result4928 := \$18958_binop_int6434364_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"2" =>
                  \$18962_res\ := work.Int.mul(\$18958_binop_int6434364_arg\(48 to 78), \$18961_v\(0 to 30));
                  \$18958_binop_int6434364_result\ := work.Int.add(\$18958_binop_int6434364_arg\(32 to 47), X"000" & X"1") & \$18962_res\ & eclat_true & 
                  work.Int.sub(\$18958_binop_int6434364_arg\(80 to 95), X"000" & X"1") & \$18958_binop_int6434364_arg\(96 to 151) & \$18958_binop_int6434364_arg\(152 to 153);
                  result4928 := \$18958_binop_int6434364_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"3" =>
                  \$v5513\ := work.Int.eq(\$18961_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v5513\(0) = '1' then
                    \$18962_res\ := "000"& X"000000" & X"0";
                    \$18958_binop_int6434364_result\ := work.Int.add(
                                                        \$18958_binop_int6434364_arg\(32 to 47), X"000" & X"1") & \$18962_res\ & eclat_true & 
                    work.Int.sub(\$18958_binop_int6434364_arg\(80 to 95), X"000" & X"1") & \$18958_binop_int6434364_arg\(96 to 151) & \$18958_binop_int6434364_arg\(152 to 153);
                    result4928 := \$18958_binop_int6434364_result\;
                    rdy4929 := eclat_true;
                    state_var5920 := IDLE4930;
                  else
                    \$18964_modulo6684356_id\ := "000001010011";
                    \$18964_modulo6684356_arg\ := work.Int.absv(\$18958_binop_int6434364_arg\(48 to 78)) & 
                    work.Int.absv(\$18961_v\(0 to 30));
                    state_var5920 := \$18964_MODULO6684356\;
                  end if;
                when X"0000000" & X"4" =>
                  \$v5516\ := work.Int.eq(\$18961_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v5516\(0) = '1' then
                    \$18962_res\ := "000"& X"000000" & X"0";
                    \$18958_binop_int6434364_result\ := work.Int.add(
                                                        \$18958_binop_int6434364_arg\(32 to 47), X"000" & X"1") & \$18962_res\ & eclat_true & 
                    work.Int.sub(\$18958_binop_int6434364_arg\(80 to 95), X"000" & X"1") & \$18958_binop_int6434364_arg\(96 to 151) & \$18958_binop_int6434364_arg\(152 to 153);
                    result4928 := \$18958_binop_int6434364_result\;
                    rdy4929 := eclat_true;
                    state_var5920 := IDLE4930;
                  else
                    \$18971_modulo6684357_id\ := "000001010101";
                    \$18971_modulo6684357_arg\ := work.Int.absv(\$18958_binop_int6434364_arg\(48 to 78)) & 
                    work.Int.absv(\$18961_v\(0 to 30));
                    state_var5920 := \$18971_MODULO6684357\;
                  end if;
                when X"0000000" & X"5" =>
                  \$18962_res\ := work.Int.land(\$18958_binop_int6434364_arg\(48 to 78), \$18961_v\(0 to 30));
                  \$18958_binop_int6434364_result\ := work.Int.add(\$18958_binop_int6434364_arg\(32 to 47), X"000" & X"1") & \$18962_res\ & eclat_true & 
                  work.Int.sub(\$18958_binop_int6434364_arg\(80 to 95), X"000" & X"1") & \$18958_binop_int6434364_arg\(96 to 151) & \$18958_binop_int6434364_arg\(152 to 153);
                  result4928 := \$18958_binop_int6434364_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"6" =>
                  \$18962_res\ := work.Int.lor(\$18958_binop_int6434364_arg\(48 to 78), \$18961_v\(0 to 30));
                  \$18958_binop_int6434364_result\ := work.Int.add(\$18958_binop_int6434364_arg\(32 to 47), X"000" & X"1") & \$18962_res\ & eclat_true & 
                  work.Int.sub(\$18958_binop_int6434364_arg\(80 to 95), X"000" & X"1") & \$18958_binop_int6434364_arg\(96 to 151) & \$18958_binop_int6434364_arg\(152 to 153);
                  result4928 := \$18958_binop_int6434364_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"7" =>
                  \$18962_res\ := work.Int.lxor(\$18958_binop_int6434364_arg\(48 to 78), \$18961_v\(0 to 30));
                  \$18958_binop_int6434364_result\ := work.Int.add(\$18958_binop_int6434364_arg\(32 to 47), X"000" & X"1") & \$18962_res\ & eclat_true & 
                  work.Int.sub(\$18958_binop_int6434364_arg\(80 to 95), X"000" & X"1") & \$18958_binop_int6434364_arg\(96 to 151) & \$18958_binop_int6434364_arg\(152 to 153);
                  result4928 := \$18958_binop_int6434364_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"8" =>
                  \$18962_res\ := work.Int.lsl(\$18958_binop_int6434364_arg\(48 to 78), \$18961_v\(0 to 30));
                  \$18958_binop_int6434364_result\ := work.Int.add(\$18958_binop_int6434364_arg\(32 to 47), X"000" & X"1") & \$18962_res\ & eclat_true & 
                  work.Int.sub(\$18958_binop_int6434364_arg\(80 to 95), X"000" & X"1") & \$18958_binop_int6434364_arg\(96 to 151) & \$18958_binop_int6434364_arg\(152 to 153);
                  result4928 := \$18958_binop_int6434364_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"9" =>
                  \$18962_res\ := work.Int.lsr(\$18958_binop_int6434364_arg\(48 to 78), \$18961_v\(0 to 30));
                  \$18958_binop_int6434364_result\ := work.Int.add(\$18958_binop_int6434364_arg\(32 to 47), X"000" & X"1") & \$18962_res\ & eclat_true & 
                  work.Int.sub(\$18958_binop_int6434364_arg\(80 to 95), X"000" & X"1") & \$18958_binop_int6434364_arg\(96 to 151) & \$18958_binop_int6434364_arg\(152 to 153);
                  result4928 := \$18958_binop_int6434364_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"a" =>
                  \$18962_res\ := work.Int.asr(\$18958_binop_int6434364_arg\(48 to 78), \$18961_v\(0 to 30));
                  \$18958_binop_int6434364_result\ := work.Int.add(\$18958_binop_int6434364_arg\(32 to 47), X"000" & X"1") & \$18962_res\ & eclat_true & 
                  work.Int.sub(\$18958_binop_int6434364_arg\(80 to 95), X"000" & X"1") & \$18958_binop_int6434364_arg\(96 to 151) & \$18958_binop_int6434364_arg\(152 to 153);
                  result4928 := \$18958_binop_int6434364_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"b" =>
                  \$18962_res\ := eclat_if(work.Int.lt(\$18958_binop_int6434364_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$18961_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.gt(\$18958_binop_int6434364_arg\(48 to 78), \$18961_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$18961_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"0" & 
                                  eclat_if(work.Int.lt(\$18958_binop_int6434364_arg\(48 to 78), \$18961_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$18958_binop_int6434364_result\ := work.Int.add(\$18958_binop_int6434364_arg\(32 to 47), X"000" & X"1") & \$18962_res\ & eclat_true & 
                  work.Int.sub(\$18958_binop_int6434364_arg\(80 to 95), X"000" & X"1") & \$18958_binop_int6434364_arg\(96 to 151) & \$18958_binop_int6434364_arg\(152 to 153);
                  result4928 := \$18958_binop_int6434364_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"c" =>
                  \$18962_res\ := eclat_if(work.Int.lt(\$18958_binop_int6434364_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$18961_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.le(\$18958_binop_int6434364_arg\(48 to 78), \$18961_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"1") & 
                                  eclat_if(work.Int.lt(\$18961_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & 
                                  eclat_if(work.Int.ge(\$18958_binop_int6434364_arg\(48 to 78), \$18961_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$18958_binop_int6434364_result\ := work.Int.add(\$18958_binop_int6434364_arg\(32 to 47), X"000" & X"1") & \$18962_res\ & eclat_true & 
                  work.Int.sub(\$18958_binop_int6434364_arg\(80 to 95), X"000" & X"1") & \$18958_binop_int6434364_arg\(96 to 151) & \$18958_binop_int6434364_arg\(152 to 153);
                  result4928 := \$18958_binop_int6434364_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when others =>
                  \$18962_res\ := "000"& X"000000" & X"0";
                  \$18958_binop_int6434364_result\ := work.Int.add(\$18958_binop_int6434364_arg\(32 to 47), X"000" & X"1") & \$18962_res\ & eclat_true & 
                  work.Int.sub(\$18958_binop_int6434364_arg\(80 to 95), X"000" & X"1") & \$18958_binop_int6434364_arg\(96 to 151) & \$18958_binop_int6434364_arg\(152 to 153);
                  result4928 := \$18958_binop_int6434364_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                end case;
              when PAUSE_GET5528 =>
                \$18980_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5527\ := \$18977_binop_int6434365_arg\(0 to 31);
                case \$v5527\ is
                when X"0000000" & X"0" =>
                  \$18981_res\ := work.Int.add(\$18977_binop_int6434365_arg\(48 to 78), \$18980_v\(0 to 30));
                  \$18977_binop_int6434365_result\ := work.Int.add(\$18977_binop_int6434365_arg\(32 to 47), X"000" & X"1") & \$18981_res\ & eclat_true & 
                  work.Int.sub(\$18977_binop_int6434365_arg\(80 to 95), X"000" & X"1") & \$18977_binop_int6434365_arg\(96 to 151) & \$18977_binop_int6434365_arg\(152 to 153);
                  result4928 := \$18977_binop_int6434365_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"1" =>
                  \$18981_res\ := work.Int.sub(\$18977_binop_int6434365_arg\(48 to 78), \$18980_v\(0 to 30));
                  \$18977_binop_int6434365_result\ := work.Int.add(\$18977_binop_int6434365_arg\(32 to 47), X"000" & X"1") & \$18981_res\ & eclat_true & 
                  work.Int.sub(\$18977_binop_int6434365_arg\(80 to 95), X"000" & X"1") & \$18977_binop_int6434365_arg\(96 to 151) & \$18977_binop_int6434365_arg\(152 to 153);
                  result4928 := \$18977_binop_int6434365_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"2" =>
                  \$18981_res\ := work.Int.mul(\$18977_binop_int6434365_arg\(48 to 78), \$18980_v\(0 to 30));
                  \$18977_binop_int6434365_result\ := work.Int.add(\$18977_binop_int6434365_arg\(32 to 47), X"000" & X"1") & \$18981_res\ & eclat_true & 
                  work.Int.sub(\$18977_binop_int6434365_arg\(80 to 95), X"000" & X"1") & \$18977_binop_int6434365_arg\(96 to 151) & \$18977_binop_int6434365_arg\(152 to 153);
                  result4928 := \$18977_binop_int6434365_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"3" =>
                  \$v5523\ := work.Int.eq(\$18980_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v5523\(0) = '1' then
                    \$18981_res\ := "000"& X"000000" & X"0";
                    \$18977_binop_int6434365_result\ := work.Int.add(
                                                        \$18977_binop_int6434365_arg\(32 to 47), X"000" & X"1") & \$18981_res\ & eclat_true & 
                    work.Int.sub(\$18977_binop_int6434365_arg\(80 to 95), X"000" & X"1") & \$18977_binop_int6434365_arg\(96 to 151) & \$18977_binop_int6434365_arg\(152 to 153);
                    result4928 := \$18977_binop_int6434365_result\;
                    rdy4929 := eclat_true;
                    state_var5920 := IDLE4930;
                  else
                    \$18983_modulo6684356_id\ := "000001011000";
                    \$18983_modulo6684356_arg\ := work.Int.absv(\$18977_binop_int6434365_arg\(48 to 78)) & 
                    work.Int.absv(\$18980_v\(0 to 30));
                    state_var5920 := \$18983_MODULO6684356\;
                  end if;
                when X"0000000" & X"4" =>
                  \$v5526\ := work.Int.eq(\$18980_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v5526\(0) = '1' then
                    \$18981_res\ := "000"& X"000000" & X"0";
                    \$18977_binop_int6434365_result\ := work.Int.add(
                                                        \$18977_binop_int6434365_arg\(32 to 47), X"000" & X"1") & \$18981_res\ & eclat_true & 
                    work.Int.sub(\$18977_binop_int6434365_arg\(80 to 95), X"000" & X"1") & \$18977_binop_int6434365_arg\(96 to 151) & \$18977_binop_int6434365_arg\(152 to 153);
                    result4928 := \$18977_binop_int6434365_result\;
                    rdy4929 := eclat_true;
                    state_var5920 := IDLE4930;
                  else
                    \$18990_modulo6684357_id\ := "000001011010";
                    \$18990_modulo6684357_arg\ := work.Int.absv(\$18977_binop_int6434365_arg\(48 to 78)) & 
                    work.Int.absv(\$18980_v\(0 to 30));
                    state_var5920 := \$18990_MODULO6684357\;
                  end if;
                when X"0000000" & X"5" =>
                  \$18981_res\ := work.Int.land(\$18977_binop_int6434365_arg\(48 to 78), \$18980_v\(0 to 30));
                  \$18977_binop_int6434365_result\ := work.Int.add(\$18977_binop_int6434365_arg\(32 to 47), X"000" & X"1") & \$18981_res\ & eclat_true & 
                  work.Int.sub(\$18977_binop_int6434365_arg\(80 to 95), X"000" & X"1") & \$18977_binop_int6434365_arg\(96 to 151) & \$18977_binop_int6434365_arg\(152 to 153);
                  result4928 := \$18977_binop_int6434365_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"6" =>
                  \$18981_res\ := work.Int.lor(\$18977_binop_int6434365_arg\(48 to 78), \$18980_v\(0 to 30));
                  \$18977_binop_int6434365_result\ := work.Int.add(\$18977_binop_int6434365_arg\(32 to 47), X"000" & X"1") & \$18981_res\ & eclat_true & 
                  work.Int.sub(\$18977_binop_int6434365_arg\(80 to 95), X"000" & X"1") & \$18977_binop_int6434365_arg\(96 to 151) & \$18977_binop_int6434365_arg\(152 to 153);
                  result4928 := \$18977_binop_int6434365_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"7" =>
                  \$18981_res\ := work.Int.lxor(\$18977_binop_int6434365_arg\(48 to 78), \$18980_v\(0 to 30));
                  \$18977_binop_int6434365_result\ := work.Int.add(\$18977_binop_int6434365_arg\(32 to 47), X"000" & X"1") & \$18981_res\ & eclat_true & 
                  work.Int.sub(\$18977_binop_int6434365_arg\(80 to 95), X"000" & X"1") & \$18977_binop_int6434365_arg\(96 to 151) & \$18977_binop_int6434365_arg\(152 to 153);
                  result4928 := \$18977_binop_int6434365_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"8" =>
                  \$18981_res\ := work.Int.lsl(\$18977_binop_int6434365_arg\(48 to 78), \$18980_v\(0 to 30));
                  \$18977_binop_int6434365_result\ := work.Int.add(\$18977_binop_int6434365_arg\(32 to 47), X"000" & X"1") & \$18981_res\ & eclat_true & 
                  work.Int.sub(\$18977_binop_int6434365_arg\(80 to 95), X"000" & X"1") & \$18977_binop_int6434365_arg\(96 to 151) & \$18977_binop_int6434365_arg\(152 to 153);
                  result4928 := \$18977_binop_int6434365_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"9" =>
                  \$18981_res\ := work.Int.lsr(\$18977_binop_int6434365_arg\(48 to 78), \$18980_v\(0 to 30));
                  \$18977_binop_int6434365_result\ := work.Int.add(\$18977_binop_int6434365_arg\(32 to 47), X"000" & X"1") & \$18981_res\ & eclat_true & 
                  work.Int.sub(\$18977_binop_int6434365_arg\(80 to 95), X"000" & X"1") & \$18977_binop_int6434365_arg\(96 to 151) & \$18977_binop_int6434365_arg\(152 to 153);
                  result4928 := \$18977_binop_int6434365_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"a" =>
                  \$18981_res\ := work.Int.asr(\$18977_binop_int6434365_arg\(48 to 78), \$18980_v\(0 to 30));
                  \$18977_binop_int6434365_result\ := work.Int.add(\$18977_binop_int6434365_arg\(32 to 47), X"000" & X"1") & \$18981_res\ & eclat_true & 
                  work.Int.sub(\$18977_binop_int6434365_arg\(80 to 95), X"000" & X"1") & \$18977_binop_int6434365_arg\(96 to 151) & \$18977_binop_int6434365_arg\(152 to 153);
                  result4928 := \$18977_binop_int6434365_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"b" =>
                  \$18981_res\ := eclat_if(work.Int.lt(\$18977_binop_int6434365_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$18980_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.gt(\$18977_binop_int6434365_arg\(48 to 78), \$18980_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$18980_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"0" & 
                                  eclat_if(work.Int.lt(\$18977_binop_int6434365_arg\(48 to 78), \$18980_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$18977_binop_int6434365_result\ := work.Int.add(\$18977_binop_int6434365_arg\(32 to 47), X"000" & X"1") & \$18981_res\ & eclat_true & 
                  work.Int.sub(\$18977_binop_int6434365_arg\(80 to 95), X"000" & X"1") & \$18977_binop_int6434365_arg\(96 to 151) & \$18977_binop_int6434365_arg\(152 to 153);
                  result4928 := \$18977_binop_int6434365_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"c" =>
                  \$18981_res\ := eclat_if(work.Int.lt(\$18977_binop_int6434365_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$18980_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.le(\$18977_binop_int6434365_arg\(48 to 78), \$18980_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"1") & 
                                  eclat_if(work.Int.lt(\$18980_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & 
                                  eclat_if(work.Int.ge(\$18977_binop_int6434365_arg\(48 to 78), \$18980_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$18977_binop_int6434365_result\ := work.Int.add(\$18977_binop_int6434365_arg\(32 to 47), X"000" & X"1") & \$18981_res\ & eclat_true & 
                  work.Int.sub(\$18977_binop_int6434365_arg\(80 to 95), X"000" & X"1") & \$18977_binop_int6434365_arg\(96 to 151) & \$18977_binop_int6434365_arg\(152 to 153);
                  result4928 := \$18977_binop_int6434365_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when others =>
                  \$18981_res\ := "000"& X"000000" & X"0";
                  \$18977_binop_int6434365_result\ := work.Int.add(\$18977_binop_int6434365_arg\(32 to 47), X"000" & X"1") & \$18981_res\ & eclat_true & 
                  work.Int.sub(\$18977_binop_int6434365_arg\(80 to 95), X"000" & X"1") & \$18977_binop_int6434365_arg\(96 to 151) & \$18977_binop_int6434365_arg\(152 to 153);
                  result4928 := \$18977_binop_int6434365_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                end case;
              when PAUSE_GET5538 =>
                \$18999_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5537\ := \$18996_binop_int6434366_arg\(0 to 31);
                case \$v5537\ is
                when X"0000000" & X"0" =>
                  \$19000_res\ := work.Int.add(\$18996_binop_int6434366_arg\(48 to 78), \$18999_v\(0 to 30));
                  \$18996_binop_int6434366_result\ := work.Int.add(\$18996_binop_int6434366_arg\(32 to 47), X"000" & X"1") & \$19000_res\ & eclat_true & 
                  work.Int.sub(\$18996_binop_int6434366_arg\(80 to 95), X"000" & X"1") & \$18996_binop_int6434366_arg\(96 to 151) & \$18996_binop_int6434366_arg\(152 to 153);
                  result4928 := \$18996_binop_int6434366_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"1" =>
                  \$19000_res\ := work.Int.sub(\$18996_binop_int6434366_arg\(48 to 78), \$18999_v\(0 to 30));
                  \$18996_binop_int6434366_result\ := work.Int.add(\$18996_binop_int6434366_arg\(32 to 47), X"000" & X"1") & \$19000_res\ & eclat_true & 
                  work.Int.sub(\$18996_binop_int6434366_arg\(80 to 95), X"000" & X"1") & \$18996_binop_int6434366_arg\(96 to 151) & \$18996_binop_int6434366_arg\(152 to 153);
                  result4928 := \$18996_binop_int6434366_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"2" =>
                  \$19000_res\ := work.Int.mul(\$18996_binop_int6434366_arg\(48 to 78), \$18999_v\(0 to 30));
                  \$18996_binop_int6434366_result\ := work.Int.add(\$18996_binop_int6434366_arg\(32 to 47), X"000" & X"1") & \$19000_res\ & eclat_true & 
                  work.Int.sub(\$18996_binop_int6434366_arg\(80 to 95), X"000" & X"1") & \$18996_binop_int6434366_arg\(96 to 151) & \$18996_binop_int6434366_arg\(152 to 153);
                  result4928 := \$18996_binop_int6434366_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"3" =>
                  \$v5533\ := work.Int.eq(\$18999_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v5533\(0) = '1' then
                    \$19000_res\ := "000"& X"000000" & X"0";
                    \$18996_binop_int6434366_result\ := work.Int.add(
                                                        \$18996_binop_int6434366_arg\(32 to 47), X"000" & X"1") & \$19000_res\ & eclat_true & 
                    work.Int.sub(\$18996_binop_int6434366_arg\(80 to 95), X"000" & X"1") & \$18996_binop_int6434366_arg\(96 to 151) & \$18996_binop_int6434366_arg\(152 to 153);
                    result4928 := \$18996_binop_int6434366_result\;
                    rdy4929 := eclat_true;
                    state_var5920 := IDLE4930;
                  else
                    \$19002_modulo6684356_id\ := "000001011101";
                    \$19002_modulo6684356_arg\ := work.Int.absv(\$18996_binop_int6434366_arg\(48 to 78)) & 
                    work.Int.absv(\$18999_v\(0 to 30));
                    state_var5920 := \$19002_MODULO6684356\;
                  end if;
                when X"0000000" & X"4" =>
                  \$v5536\ := work.Int.eq(\$18999_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v5536\(0) = '1' then
                    \$19000_res\ := "000"& X"000000" & X"0";
                    \$18996_binop_int6434366_result\ := work.Int.add(
                                                        \$18996_binop_int6434366_arg\(32 to 47), X"000" & X"1") & \$19000_res\ & eclat_true & 
                    work.Int.sub(\$18996_binop_int6434366_arg\(80 to 95), X"000" & X"1") & \$18996_binop_int6434366_arg\(96 to 151) & \$18996_binop_int6434366_arg\(152 to 153);
                    result4928 := \$18996_binop_int6434366_result\;
                    rdy4929 := eclat_true;
                    state_var5920 := IDLE4930;
                  else
                    \$19009_modulo6684357_id\ := "000001011111";
                    \$19009_modulo6684357_arg\ := work.Int.absv(\$18996_binop_int6434366_arg\(48 to 78)) & 
                    work.Int.absv(\$18999_v\(0 to 30));
                    state_var5920 := \$19009_MODULO6684357\;
                  end if;
                when X"0000000" & X"5" =>
                  \$19000_res\ := work.Int.land(\$18996_binop_int6434366_arg\(48 to 78), \$18999_v\(0 to 30));
                  \$18996_binop_int6434366_result\ := work.Int.add(\$18996_binop_int6434366_arg\(32 to 47), X"000" & X"1") & \$19000_res\ & eclat_true & 
                  work.Int.sub(\$18996_binop_int6434366_arg\(80 to 95), X"000" & X"1") & \$18996_binop_int6434366_arg\(96 to 151) & \$18996_binop_int6434366_arg\(152 to 153);
                  result4928 := \$18996_binop_int6434366_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"6" =>
                  \$19000_res\ := work.Int.lor(\$18996_binop_int6434366_arg\(48 to 78), \$18999_v\(0 to 30));
                  \$18996_binop_int6434366_result\ := work.Int.add(\$18996_binop_int6434366_arg\(32 to 47), X"000" & X"1") & \$19000_res\ & eclat_true & 
                  work.Int.sub(\$18996_binop_int6434366_arg\(80 to 95), X"000" & X"1") & \$18996_binop_int6434366_arg\(96 to 151) & \$18996_binop_int6434366_arg\(152 to 153);
                  result4928 := \$18996_binop_int6434366_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"7" =>
                  \$19000_res\ := work.Int.lxor(\$18996_binop_int6434366_arg\(48 to 78), \$18999_v\(0 to 30));
                  \$18996_binop_int6434366_result\ := work.Int.add(\$18996_binop_int6434366_arg\(32 to 47), X"000" & X"1") & \$19000_res\ & eclat_true & 
                  work.Int.sub(\$18996_binop_int6434366_arg\(80 to 95), X"000" & X"1") & \$18996_binop_int6434366_arg\(96 to 151) & \$18996_binop_int6434366_arg\(152 to 153);
                  result4928 := \$18996_binop_int6434366_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"8" =>
                  \$19000_res\ := work.Int.lsl(\$18996_binop_int6434366_arg\(48 to 78), \$18999_v\(0 to 30));
                  \$18996_binop_int6434366_result\ := work.Int.add(\$18996_binop_int6434366_arg\(32 to 47), X"000" & X"1") & \$19000_res\ & eclat_true & 
                  work.Int.sub(\$18996_binop_int6434366_arg\(80 to 95), X"000" & X"1") & \$18996_binop_int6434366_arg\(96 to 151) & \$18996_binop_int6434366_arg\(152 to 153);
                  result4928 := \$18996_binop_int6434366_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"9" =>
                  \$19000_res\ := work.Int.lsr(\$18996_binop_int6434366_arg\(48 to 78), \$18999_v\(0 to 30));
                  \$18996_binop_int6434366_result\ := work.Int.add(\$18996_binop_int6434366_arg\(32 to 47), X"000" & X"1") & \$19000_res\ & eclat_true & 
                  work.Int.sub(\$18996_binop_int6434366_arg\(80 to 95), X"000" & X"1") & \$18996_binop_int6434366_arg\(96 to 151) & \$18996_binop_int6434366_arg\(152 to 153);
                  result4928 := \$18996_binop_int6434366_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"a" =>
                  \$19000_res\ := work.Int.asr(\$18996_binop_int6434366_arg\(48 to 78), \$18999_v\(0 to 30));
                  \$18996_binop_int6434366_result\ := work.Int.add(\$18996_binop_int6434366_arg\(32 to 47), X"000" & X"1") & \$19000_res\ & eclat_true & 
                  work.Int.sub(\$18996_binop_int6434366_arg\(80 to 95), X"000" & X"1") & \$18996_binop_int6434366_arg\(96 to 151) & \$18996_binop_int6434366_arg\(152 to 153);
                  result4928 := \$18996_binop_int6434366_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"b" =>
                  \$19000_res\ := eclat_if(work.Int.lt(\$18996_binop_int6434366_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$18999_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.gt(\$18996_binop_int6434366_arg\(48 to 78), \$18999_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$18999_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"0" & 
                                  eclat_if(work.Int.lt(\$18996_binop_int6434366_arg\(48 to 78), \$18999_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$18996_binop_int6434366_result\ := work.Int.add(\$18996_binop_int6434366_arg\(32 to 47), X"000" & X"1") & \$19000_res\ & eclat_true & 
                  work.Int.sub(\$18996_binop_int6434366_arg\(80 to 95), X"000" & X"1") & \$18996_binop_int6434366_arg\(96 to 151) & \$18996_binop_int6434366_arg\(152 to 153);
                  result4928 := \$18996_binop_int6434366_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"c" =>
                  \$19000_res\ := eclat_if(work.Int.lt(\$18996_binop_int6434366_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$18999_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.le(\$18996_binop_int6434366_arg\(48 to 78), \$18999_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"1") & 
                                  eclat_if(work.Int.lt(\$18999_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & 
                                  eclat_if(work.Int.ge(\$18996_binop_int6434366_arg\(48 to 78), \$18999_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$18996_binop_int6434366_result\ := work.Int.add(\$18996_binop_int6434366_arg\(32 to 47), X"000" & X"1") & \$19000_res\ & eclat_true & 
                  work.Int.sub(\$18996_binop_int6434366_arg\(80 to 95), X"000" & X"1") & \$18996_binop_int6434366_arg\(96 to 151) & \$18996_binop_int6434366_arg\(152 to 153);
                  result4928 := \$18996_binop_int6434366_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when others =>
                  \$19000_res\ := "000"& X"000000" & X"0";
                  \$18996_binop_int6434366_result\ := work.Int.add(\$18996_binop_int6434366_arg\(32 to 47), X"000" & X"1") & \$19000_res\ & eclat_true & 
                  work.Int.sub(\$18996_binop_int6434366_arg\(80 to 95), X"000" & X"1") & \$18996_binop_int6434366_arg\(96 to 151) & \$18996_binop_int6434366_arg\(152 to 153);
                  result4928 := \$18996_binop_int6434366_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                end case;
              when PAUSE_GET5548 =>
                \$19018_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5547\ := \$19015_binop_int6434367_arg\(0 to 31);
                case \$v5547\ is
                when X"0000000" & X"0" =>
                  \$19019_res\ := work.Int.add(\$19015_binop_int6434367_arg\(48 to 78), \$19018_v\(0 to 30));
                  \$19015_binop_int6434367_result\ := work.Int.add(\$19015_binop_int6434367_arg\(32 to 47), X"000" & X"1") & \$19019_res\ & eclat_true & 
                  work.Int.sub(\$19015_binop_int6434367_arg\(80 to 95), X"000" & X"1") & \$19015_binop_int6434367_arg\(96 to 151) & \$19015_binop_int6434367_arg\(152 to 153);
                  result4928 := \$19015_binop_int6434367_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"1" =>
                  \$19019_res\ := work.Int.sub(\$19015_binop_int6434367_arg\(48 to 78), \$19018_v\(0 to 30));
                  \$19015_binop_int6434367_result\ := work.Int.add(\$19015_binop_int6434367_arg\(32 to 47), X"000" & X"1") & \$19019_res\ & eclat_true & 
                  work.Int.sub(\$19015_binop_int6434367_arg\(80 to 95), X"000" & X"1") & \$19015_binop_int6434367_arg\(96 to 151) & \$19015_binop_int6434367_arg\(152 to 153);
                  result4928 := \$19015_binop_int6434367_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"2" =>
                  \$19019_res\ := work.Int.mul(\$19015_binop_int6434367_arg\(48 to 78), \$19018_v\(0 to 30));
                  \$19015_binop_int6434367_result\ := work.Int.add(\$19015_binop_int6434367_arg\(32 to 47), X"000" & X"1") & \$19019_res\ & eclat_true & 
                  work.Int.sub(\$19015_binop_int6434367_arg\(80 to 95), X"000" & X"1") & \$19015_binop_int6434367_arg\(96 to 151) & \$19015_binop_int6434367_arg\(152 to 153);
                  result4928 := \$19015_binop_int6434367_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"3" =>
                  \$v5543\ := work.Int.eq(\$19018_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v5543\(0) = '1' then
                    \$19019_res\ := "000"& X"000000" & X"0";
                    \$19015_binop_int6434367_result\ := work.Int.add(
                                                        \$19015_binop_int6434367_arg\(32 to 47), X"000" & X"1") & \$19019_res\ & eclat_true & 
                    work.Int.sub(\$19015_binop_int6434367_arg\(80 to 95), X"000" & X"1") & \$19015_binop_int6434367_arg\(96 to 151) & \$19015_binop_int6434367_arg\(152 to 153);
                    result4928 := \$19015_binop_int6434367_result\;
                    rdy4929 := eclat_true;
                    state_var5920 := IDLE4930;
                  else
                    \$19021_modulo6684356_id\ := "000001100010";
                    \$19021_modulo6684356_arg\ := work.Int.absv(\$19015_binop_int6434367_arg\(48 to 78)) & 
                    work.Int.absv(\$19018_v\(0 to 30));
                    state_var5920 := \$19021_MODULO6684356\;
                  end if;
                when X"0000000" & X"4" =>
                  \$v5546\ := work.Int.eq(\$19018_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v5546\(0) = '1' then
                    \$19019_res\ := "000"& X"000000" & X"0";
                    \$19015_binop_int6434367_result\ := work.Int.add(
                                                        \$19015_binop_int6434367_arg\(32 to 47), X"000" & X"1") & \$19019_res\ & eclat_true & 
                    work.Int.sub(\$19015_binop_int6434367_arg\(80 to 95), X"000" & X"1") & \$19015_binop_int6434367_arg\(96 to 151) & \$19015_binop_int6434367_arg\(152 to 153);
                    result4928 := \$19015_binop_int6434367_result\;
                    rdy4929 := eclat_true;
                    state_var5920 := IDLE4930;
                  else
                    \$19028_modulo6684357_id\ := "000001100100";
                    \$19028_modulo6684357_arg\ := work.Int.absv(\$19015_binop_int6434367_arg\(48 to 78)) & 
                    work.Int.absv(\$19018_v\(0 to 30));
                    state_var5920 := \$19028_MODULO6684357\;
                  end if;
                when X"0000000" & X"5" =>
                  \$19019_res\ := work.Int.land(\$19015_binop_int6434367_arg\(48 to 78), \$19018_v\(0 to 30));
                  \$19015_binop_int6434367_result\ := work.Int.add(\$19015_binop_int6434367_arg\(32 to 47), X"000" & X"1") & \$19019_res\ & eclat_true & 
                  work.Int.sub(\$19015_binop_int6434367_arg\(80 to 95), X"000" & X"1") & \$19015_binop_int6434367_arg\(96 to 151) & \$19015_binop_int6434367_arg\(152 to 153);
                  result4928 := \$19015_binop_int6434367_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"6" =>
                  \$19019_res\ := work.Int.lor(\$19015_binop_int6434367_arg\(48 to 78), \$19018_v\(0 to 30));
                  \$19015_binop_int6434367_result\ := work.Int.add(\$19015_binop_int6434367_arg\(32 to 47), X"000" & X"1") & \$19019_res\ & eclat_true & 
                  work.Int.sub(\$19015_binop_int6434367_arg\(80 to 95), X"000" & X"1") & \$19015_binop_int6434367_arg\(96 to 151) & \$19015_binop_int6434367_arg\(152 to 153);
                  result4928 := \$19015_binop_int6434367_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"7" =>
                  \$19019_res\ := work.Int.lxor(\$19015_binop_int6434367_arg\(48 to 78), \$19018_v\(0 to 30));
                  \$19015_binop_int6434367_result\ := work.Int.add(\$19015_binop_int6434367_arg\(32 to 47), X"000" & X"1") & \$19019_res\ & eclat_true & 
                  work.Int.sub(\$19015_binop_int6434367_arg\(80 to 95), X"000" & X"1") & \$19015_binop_int6434367_arg\(96 to 151) & \$19015_binop_int6434367_arg\(152 to 153);
                  result4928 := \$19015_binop_int6434367_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"8" =>
                  \$19019_res\ := work.Int.lsl(\$19015_binop_int6434367_arg\(48 to 78), \$19018_v\(0 to 30));
                  \$19015_binop_int6434367_result\ := work.Int.add(\$19015_binop_int6434367_arg\(32 to 47), X"000" & X"1") & \$19019_res\ & eclat_true & 
                  work.Int.sub(\$19015_binop_int6434367_arg\(80 to 95), X"000" & X"1") & \$19015_binop_int6434367_arg\(96 to 151) & \$19015_binop_int6434367_arg\(152 to 153);
                  result4928 := \$19015_binop_int6434367_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"9" =>
                  \$19019_res\ := work.Int.lsr(\$19015_binop_int6434367_arg\(48 to 78), \$19018_v\(0 to 30));
                  \$19015_binop_int6434367_result\ := work.Int.add(\$19015_binop_int6434367_arg\(32 to 47), X"000" & X"1") & \$19019_res\ & eclat_true & 
                  work.Int.sub(\$19015_binop_int6434367_arg\(80 to 95), X"000" & X"1") & \$19015_binop_int6434367_arg\(96 to 151) & \$19015_binop_int6434367_arg\(152 to 153);
                  result4928 := \$19015_binop_int6434367_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"a" =>
                  \$19019_res\ := work.Int.asr(\$19015_binop_int6434367_arg\(48 to 78), \$19018_v\(0 to 30));
                  \$19015_binop_int6434367_result\ := work.Int.add(\$19015_binop_int6434367_arg\(32 to 47), X"000" & X"1") & \$19019_res\ & eclat_true & 
                  work.Int.sub(\$19015_binop_int6434367_arg\(80 to 95), X"000" & X"1") & \$19015_binop_int6434367_arg\(96 to 151) & \$19015_binop_int6434367_arg\(152 to 153);
                  result4928 := \$19015_binop_int6434367_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"b" =>
                  \$19019_res\ := eclat_if(work.Int.lt(\$19015_binop_int6434367_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$19018_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.gt(\$19015_binop_int6434367_arg\(48 to 78), \$19018_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$19018_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"0" & 
                                  eclat_if(work.Int.lt(\$19015_binop_int6434367_arg\(48 to 78), \$19018_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$19015_binop_int6434367_result\ := work.Int.add(\$19015_binop_int6434367_arg\(32 to 47), X"000" & X"1") & \$19019_res\ & eclat_true & 
                  work.Int.sub(\$19015_binop_int6434367_arg\(80 to 95), X"000" & X"1") & \$19015_binop_int6434367_arg\(96 to 151) & \$19015_binop_int6434367_arg\(152 to 153);
                  result4928 := \$19015_binop_int6434367_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"c" =>
                  \$19019_res\ := eclat_if(work.Int.lt(\$19015_binop_int6434367_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$19018_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.le(\$19015_binop_int6434367_arg\(48 to 78), \$19018_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"1") & 
                                  eclat_if(work.Int.lt(\$19018_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & 
                                  eclat_if(work.Int.ge(\$19015_binop_int6434367_arg\(48 to 78), \$19018_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$19015_binop_int6434367_result\ := work.Int.add(\$19015_binop_int6434367_arg\(32 to 47), X"000" & X"1") & \$19019_res\ & eclat_true & 
                  work.Int.sub(\$19015_binop_int6434367_arg\(80 to 95), X"000" & X"1") & \$19015_binop_int6434367_arg\(96 to 151) & \$19015_binop_int6434367_arg\(152 to 153);
                  result4928 := \$19015_binop_int6434367_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when others =>
                  \$19019_res\ := "000"& X"000000" & X"0";
                  \$19015_binop_int6434367_result\ := work.Int.add(\$19015_binop_int6434367_arg\(32 to 47), X"000" & X"1") & \$19019_res\ & eclat_true & 
                  work.Int.sub(\$19015_binop_int6434367_arg\(80 to 95), X"000" & X"1") & \$19015_binop_int6434367_arg\(96 to 151) & \$19015_binop_int6434367_arg\(152 to 153);
                  result4928 := \$19015_binop_int6434367_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                end case;
              when PAUSE_GET5558 =>
                \$19037_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5557\ := \$19034_binop_int6434368_arg\(0 to 31);
                case \$v5557\ is
                when X"0000000" & X"0" =>
                  \$19038_res\ := work.Int.add(\$19034_binop_int6434368_arg\(48 to 78), \$19037_v\(0 to 30));
                  \$19034_binop_int6434368_result\ := work.Int.add(\$19034_binop_int6434368_arg\(32 to 47), X"000" & X"1") & \$19038_res\ & eclat_true & 
                  work.Int.sub(\$19034_binop_int6434368_arg\(80 to 95), X"000" & X"1") & \$19034_binop_int6434368_arg\(96 to 151) & \$19034_binop_int6434368_arg\(152 to 153);
                  result4928 := \$19034_binop_int6434368_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"1" =>
                  \$19038_res\ := work.Int.sub(\$19034_binop_int6434368_arg\(48 to 78), \$19037_v\(0 to 30));
                  \$19034_binop_int6434368_result\ := work.Int.add(\$19034_binop_int6434368_arg\(32 to 47), X"000" & X"1") & \$19038_res\ & eclat_true & 
                  work.Int.sub(\$19034_binop_int6434368_arg\(80 to 95), X"000" & X"1") & \$19034_binop_int6434368_arg\(96 to 151) & \$19034_binop_int6434368_arg\(152 to 153);
                  result4928 := \$19034_binop_int6434368_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"2" =>
                  \$19038_res\ := work.Int.mul(\$19034_binop_int6434368_arg\(48 to 78), \$19037_v\(0 to 30));
                  \$19034_binop_int6434368_result\ := work.Int.add(\$19034_binop_int6434368_arg\(32 to 47), X"000" & X"1") & \$19038_res\ & eclat_true & 
                  work.Int.sub(\$19034_binop_int6434368_arg\(80 to 95), X"000" & X"1") & \$19034_binop_int6434368_arg\(96 to 151) & \$19034_binop_int6434368_arg\(152 to 153);
                  result4928 := \$19034_binop_int6434368_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"3" =>
                  \$v5553\ := work.Int.eq(\$19037_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v5553\(0) = '1' then
                    \$19038_res\ := "000"& X"000000" & X"0";
                    \$19034_binop_int6434368_result\ := work.Int.add(
                                                        \$19034_binop_int6434368_arg\(32 to 47), X"000" & X"1") & \$19038_res\ & eclat_true & 
                    work.Int.sub(\$19034_binop_int6434368_arg\(80 to 95), X"000" & X"1") & \$19034_binop_int6434368_arg\(96 to 151) & \$19034_binop_int6434368_arg\(152 to 153);
                    result4928 := \$19034_binop_int6434368_result\;
                    rdy4929 := eclat_true;
                    state_var5920 := IDLE4930;
                  else
                    \$19040_modulo6684356_id\ := "000001100111";
                    \$19040_modulo6684356_arg\ := work.Int.absv(\$19034_binop_int6434368_arg\(48 to 78)) & 
                    work.Int.absv(\$19037_v\(0 to 30));
                    state_var5920 := \$19040_MODULO6684356\;
                  end if;
                when X"0000000" & X"4" =>
                  \$v5556\ := work.Int.eq(\$19037_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v5556\(0) = '1' then
                    \$19038_res\ := "000"& X"000000" & X"0";
                    \$19034_binop_int6434368_result\ := work.Int.add(
                                                        \$19034_binop_int6434368_arg\(32 to 47), X"000" & X"1") & \$19038_res\ & eclat_true & 
                    work.Int.sub(\$19034_binop_int6434368_arg\(80 to 95), X"000" & X"1") & \$19034_binop_int6434368_arg\(96 to 151) & \$19034_binop_int6434368_arg\(152 to 153);
                    result4928 := \$19034_binop_int6434368_result\;
                    rdy4929 := eclat_true;
                    state_var5920 := IDLE4930;
                  else
                    \$19047_modulo6684357_id\ := "000001101001";
                    \$19047_modulo6684357_arg\ := work.Int.absv(\$19034_binop_int6434368_arg\(48 to 78)) & 
                    work.Int.absv(\$19037_v\(0 to 30));
                    state_var5920 := \$19047_MODULO6684357\;
                  end if;
                when X"0000000" & X"5" =>
                  \$19038_res\ := work.Int.land(\$19034_binop_int6434368_arg\(48 to 78), \$19037_v\(0 to 30));
                  \$19034_binop_int6434368_result\ := work.Int.add(\$19034_binop_int6434368_arg\(32 to 47), X"000" & X"1") & \$19038_res\ & eclat_true & 
                  work.Int.sub(\$19034_binop_int6434368_arg\(80 to 95), X"000" & X"1") & \$19034_binop_int6434368_arg\(96 to 151) & \$19034_binop_int6434368_arg\(152 to 153);
                  result4928 := \$19034_binop_int6434368_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"6" =>
                  \$19038_res\ := work.Int.lor(\$19034_binop_int6434368_arg\(48 to 78), \$19037_v\(0 to 30));
                  \$19034_binop_int6434368_result\ := work.Int.add(\$19034_binop_int6434368_arg\(32 to 47), X"000" & X"1") & \$19038_res\ & eclat_true & 
                  work.Int.sub(\$19034_binop_int6434368_arg\(80 to 95), X"000" & X"1") & \$19034_binop_int6434368_arg\(96 to 151) & \$19034_binop_int6434368_arg\(152 to 153);
                  result4928 := \$19034_binop_int6434368_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"7" =>
                  \$19038_res\ := work.Int.lxor(\$19034_binop_int6434368_arg\(48 to 78), \$19037_v\(0 to 30));
                  \$19034_binop_int6434368_result\ := work.Int.add(\$19034_binop_int6434368_arg\(32 to 47), X"000" & X"1") & \$19038_res\ & eclat_true & 
                  work.Int.sub(\$19034_binop_int6434368_arg\(80 to 95), X"000" & X"1") & \$19034_binop_int6434368_arg\(96 to 151) & \$19034_binop_int6434368_arg\(152 to 153);
                  result4928 := \$19034_binop_int6434368_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"8" =>
                  \$19038_res\ := work.Int.lsl(\$19034_binop_int6434368_arg\(48 to 78), \$19037_v\(0 to 30));
                  \$19034_binop_int6434368_result\ := work.Int.add(\$19034_binop_int6434368_arg\(32 to 47), X"000" & X"1") & \$19038_res\ & eclat_true & 
                  work.Int.sub(\$19034_binop_int6434368_arg\(80 to 95), X"000" & X"1") & \$19034_binop_int6434368_arg\(96 to 151) & \$19034_binop_int6434368_arg\(152 to 153);
                  result4928 := \$19034_binop_int6434368_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"9" =>
                  \$19038_res\ := work.Int.lsr(\$19034_binop_int6434368_arg\(48 to 78), \$19037_v\(0 to 30));
                  \$19034_binop_int6434368_result\ := work.Int.add(\$19034_binop_int6434368_arg\(32 to 47), X"000" & X"1") & \$19038_res\ & eclat_true & 
                  work.Int.sub(\$19034_binop_int6434368_arg\(80 to 95), X"000" & X"1") & \$19034_binop_int6434368_arg\(96 to 151) & \$19034_binop_int6434368_arg\(152 to 153);
                  result4928 := \$19034_binop_int6434368_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"a" =>
                  \$19038_res\ := work.Int.asr(\$19034_binop_int6434368_arg\(48 to 78), \$19037_v\(0 to 30));
                  \$19034_binop_int6434368_result\ := work.Int.add(\$19034_binop_int6434368_arg\(32 to 47), X"000" & X"1") & \$19038_res\ & eclat_true & 
                  work.Int.sub(\$19034_binop_int6434368_arg\(80 to 95), X"000" & X"1") & \$19034_binop_int6434368_arg\(96 to 151) & \$19034_binop_int6434368_arg\(152 to 153);
                  result4928 := \$19034_binop_int6434368_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"b" =>
                  \$19038_res\ := eclat_if(work.Int.lt(\$19034_binop_int6434368_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$19037_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.gt(\$19034_binop_int6434368_arg\(48 to 78), \$19037_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$19037_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"0" & 
                                  eclat_if(work.Int.lt(\$19034_binop_int6434368_arg\(48 to 78), \$19037_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$19034_binop_int6434368_result\ := work.Int.add(\$19034_binop_int6434368_arg\(32 to 47), X"000" & X"1") & \$19038_res\ & eclat_true & 
                  work.Int.sub(\$19034_binop_int6434368_arg\(80 to 95), X"000" & X"1") & \$19034_binop_int6434368_arg\(96 to 151) & \$19034_binop_int6434368_arg\(152 to 153);
                  result4928 := \$19034_binop_int6434368_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"c" =>
                  \$19038_res\ := eclat_if(work.Int.lt(\$19034_binop_int6434368_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$19037_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.le(\$19034_binop_int6434368_arg\(48 to 78), \$19037_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"1") & 
                                  eclat_if(work.Int.lt(\$19037_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & 
                                  eclat_if(work.Int.ge(\$19034_binop_int6434368_arg\(48 to 78), \$19037_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$19034_binop_int6434368_result\ := work.Int.add(\$19034_binop_int6434368_arg\(32 to 47), X"000" & X"1") & \$19038_res\ & eclat_true & 
                  work.Int.sub(\$19034_binop_int6434368_arg\(80 to 95), X"000" & X"1") & \$19034_binop_int6434368_arg\(96 to 151) & \$19034_binop_int6434368_arg\(152 to 153);
                  result4928 := \$19034_binop_int6434368_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when others =>
                  \$19038_res\ := "000"& X"000000" & X"0";
                  \$19034_binop_int6434368_result\ := work.Int.add(\$19034_binop_int6434368_arg\(32 to 47), X"000" & X"1") & \$19038_res\ & eclat_true & 
                  work.Int.sub(\$19034_binop_int6434368_arg\(80 to 95), X"000" & X"1") & \$19034_binop_int6434368_arg\(96 to 151) & \$19034_binop_int6434368_arg\(152 to 153);
                  result4928 := \$19034_binop_int6434368_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                end case;
              when PAUSE_GET5568 =>
                \$19056_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5567\ := \$19053_binop_int6434369_arg\(0 to 31);
                case \$v5567\ is
                when X"0000000" & X"0" =>
                  \$19057_res\ := work.Int.add(\$19053_binop_int6434369_arg\(48 to 78), \$19056_v\(0 to 30));
                  \$19053_binop_int6434369_result\ := work.Int.add(\$19053_binop_int6434369_arg\(32 to 47), X"000" & X"1") & \$19057_res\ & eclat_true & 
                  work.Int.sub(\$19053_binop_int6434369_arg\(80 to 95), X"000" & X"1") & \$19053_binop_int6434369_arg\(96 to 151) & \$19053_binop_int6434369_arg\(152 to 153);
                  result4928 := \$19053_binop_int6434369_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"1" =>
                  \$19057_res\ := work.Int.sub(\$19053_binop_int6434369_arg\(48 to 78), \$19056_v\(0 to 30));
                  \$19053_binop_int6434369_result\ := work.Int.add(\$19053_binop_int6434369_arg\(32 to 47), X"000" & X"1") & \$19057_res\ & eclat_true & 
                  work.Int.sub(\$19053_binop_int6434369_arg\(80 to 95), X"000" & X"1") & \$19053_binop_int6434369_arg\(96 to 151) & \$19053_binop_int6434369_arg\(152 to 153);
                  result4928 := \$19053_binop_int6434369_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"2" =>
                  \$19057_res\ := work.Int.mul(\$19053_binop_int6434369_arg\(48 to 78), \$19056_v\(0 to 30));
                  \$19053_binop_int6434369_result\ := work.Int.add(\$19053_binop_int6434369_arg\(32 to 47), X"000" & X"1") & \$19057_res\ & eclat_true & 
                  work.Int.sub(\$19053_binop_int6434369_arg\(80 to 95), X"000" & X"1") & \$19053_binop_int6434369_arg\(96 to 151) & \$19053_binop_int6434369_arg\(152 to 153);
                  result4928 := \$19053_binop_int6434369_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"3" =>
                  \$v5563\ := work.Int.eq(\$19056_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v5563\(0) = '1' then
                    \$19057_res\ := "000"& X"000000" & X"0";
                    \$19053_binop_int6434369_result\ := work.Int.add(
                                                        \$19053_binop_int6434369_arg\(32 to 47), X"000" & X"1") & \$19057_res\ & eclat_true & 
                    work.Int.sub(\$19053_binop_int6434369_arg\(80 to 95), X"000" & X"1") & \$19053_binop_int6434369_arg\(96 to 151) & \$19053_binop_int6434369_arg\(152 to 153);
                    result4928 := \$19053_binop_int6434369_result\;
                    rdy4929 := eclat_true;
                    state_var5920 := IDLE4930;
                  else
                    \$19059_modulo6684356_id\ := "000001101100";
                    \$19059_modulo6684356_arg\ := work.Int.absv(\$19053_binop_int6434369_arg\(48 to 78)) & 
                    work.Int.absv(\$19056_v\(0 to 30));
                    state_var5920 := \$19059_MODULO6684356\;
                  end if;
                when X"0000000" & X"4" =>
                  \$v5566\ := work.Int.eq(\$19056_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v5566\(0) = '1' then
                    \$19057_res\ := "000"& X"000000" & X"0";
                    \$19053_binop_int6434369_result\ := work.Int.add(
                                                        \$19053_binop_int6434369_arg\(32 to 47), X"000" & X"1") & \$19057_res\ & eclat_true & 
                    work.Int.sub(\$19053_binop_int6434369_arg\(80 to 95), X"000" & X"1") & \$19053_binop_int6434369_arg\(96 to 151) & \$19053_binop_int6434369_arg\(152 to 153);
                    result4928 := \$19053_binop_int6434369_result\;
                    rdy4929 := eclat_true;
                    state_var5920 := IDLE4930;
                  else
                    \$19066_modulo6684357_id\ := "000001101110";
                    \$19066_modulo6684357_arg\ := work.Int.absv(\$19053_binop_int6434369_arg\(48 to 78)) & 
                    work.Int.absv(\$19056_v\(0 to 30));
                    state_var5920 := \$19066_MODULO6684357\;
                  end if;
                when X"0000000" & X"5" =>
                  \$19057_res\ := work.Int.land(\$19053_binop_int6434369_arg\(48 to 78), \$19056_v\(0 to 30));
                  \$19053_binop_int6434369_result\ := work.Int.add(\$19053_binop_int6434369_arg\(32 to 47), X"000" & X"1") & \$19057_res\ & eclat_true & 
                  work.Int.sub(\$19053_binop_int6434369_arg\(80 to 95), X"000" & X"1") & \$19053_binop_int6434369_arg\(96 to 151) & \$19053_binop_int6434369_arg\(152 to 153);
                  result4928 := \$19053_binop_int6434369_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"6" =>
                  \$19057_res\ := work.Int.lor(\$19053_binop_int6434369_arg\(48 to 78), \$19056_v\(0 to 30));
                  \$19053_binop_int6434369_result\ := work.Int.add(\$19053_binop_int6434369_arg\(32 to 47), X"000" & X"1") & \$19057_res\ & eclat_true & 
                  work.Int.sub(\$19053_binop_int6434369_arg\(80 to 95), X"000" & X"1") & \$19053_binop_int6434369_arg\(96 to 151) & \$19053_binop_int6434369_arg\(152 to 153);
                  result4928 := \$19053_binop_int6434369_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"7" =>
                  \$19057_res\ := work.Int.lxor(\$19053_binop_int6434369_arg\(48 to 78), \$19056_v\(0 to 30));
                  \$19053_binop_int6434369_result\ := work.Int.add(\$19053_binop_int6434369_arg\(32 to 47), X"000" & X"1") & \$19057_res\ & eclat_true & 
                  work.Int.sub(\$19053_binop_int6434369_arg\(80 to 95), X"000" & X"1") & \$19053_binop_int6434369_arg\(96 to 151) & \$19053_binop_int6434369_arg\(152 to 153);
                  result4928 := \$19053_binop_int6434369_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"8" =>
                  \$19057_res\ := work.Int.lsl(\$19053_binop_int6434369_arg\(48 to 78), \$19056_v\(0 to 30));
                  \$19053_binop_int6434369_result\ := work.Int.add(\$19053_binop_int6434369_arg\(32 to 47), X"000" & X"1") & \$19057_res\ & eclat_true & 
                  work.Int.sub(\$19053_binop_int6434369_arg\(80 to 95), X"000" & X"1") & \$19053_binop_int6434369_arg\(96 to 151) & \$19053_binop_int6434369_arg\(152 to 153);
                  result4928 := \$19053_binop_int6434369_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"9" =>
                  \$19057_res\ := work.Int.lsr(\$19053_binop_int6434369_arg\(48 to 78), \$19056_v\(0 to 30));
                  \$19053_binop_int6434369_result\ := work.Int.add(\$19053_binop_int6434369_arg\(32 to 47), X"000" & X"1") & \$19057_res\ & eclat_true & 
                  work.Int.sub(\$19053_binop_int6434369_arg\(80 to 95), X"000" & X"1") & \$19053_binop_int6434369_arg\(96 to 151) & \$19053_binop_int6434369_arg\(152 to 153);
                  result4928 := \$19053_binop_int6434369_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"a" =>
                  \$19057_res\ := work.Int.asr(\$19053_binop_int6434369_arg\(48 to 78), \$19056_v\(0 to 30));
                  \$19053_binop_int6434369_result\ := work.Int.add(\$19053_binop_int6434369_arg\(32 to 47), X"000" & X"1") & \$19057_res\ & eclat_true & 
                  work.Int.sub(\$19053_binop_int6434369_arg\(80 to 95), X"000" & X"1") & \$19053_binop_int6434369_arg\(96 to 151) & \$19053_binop_int6434369_arg\(152 to 153);
                  result4928 := \$19053_binop_int6434369_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"b" =>
                  \$19057_res\ := eclat_if(work.Int.lt(\$19053_binop_int6434369_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$19056_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.gt(\$19053_binop_int6434369_arg\(48 to 78), \$19056_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$19056_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"0" & 
                                  eclat_if(work.Int.lt(\$19053_binop_int6434369_arg\(48 to 78), \$19056_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$19053_binop_int6434369_result\ := work.Int.add(\$19053_binop_int6434369_arg\(32 to 47), X"000" & X"1") & \$19057_res\ & eclat_true & 
                  work.Int.sub(\$19053_binop_int6434369_arg\(80 to 95), X"000" & X"1") & \$19053_binop_int6434369_arg\(96 to 151) & \$19053_binop_int6434369_arg\(152 to 153);
                  result4928 := \$19053_binop_int6434369_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"c" =>
                  \$19057_res\ := eclat_if(work.Int.lt(\$19053_binop_int6434369_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$19056_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.le(\$19053_binop_int6434369_arg\(48 to 78), \$19056_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"1") & 
                                  eclat_if(work.Int.lt(\$19056_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & 
                                  eclat_if(work.Int.ge(\$19053_binop_int6434369_arg\(48 to 78), \$19056_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$19053_binop_int6434369_result\ := work.Int.add(\$19053_binop_int6434369_arg\(32 to 47), X"000" & X"1") & \$19057_res\ & eclat_true & 
                  work.Int.sub(\$19053_binop_int6434369_arg\(80 to 95), X"000" & X"1") & \$19053_binop_int6434369_arg\(96 to 151) & \$19053_binop_int6434369_arg\(152 to 153);
                  result4928 := \$19053_binop_int6434369_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when others =>
                  \$19057_res\ := "000"& X"000000" & X"0";
                  \$19053_binop_int6434369_result\ := work.Int.add(\$19053_binop_int6434369_arg\(32 to 47), X"000" & X"1") & \$19057_res\ & eclat_true & 
                  work.Int.sub(\$19053_binop_int6434369_arg\(80 to 95), X"000" & X"1") & \$19053_binop_int6434369_arg\(96 to 151) & \$19053_binop_int6434369_arg\(152 to 153);
                  result4928 := \$19053_binop_int6434369_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                end case;
              when PAUSE_GET5578 =>
                \$19075_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5577\ := \$19072_binop_int6434370_arg\(0 to 31);
                case \$v5577\ is
                when X"0000000" & X"0" =>
                  \$19076_res\ := work.Int.add(\$19072_binop_int6434370_arg\(48 to 78), \$19075_v\(0 to 30));
                  \$19072_binop_int6434370_result\ := work.Int.add(\$19072_binop_int6434370_arg\(32 to 47), X"000" & X"1") & \$19076_res\ & eclat_true & 
                  work.Int.sub(\$19072_binop_int6434370_arg\(80 to 95), X"000" & X"1") & \$19072_binop_int6434370_arg\(96 to 151) & \$19072_binop_int6434370_arg\(152 to 153);
                  result4928 := \$19072_binop_int6434370_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"1" =>
                  \$19076_res\ := work.Int.sub(\$19072_binop_int6434370_arg\(48 to 78), \$19075_v\(0 to 30));
                  \$19072_binop_int6434370_result\ := work.Int.add(\$19072_binop_int6434370_arg\(32 to 47), X"000" & X"1") & \$19076_res\ & eclat_true & 
                  work.Int.sub(\$19072_binop_int6434370_arg\(80 to 95), X"000" & X"1") & \$19072_binop_int6434370_arg\(96 to 151) & \$19072_binop_int6434370_arg\(152 to 153);
                  result4928 := \$19072_binop_int6434370_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"2" =>
                  \$19076_res\ := work.Int.mul(\$19072_binop_int6434370_arg\(48 to 78), \$19075_v\(0 to 30));
                  \$19072_binop_int6434370_result\ := work.Int.add(\$19072_binop_int6434370_arg\(32 to 47), X"000" & X"1") & \$19076_res\ & eclat_true & 
                  work.Int.sub(\$19072_binop_int6434370_arg\(80 to 95), X"000" & X"1") & \$19072_binop_int6434370_arg\(96 to 151) & \$19072_binop_int6434370_arg\(152 to 153);
                  result4928 := \$19072_binop_int6434370_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"3" =>
                  \$v5573\ := work.Int.eq(\$19075_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v5573\(0) = '1' then
                    \$19076_res\ := "000"& X"000000" & X"0";
                    \$19072_binop_int6434370_result\ := work.Int.add(
                                                        \$19072_binop_int6434370_arg\(32 to 47), X"000" & X"1") & \$19076_res\ & eclat_true & 
                    work.Int.sub(\$19072_binop_int6434370_arg\(80 to 95), X"000" & X"1") & \$19072_binop_int6434370_arg\(96 to 151) & \$19072_binop_int6434370_arg\(152 to 153);
                    result4928 := \$19072_binop_int6434370_result\;
                    rdy4929 := eclat_true;
                    state_var5920 := IDLE4930;
                  else
                    \$19078_modulo6684356_id\ := "000001110001";
                    \$19078_modulo6684356_arg\ := work.Int.absv(\$19072_binop_int6434370_arg\(48 to 78)) & 
                    work.Int.absv(\$19075_v\(0 to 30));
                    state_var5920 := \$19078_MODULO6684356\;
                  end if;
                when X"0000000" & X"4" =>
                  \$v5576\ := work.Int.eq(\$19075_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v5576\(0) = '1' then
                    \$19076_res\ := "000"& X"000000" & X"0";
                    \$19072_binop_int6434370_result\ := work.Int.add(
                                                        \$19072_binop_int6434370_arg\(32 to 47), X"000" & X"1") & \$19076_res\ & eclat_true & 
                    work.Int.sub(\$19072_binop_int6434370_arg\(80 to 95), X"000" & X"1") & \$19072_binop_int6434370_arg\(96 to 151) & \$19072_binop_int6434370_arg\(152 to 153);
                    result4928 := \$19072_binop_int6434370_result\;
                    rdy4929 := eclat_true;
                    state_var5920 := IDLE4930;
                  else
                    \$19085_modulo6684357_id\ := "000001110011";
                    \$19085_modulo6684357_arg\ := work.Int.absv(\$19072_binop_int6434370_arg\(48 to 78)) & 
                    work.Int.absv(\$19075_v\(0 to 30));
                    state_var5920 := \$19085_MODULO6684357\;
                  end if;
                when X"0000000" & X"5" =>
                  \$19076_res\ := work.Int.land(\$19072_binop_int6434370_arg\(48 to 78), \$19075_v\(0 to 30));
                  \$19072_binop_int6434370_result\ := work.Int.add(\$19072_binop_int6434370_arg\(32 to 47), X"000" & X"1") & \$19076_res\ & eclat_true & 
                  work.Int.sub(\$19072_binop_int6434370_arg\(80 to 95), X"000" & X"1") & \$19072_binop_int6434370_arg\(96 to 151) & \$19072_binop_int6434370_arg\(152 to 153);
                  result4928 := \$19072_binop_int6434370_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"6" =>
                  \$19076_res\ := work.Int.lor(\$19072_binop_int6434370_arg\(48 to 78), \$19075_v\(0 to 30));
                  \$19072_binop_int6434370_result\ := work.Int.add(\$19072_binop_int6434370_arg\(32 to 47), X"000" & X"1") & \$19076_res\ & eclat_true & 
                  work.Int.sub(\$19072_binop_int6434370_arg\(80 to 95), X"000" & X"1") & \$19072_binop_int6434370_arg\(96 to 151) & \$19072_binop_int6434370_arg\(152 to 153);
                  result4928 := \$19072_binop_int6434370_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"7" =>
                  \$19076_res\ := work.Int.lxor(\$19072_binop_int6434370_arg\(48 to 78), \$19075_v\(0 to 30));
                  \$19072_binop_int6434370_result\ := work.Int.add(\$19072_binop_int6434370_arg\(32 to 47), X"000" & X"1") & \$19076_res\ & eclat_true & 
                  work.Int.sub(\$19072_binop_int6434370_arg\(80 to 95), X"000" & X"1") & \$19072_binop_int6434370_arg\(96 to 151) & \$19072_binop_int6434370_arg\(152 to 153);
                  result4928 := \$19072_binop_int6434370_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"8" =>
                  \$19076_res\ := work.Int.lsl(\$19072_binop_int6434370_arg\(48 to 78), \$19075_v\(0 to 30));
                  \$19072_binop_int6434370_result\ := work.Int.add(\$19072_binop_int6434370_arg\(32 to 47), X"000" & X"1") & \$19076_res\ & eclat_true & 
                  work.Int.sub(\$19072_binop_int6434370_arg\(80 to 95), X"000" & X"1") & \$19072_binop_int6434370_arg\(96 to 151) & \$19072_binop_int6434370_arg\(152 to 153);
                  result4928 := \$19072_binop_int6434370_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"9" =>
                  \$19076_res\ := work.Int.lsr(\$19072_binop_int6434370_arg\(48 to 78), \$19075_v\(0 to 30));
                  \$19072_binop_int6434370_result\ := work.Int.add(\$19072_binop_int6434370_arg\(32 to 47), X"000" & X"1") & \$19076_res\ & eclat_true & 
                  work.Int.sub(\$19072_binop_int6434370_arg\(80 to 95), X"000" & X"1") & \$19072_binop_int6434370_arg\(96 to 151) & \$19072_binop_int6434370_arg\(152 to 153);
                  result4928 := \$19072_binop_int6434370_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"a" =>
                  \$19076_res\ := work.Int.asr(\$19072_binop_int6434370_arg\(48 to 78), \$19075_v\(0 to 30));
                  \$19072_binop_int6434370_result\ := work.Int.add(\$19072_binop_int6434370_arg\(32 to 47), X"000" & X"1") & \$19076_res\ & eclat_true & 
                  work.Int.sub(\$19072_binop_int6434370_arg\(80 to 95), X"000" & X"1") & \$19072_binop_int6434370_arg\(96 to 151) & \$19072_binop_int6434370_arg\(152 to 153);
                  result4928 := \$19072_binop_int6434370_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"b" =>
                  \$19076_res\ := eclat_if(work.Int.lt(\$19072_binop_int6434370_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$19075_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.gt(\$19072_binop_int6434370_arg\(48 to 78), \$19075_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$19075_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"0" & 
                                  eclat_if(work.Int.lt(\$19072_binop_int6434370_arg\(48 to 78), \$19075_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$19072_binop_int6434370_result\ := work.Int.add(\$19072_binop_int6434370_arg\(32 to 47), X"000" & X"1") & \$19076_res\ & eclat_true & 
                  work.Int.sub(\$19072_binop_int6434370_arg\(80 to 95), X"000" & X"1") & \$19072_binop_int6434370_arg\(96 to 151) & \$19072_binop_int6434370_arg\(152 to 153);
                  result4928 := \$19072_binop_int6434370_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"c" =>
                  \$19076_res\ := eclat_if(work.Int.lt(\$19072_binop_int6434370_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$19075_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.le(\$19072_binop_int6434370_arg\(48 to 78), \$19075_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"1") & 
                                  eclat_if(work.Int.lt(\$19075_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & 
                                  eclat_if(work.Int.ge(\$19072_binop_int6434370_arg\(48 to 78), \$19075_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$19072_binop_int6434370_result\ := work.Int.add(\$19072_binop_int6434370_arg\(32 to 47), X"000" & X"1") & \$19076_res\ & eclat_true & 
                  work.Int.sub(\$19072_binop_int6434370_arg\(80 to 95), X"000" & X"1") & \$19072_binop_int6434370_arg\(96 to 151) & \$19072_binop_int6434370_arg\(152 to 153);
                  result4928 := \$19072_binop_int6434370_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when others =>
                  \$19076_res\ := "000"& X"000000" & X"0";
                  \$19072_binop_int6434370_result\ := work.Int.add(\$19072_binop_int6434370_arg\(32 to 47), X"000" & X"1") & \$19076_res\ & eclat_true & 
                  work.Int.sub(\$19072_binop_int6434370_arg\(80 to 95), X"000" & X"1") & \$19072_binop_int6434370_arg\(96 to 151) & \$19072_binop_int6434370_arg\(152 to 153);
                  result4928 := \$19072_binop_int6434370_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                end case;
              when PAUSE_GET5588 =>
                \$19094_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5587\ := \$19091_binop_int6434371_arg\(0 to 31);
                case \$v5587\ is
                when X"0000000" & X"0" =>
                  \$19095_res\ := work.Int.add(\$19091_binop_int6434371_arg\(48 to 78), \$19094_v\(0 to 30));
                  \$19091_binop_int6434371_result\ := work.Int.add(\$19091_binop_int6434371_arg\(32 to 47), X"000" & X"1") & \$19095_res\ & eclat_true & 
                  work.Int.sub(\$19091_binop_int6434371_arg\(80 to 95), X"000" & X"1") & \$19091_binop_int6434371_arg\(96 to 151) & \$19091_binop_int6434371_arg\(152 to 153);
                  result4928 := \$19091_binop_int6434371_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"1" =>
                  \$19095_res\ := work.Int.sub(\$19091_binop_int6434371_arg\(48 to 78), \$19094_v\(0 to 30));
                  \$19091_binop_int6434371_result\ := work.Int.add(\$19091_binop_int6434371_arg\(32 to 47), X"000" & X"1") & \$19095_res\ & eclat_true & 
                  work.Int.sub(\$19091_binop_int6434371_arg\(80 to 95), X"000" & X"1") & \$19091_binop_int6434371_arg\(96 to 151) & \$19091_binop_int6434371_arg\(152 to 153);
                  result4928 := \$19091_binop_int6434371_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"2" =>
                  \$19095_res\ := work.Int.mul(\$19091_binop_int6434371_arg\(48 to 78), \$19094_v\(0 to 30));
                  \$19091_binop_int6434371_result\ := work.Int.add(\$19091_binop_int6434371_arg\(32 to 47), X"000" & X"1") & \$19095_res\ & eclat_true & 
                  work.Int.sub(\$19091_binop_int6434371_arg\(80 to 95), X"000" & X"1") & \$19091_binop_int6434371_arg\(96 to 151) & \$19091_binop_int6434371_arg\(152 to 153);
                  result4928 := \$19091_binop_int6434371_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"3" =>
                  \$v5583\ := work.Int.eq(\$19094_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v5583\(0) = '1' then
                    \$19095_res\ := "000"& X"000000" & X"0";
                    \$19091_binop_int6434371_result\ := work.Int.add(
                                                        \$19091_binop_int6434371_arg\(32 to 47), X"000" & X"1") & \$19095_res\ & eclat_true & 
                    work.Int.sub(\$19091_binop_int6434371_arg\(80 to 95), X"000" & X"1") & \$19091_binop_int6434371_arg\(96 to 151) & \$19091_binop_int6434371_arg\(152 to 153);
                    result4928 := \$19091_binop_int6434371_result\;
                    rdy4929 := eclat_true;
                    state_var5920 := IDLE4930;
                  else
                    \$19097_modulo6684356_id\ := "000001110110";
                    \$19097_modulo6684356_arg\ := work.Int.absv(\$19091_binop_int6434371_arg\(48 to 78)) & 
                    work.Int.absv(\$19094_v\(0 to 30));
                    state_var5920 := \$19097_MODULO6684356\;
                  end if;
                when X"0000000" & X"4" =>
                  \$v5586\ := work.Int.eq(\$19094_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v5586\(0) = '1' then
                    \$19095_res\ := "000"& X"000000" & X"0";
                    \$19091_binop_int6434371_result\ := work.Int.add(
                                                        \$19091_binop_int6434371_arg\(32 to 47), X"000" & X"1") & \$19095_res\ & eclat_true & 
                    work.Int.sub(\$19091_binop_int6434371_arg\(80 to 95), X"000" & X"1") & \$19091_binop_int6434371_arg\(96 to 151) & \$19091_binop_int6434371_arg\(152 to 153);
                    result4928 := \$19091_binop_int6434371_result\;
                    rdy4929 := eclat_true;
                    state_var5920 := IDLE4930;
                  else
                    \$19104_modulo6684357_id\ := "000001111000";
                    \$19104_modulo6684357_arg\ := work.Int.absv(\$19091_binop_int6434371_arg\(48 to 78)) & 
                    work.Int.absv(\$19094_v\(0 to 30));
                    state_var5920 := \$19104_MODULO6684357\;
                  end if;
                when X"0000000" & X"5" =>
                  \$19095_res\ := work.Int.land(\$19091_binop_int6434371_arg\(48 to 78), \$19094_v\(0 to 30));
                  \$19091_binop_int6434371_result\ := work.Int.add(\$19091_binop_int6434371_arg\(32 to 47), X"000" & X"1") & \$19095_res\ & eclat_true & 
                  work.Int.sub(\$19091_binop_int6434371_arg\(80 to 95), X"000" & X"1") & \$19091_binop_int6434371_arg\(96 to 151) & \$19091_binop_int6434371_arg\(152 to 153);
                  result4928 := \$19091_binop_int6434371_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"6" =>
                  \$19095_res\ := work.Int.lor(\$19091_binop_int6434371_arg\(48 to 78), \$19094_v\(0 to 30));
                  \$19091_binop_int6434371_result\ := work.Int.add(\$19091_binop_int6434371_arg\(32 to 47), X"000" & X"1") & \$19095_res\ & eclat_true & 
                  work.Int.sub(\$19091_binop_int6434371_arg\(80 to 95), X"000" & X"1") & \$19091_binop_int6434371_arg\(96 to 151) & \$19091_binop_int6434371_arg\(152 to 153);
                  result4928 := \$19091_binop_int6434371_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"7" =>
                  \$19095_res\ := work.Int.lxor(\$19091_binop_int6434371_arg\(48 to 78), \$19094_v\(0 to 30));
                  \$19091_binop_int6434371_result\ := work.Int.add(\$19091_binop_int6434371_arg\(32 to 47), X"000" & X"1") & \$19095_res\ & eclat_true & 
                  work.Int.sub(\$19091_binop_int6434371_arg\(80 to 95), X"000" & X"1") & \$19091_binop_int6434371_arg\(96 to 151) & \$19091_binop_int6434371_arg\(152 to 153);
                  result4928 := \$19091_binop_int6434371_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"8" =>
                  \$19095_res\ := work.Int.lsl(\$19091_binop_int6434371_arg\(48 to 78), \$19094_v\(0 to 30));
                  \$19091_binop_int6434371_result\ := work.Int.add(\$19091_binop_int6434371_arg\(32 to 47), X"000" & X"1") & \$19095_res\ & eclat_true & 
                  work.Int.sub(\$19091_binop_int6434371_arg\(80 to 95), X"000" & X"1") & \$19091_binop_int6434371_arg\(96 to 151) & \$19091_binop_int6434371_arg\(152 to 153);
                  result4928 := \$19091_binop_int6434371_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"9" =>
                  \$19095_res\ := work.Int.lsr(\$19091_binop_int6434371_arg\(48 to 78), \$19094_v\(0 to 30));
                  \$19091_binop_int6434371_result\ := work.Int.add(\$19091_binop_int6434371_arg\(32 to 47), X"000" & X"1") & \$19095_res\ & eclat_true & 
                  work.Int.sub(\$19091_binop_int6434371_arg\(80 to 95), X"000" & X"1") & \$19091_binop_int6434371_arg\(96 to 151) & \$19091_binop_int6434371_arg\(152 to 153);
                  result4928 := \$19091_binop_int6434371_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"a" =>
                  \$19095_res\ := work.Int.asr(\$19091_binop_int6434371_arg\(48 to 78), \$19094_v\(0 to 30));
                  \$19091_binop_int6434371_result\ := work.Int.add(\$19091_binop_int6434371_arg\(32 to 47), X"000" & X"1") & \$19095_res\ & eclat_true & 
                  work.Int.sub(\$19091_binop_int6434371_arg\(80 to 95), X"000" & X"1") & \$19091_binop_int6434371_arg\(96 to 151) & \$19091_binop_int6434371_arg\(152 to 153);
                  result4928 := \$19091_binop_int6434371_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"b" =>
                  \$19095_res\ := eclat_if(work.Int.lt(\$19091_binop_int6434371_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$19094_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.gt(\$19091_binop_int6434371_arg\(48 to 78), \$19094_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$19094_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"0" & 
                                  eclat_if(work.Int.lt(\$19091_binop_int6434371_arg\(48 to 78), \$19094_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$19091_binop_int6434371_result\ := work.Int.add(\$19091_binop_int6434371_arg\(32 to 47), X"000" & X"1") & \$19095_res\ & eclat_true & 
                  work.Int.sub(\$19091_binop_int6434371_arg\(80 to 95), X"000" & X"1") & \$19091_binop_int6434371_arg\(96 to 151) & \$19091_binop_int6434371_arg\(152 to 153);
                  result4928 := \$19091_binop_int6434371_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"c" =>
                  \$19095_res\ := eclat_if(work.Int.lt(\$19091_binop_int6434371_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$19094_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.le(\$19091_binop_int6434371_arg\(48 to 78), \$19094_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"1") & 
                                  eclat_if(work.Int.lt(\$19094_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & 
                                  eclat_if(work.Int.ge(\$19091_binop_int6434371_arg\(48 to 78), \$19094_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$19091_binop_int6434371_result\ := work.Int.add(\$19091_binop_int6434371_arg\(32 to 47), X"000" & X"1") & \$19095_res\ & eclat_true & 
                  work.Int.sub(\$19091_binop_int6434371_arg\(80 to 95), X"000" & X"1") & \$19091_binop_int6434371_arg\(96 to 151) & \$19091_binop_int6434371_arg\(152 to 153);
                  result4928 := \$19091_binop_int6434371_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when others =>
                  \$19095_res\ := "000"& X"000000" & X"0";
                  \$19091_binop_int6434371_result\ := work.Int.add(\$19091_binop_int6434371_arg\(32 to 47), X"000" & X"1") & \$19095_res\ & eclat_true & 
                  work.Int.sub(\$19091_binop_int6434371_arg\(80 to 95), X"000" & X"1") & \$19091_binop_int6434371_arg\(96 to 151) & \$19091_binop_int6434371_arg\(152 to 153);
                  result4928 := \$19091_binop_int6434371_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                end case;
              when PAUSE_GET5598 =>
                \$19119_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5597\ := \$19116_binop_int6434373_arg\(0 to 31);
                case \$v5597\ is
                when X"0000000" & X"0" =>
                  \$19120_res\ := work.Int.add(\$19116_binop_int6434373_arg\(48 to 78), \$19119_v\(0 to 30));
                  \$19116_binop_int6434373_result\ := work.Int.add(\$19116_binop_int6434373_arg\(32 to 47), X"000" & X"1") & \$19120_res\ & eclat_true & 
                  work.Int.sub(\$19116_binop_int6434373_arg\(80 to 95), X"000" & X"1") & \$19116_binop_int6434373_arg\(96 to 151) & \$19116_binop_int6434373_arg\(152 to 153);
                  result4928 := \$19116_binop_int6434373_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"1" =>
                  \$19120_res\ := work.Int.sub(\$19116_binop_int6434373_arg\(48 to 78), \$19119_v\(0 to 30));
                  \$19116_binop_int6434373_result\ := work.Int.add(\$19116_binop_int6434373_arg\(32 to 47), X"000" & X"1") & \$19120_res\ & eclat_true & 
                  work.Int.sub(\$19116_binop_int6434373_arg\(80 to 95), X"000" & X"1") & \$19116_binop_int6434373_arg\(96 to 151) & \$19116_binop_int6434373_arg\(152 to 153);
                  result4928 := \$19116_binop_int6434373_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"2" =>
                  \$19120_res\ := work.Int.mul(\$19116_binop_int6434373_arg\(48 to 78), \$19119_v\(0 to 30));
                  \$19116_binop_int6434373_result\ := work.Int.add(\$19116_binop_int6434373_arg\(32 to 47), X"000" & X"1") & \$19120_res\ & eclat_true & 
                  work.Int.sub(\$19116_binop_int6434373_arg\(80 to 95), X"000" & X"1") & \$19116_binop_int6434373_arg\(96 to 151) & \$19116_binop_int6434373_arg\(152 to 153);
                  result4928 := \$19116_binop_int6434373_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"3" =>
                  \$v5593\ := work.Int.eq(\$19119_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v5593\(0) = '1' then
                    \$19120_res\ := "000"& X"000000" & X"0";
                    \$19116_binop_int6434373_result\ := work.Int.add(
                                                        \$19116_binop_int6434373_arg\(32 to 47), X"000" & X"1") & \$19120_res\ & eclat_true & 
                    work.Int.sub(\$19116_binop_int6434373_arg\(80 to 95), X"000" & X"1") & \$19116_binop_int6434373_arg\(96 to 151) & \$19116_binop_int6434373_arg\(152 to 153);
                    result4928 := \$19116_binop_int6434373_result\;
                    rdy4929 := eclat_true;
                    state_var5920 := IDLE4930;
                  else
                    \$19122_modulo6684356_id\ := "000001111100";
                    \$19122_modulo6684356_arg\ := work.Int.absv(\$19116_binop_int6434373_arg\(48 to 78)) & 
                    work.Int.absv(\$19119_v\(0 to 30));
                    state_var5920 := \$19122_MODULO6684356\;
                  end if;
                when X"0000000" & X"4" =>
                  \$v5596\ := work.Int.eq(\$19119_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v5596\(0) = '1' then
                    \$19120_res\ := "000"& X"000000" & X"0";
                    \$19116_binop_int6434373_result\ := work.Int.add(
                                                        \$19116_binop_int6434373_arg\(32 to 47), X"000" & X"1") & \$19120_res\ & eclat_true & 
                    work.Int.sub(\$19116_binop_int6434373_arg\(80 to 95), X"000" & X"1") & \$19116_binop_int6434373_arg\(96 to 151) & \$19116_binop_int6434373_arg\(152 to 153);
                    result4928 := \$19116_binop_int6434373_result\;
                    rdy4929 := eclat_true;
                    state_var5920 := IDLE4930;
                  else
                    \$19129_modulo6684357_id\ := "000001111110";
                    \$19129_modulo6684357_arg\ := work.Int.absv(\$19116_binop_int6434373_arg\(48 to 78)) & 
                    work.Int.absv(\$19119_v\(0 to 30));
                    state_var5920 := \$19129_MODULO6684357\;
                  end if;
                when X"0000000" & X"5" =>
                  \$19120_res\ := work.Int.land(\$19116_binop_int6434373_arg\(48 to 78), \$19119_v\(0 to 30));
                  \$19116_binop_int6434373_result\ := work.Int.add(\$19116_binop_int6434373_arg\(32 to 47), X"000" & X"1") & \$19120_res\ & eclat_true & 
                  work.Int.sub(\$19116_binop_int6434373_arg\(80 to 95), X"000" & X"1") & \$19116_binop_int6434373_arg\(96 to 151) & \$19116_binop_int6434373_arg\(152 to 153);
                  result4928 := \$19116_binop_int6434373_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"6" =>
                  \$19120_res\ := work.Int.lor(\$19116_binop_int6434373_arg\(48 to 78), \$19119_v\(0 to 30));
                  \$19116_binop_int6434373_result\ := work.Int.add(\$19116_binop_int6434373_arg\(32 to 47), X"000" & X"1") & \$19120_res\ & eclat_true & 
                  work.Int.sub(\$19116_binop_int6434373_arg\(80 to 95), X"000" & X"1") & \$19116_binop_int6434373_arg\(96 to 151) & \$19116_binop_int6434373_arg\(152 to 153);
                  result4928 := \$19116_binop_int6434373_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"7" =>
                  \$19120_res\ := work.Int.lxor(\$19116_binop_int6434373_arg\(48 to 78), \$19119_v\(0 to 30));
                  \$19116_binop_int6434373_result\ := work.Int.add(\$19116_binop_int6434373_arg\(32 to 47), X"000" & X"1") & \$19120_res\ & eclat_true & 
                  work.Int.sub(\$19116_binop_int6434373_arg\(80 to 95), X"000" & X"1") & \$19116_binop_int6434373_arg\(96 to 151) & \$19116_binop_int6434373_arg\(152 to 153);
                  result4928 := \$19116_binop_int6434373_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"8" =>
                  \$19120_res\ := work.Int.lsl(\$19116_binop_int6434373_arg\(48 to 78), \$19119_v\(0 to 30));
                  \$19116_binop_int6434373_result\ := work.Int.add(\$19116_binop_int6434373_arg\(32 to 47), X"000" & X"1") & \$19120_res\ & eclat_true & 
                  work.Int.sub(\$19116_binop_int6434373_arg\(80 to 95), X"000" & X"1") & \$19116_binop_int6434373_arg\(96 to 151) & \$19116_binop_int6434373_arg\(152 to 153);
                  result4928 := \$19116_binop_int6434373_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"9" =>
                  \$19120_res\ := work.Int.lsr(\$19116_binop_int6434373_arg\(48 to 78), \$19119_v\(0 to 30));
                  \$19116_binop_int6434373_result\ := work.Int.add(\$19116_binop_int6434373_arg\(32 to 47), X"000" & X"1") & \$19120_res\ & eclat_true & 
                  work.Int.sub(\$19116_binop_int6434373_arg\(80 to 95), X"000" & X"1") & \$19116_binop_int6434373_arg\(96 to 151) & \$19116_binop_int6434373_arg\(152 to 153);
                  result4928 := \$19116_binop_int6434373_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"a" =>
                  \$19120_res\ := work.Int.asr(\$19116_binop_int6434373_arg\(48 to 78), \$19119_v\(0 to 30));
                  \$19116_binop_int6434373_result\ := work.Int.add(\$19116_binop_int6434373_arg\(32 to 47), X"000" & X"1") & \$19120_res\ & eclat_true & 
                  work.Int.sub(\$19116_binop_int6434373_arg\(80 to 95), X"000" & X"1") & \$19116_binop_int6434373_arg\(96 to 151) & \$19116_binop_int6434373_arg\(152 to 153);
                  result4928 := \$19116_binop_int6434373_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"b" =>
                  \$19120_res\ := eclat_if(work.Int.lt(\$19116_binop_int6434373_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$19119_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.gt(\$19116_binop_int6434373_arg\(48 to 78), \$19119_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$19119_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"0" & 
                                  eclat_if(work.Int.lt(\$19116_binop_int6434373_arg\(48 to 78), \$19119_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$19116_binop_int6434373_result\ := work.Int.add(\$19116_binop_int6434373_arg\(32 to 47), X"000" & X"1") & \$19120_res\ & eclat_true & 
                  work.Int.sub(\$19116_binop_int6434373_arg\(80 to 95), X"000" & X"1") & \$19116_binop_int6434373_arg\(96 to 151) & \$19116_binop_int6434373_arg\(152 to 153);
                  result4928 := \$19116_binop_int6434373_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"c" =>
                  \$19120_res\ := eclat_if(work.Int.lt(\$19116_binop_int6434373_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$19119_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.le(\$19116_binop_int6434373_arg\(48 to 78), \$19119_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"1") & 
                                  eclat_if(work.Int.lt(\$19119_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & 
                                  eclat_if(work.Int.ge(\$19116_binop_int6434373_arg\(48 to 78), \$19119_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$19116_binop_int6434373_result\ := work.Int.add(\$19116_binop_int6434373_arg\(32 to 47), X"000" & X"1") & \$19120_res\ & eclat_true & 
                  work.Int.sub(\$19116_binop_int6434373_arg\(80 to 95), X"000" & X"1") & \$19116_binop_int6434373_arg\(96 to 151) & \$19116_binop_int6434373_arg\(152 to 153);
                  result4928 := \$19116_binop_int6434373_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when others =>
                  \$19120_res\ := "000"& X"000000" & X"0";
                  \$19116_binop_int6434373_result\ := work.Int.add(\$19116_binop_int6434373_arg\(32 to 47), X"000" & X"1") & \$19120_res\ & eclat_true & 
                  work.Int.sub(\$19116_binop_int6434373_arg\(80 to 95), X"000" & X"1") & \$19116_binop_int6434373_arg\(96 to 151) & \$19116_binop_int6434373_arg\(152 to 153);
                  result4928 := \$19116_binop_int6434373_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                end case;
              when PAUSE_GET5608 =>
                \$19138_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5607\ := \$19135_binop_int6434374_arg\(0 to 31);
                case \$v5607\ is
                when X"0000000" & X"0" =>
                  \$19139_res\ := work.Int.add(\$19135_binop_int6434374_arg\(48 to 78), \$19138_v\(0 to 30));
                  \$19135_binop_int6434374_result\ := work.Int.add(\$19135_binop_int6434374_arg\(32 to 47), X"000" & X"1") & \$19139_res\ & eclat_true & 
                  work.Int.sub(\$19135_binop_int6434374_arg\(80 to 95), X"000" & X"1") & \$19135_binop_int6434374_arg\(96 to 151) & \$19135_binop_int6434374_arg\(152 to 153);
                  result4928 := \$19135_binop_int6434374_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"1" =>
                  \$19139_res\ := work.Int.sub(\$19135_binop_int6434374_arg\(48 to 78), \$19138_v\(0 to 30));
                  \$19135_binop_int6434374_result\ := work.Int.add(\$19135_binop_int6434374_arg\(32 to 47), X"000" & X"1") & \$19139_res\ & eclat_true & 
                  work.Int.sub(\$19135_binop_int6434374_arg\(80 to 95), X"000" & X"1") & \$19135_binop_int6434374_arg\(96 to 151) & \$19135_binop_int6434374_arg\(152 to 153);
                  result4928 := \$19135_binop_int6434374_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"2" =>
                  \$19139_res\ := work.Int.mul(\$19135_binop_int6434374_arg\(48 to 78), \$19138_v\(0 to 30));
                  \$19135_binop_int6434374_result\ := work.Int.add(\$19135_binop_int6434374_arg\(32 to 47), X"000" & X"1") & \$19139_res\ & eclat_true & 
                  work.Int.sub(\$19135_binop_int6434374_arg\(80 to 95), X"000" & X"1") & \$19135_binop_int6434374_arg\(96 to 151) & \$19135_binop_int6434374_arg\(152 to 153);
                  result4928 := \$19135_binop_int6434374_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"3" =>
                  \$v5603\ := work.Int.eq(\$19138_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v5603\(0) = '1' then
                    \$19139_res\ := "000"& X"000000" & X"0";
                    \$19135_binop_int6434374_result\ := work.Int.add(
                                                        \$19135_binop_int6434374_arg\(32 to 47), X"000" & X"1") & \$19139_res\ & eclat_true & 
                    work.Int.sub(\$19135_binop_int6434374_arg\(80 to 95), X"000" & X"1") & \$19135_binop_int6434374_arg\(96 to 151) & \$19135_binop_int6434374_arg\(152 to 153);
                    result4928 := \$19135_binop_int6434374_result\;
                    rdy4929 := eclat_true;
                    state_var5920 := IDLE4930;
                  else
                    \$19141_modulo6684356_id\ := "000010000001";
                    \$19141_modulo6684356_arg\ := work.Int.absv(\$19135_binop_int6434374_arg\(48 to 78)) & 
                    work.Int.absv(\$19138_v\(0 to 30));
                    state_var5920 := \$19141_MODULO6684356\;
                  end if;
                when X"0000000" & X"4" =>
                  \$v5606\ := work.Int.eq(\$19138_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v5606\(0) = '1' then
                    \$19139_res\ := "000"& X"000000" & X"0";
                    \$19135_binop_int6434374_result\ := work.Int.add(
                                                        \$19135_binop_int6434374_arg\(32 to 47), X"000" & X"1") & \$19139_res\ & eclat_true & 
                    work.Int.sub(\$19135_binop_int6434374_arg\(80 to 95), X"000" & X"1") & \$19135_binop_int6434374_arg\(96 to 151) & \$19135_binop_int6434374_arg\(152 to 153);
                    result4928 := \$19135_binop_int6434374_result\;
                    rdy4929 := eclat_true;
                    state_var5920 := IDLE4930;
                  else
                    \$19148_modulo6684357_id\ := "000010000011";
                    \$19148_modulo6684357_arg\ := work.Int.absv(\$19135_binop_int6434374_arg\(48 to 78)) & 
                    work.Int.absv(\$19138_v\(0 to 30));
                    state_var5920 := \$19148_MODULO6684357\;
                  end if;
                when X"0000000" & X"5" =>
                  \$19139_res\ := work.Int.land(\$19135_binop_int6434374_arg\(48 to 78), \$19138_v\(0 to 30));
                  \$19135_binop_int6434374_result\ := work.Int.add(\$19135_binop_int6434374_arg\(32 to 47), X"000" & X"1") & \$19139_res\ & eclat_true & 
                  work.Int.sub(\$19135_binop_int6434374_arg\(80 to 95), X"000" & X"1") & \$19135_binop_int6434374_arg\(96 to 151) & \$19135_binop_int6434374_arg\(152 to 153);
                  result4928 := \$19135_binop_int6434374_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"6" =>
                  \$19139_res\ := work.Int.lor(\$19135_binop_int6434374_arg\(48 to 78), \$19138_v\(0 to 30));
                  \$19135_binop_int6434374_result\ := work.Int.add(\$19135_binop_int6434374_arg\(32 to 47), X"000" & X"1") & \$19139_res\ & eclat_true & 
                  work.Int.sub(\$19135_binop_int6434374_arg\(80 to 95), X"000" & X"1") & \$19135_binop_int6434374_arg\(96 to 151) & \$19135_binop_int6434374_arg\(152 to 153);
                  result4928 := \$19135_binop_int6434374_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"7" =>
                  \$19139_res\ := work.Int.lxor(\$19135_binop_int6434374_arg\(48 to 78), \$19138_v\(0 to 30));
                  \$19135_binop_int6434374_result\ := work.Int.add(\$19135_binop_int6434374_arg\(32 to 47), X"000" & X"1") & \$19139_res\ & eclat_true & 
                  work.Int.sub(\$19135_binop_int6434374_arg\(80 to 95), X"000" & X"1") & \$19135_binop_int6434374_arg\(96 to 151) & \$19135_binop_int6434374_arg\(152 to 153);
                  result4928 := \$19135_binop_int6434374_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"8" =>
                  \$19139_res\ := work.Int.lsl(\$19135_binop_int6434374_arg\(48 to 78), \$19138_v\(0 to 30));
                  \$19135_binop_int6434374_result\ := work.Int.add(\$19135_binop_int6434374_arg\(32 to 47), X"000" & X"1") & \$19139_res\ & eclat_true & 
                  work.Int.sub(\$19135_binop_int6434374_arg\(80 to 95), X"000" & X"1") & \$19135_binop_int6434374_arg\(96 to 151) & \$19135_binop_int6434374_arg\(152 to 153);
                  result4928 := \$19135_binop_int6434374_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"9" =>
                  \$19139_res\ := work.Int.lsr(\$19135_binop_int6434374_arg\(48 to 78), \$19138_v\(0 to 30));
                  \$19135_binop_int6434374_result\ := work.Int.add(\$19135_binop_int6434374_arg\(32 to 47), X"000" & X"1") & \$19139_res\ & eclat_true & 
                  work.Int.sub(\$19135_binop_int6434374_arg\(80 to 95), X"000" & X"1") & \$19135_binop_int6434374_arg\(96 to 151) & \$19135_binop_int6434374_arg\(152 to 153);
                  result4928 := \$19135_binop_int6434374_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"a" =>
                  \$19139_res\ := work.Int.asr(\$19135_binop_int6434374_arg\(48 to 78), \$19138_v\(0 to 30));
                  \$19135_binop_int6434374_result\ := work.Int.add(\$19135_binop_int6434374_arg\(32 to 47), X"000" & X"1") & \$19139_res\ & eclat_true & 
                  work.Int.sub(\$19135_binop_int6434374_arg\(80 to 95), X"000" & X"1") & \$19135_binop_int6434374_arg\(96 to 151) & \$19135_binop_int6434374_arg\(152 to 153);
                  result4928 := \$19135_binop_int6434374_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"b" =>
                  \$19139_res\ := eclat_if(work.Int.lt(\$19135_binop_int6434374_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$19138_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.gt(\$19135_binop_int6434374_arg\(48 to 78), \$19138_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$19138_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"0" & 
                                  eclat_if(work.Int.lt(\$19135_binop_int6434374_arg\(48 to 78), \$19138_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$19135_binop_int6434374_result\ := work.Int.add(\$19135_binop_int6434374_arg\(32 to 47), X"000" & X"1") & \$19139_res\ & eclat_true & 
                  work.Int.sub(\$19135_binop_int6434374_arg\(80 to 95), X"000" & X"1") & \$19135_binop_int6434374_arg\(96 to 151) & \$19135_binop_int6434374_arg\(152 to 153);
                  result4928 := \$19135_binop_int6434374_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when X"0000000" & X"c" =>
                  \$19139_res\ := eclat_if(work.Int.lt(\$19135_binop_int6434374_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$19138_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.le(\$19135_binop_int6434374_arg\(48 to 78), \$19138_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"1") & 
                                  eclat_if(work.Int.lt(\$19138_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & 
                                  eclat_if(work.Int.ge(\$19135_binop_int6434374_arg\(48 to 78), \$19138_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$19135_binop_int6434374_result\ := work.Int.add(\$19135_binop_int6434374_arg\(32 to 47), X"000" & X"1") & \$19139_res\ & eclat_true & 
                  work.Int.sub(\$19135_binop_int6434374_arg\(80 to 95), X"000" & X"1") & \$19135_binop_int6434374_arg\(96 to 151) & \$19135_binop_int6434374_arg\(152 to 153);
                  result4928 := \$19135_binop_int6434374_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when others =>
                  \$19139_res\ := "000"& X"000000" & X"0";
                  \$19135_binop_int6434374_result\ := work.Int.add(\$19135_binop_int6434374_arg\(32 to 47), X"000" & X"1") & \$19139_res\ & eclat_true & 
                  work.Int.sub(\$19135_binop_int6434374_arg\(80 to 95), X"000" & X"1") & \$19135_binop_int6434374_arg\(96 to 151) & \$19135_binop_int6434374_arg\(152 to 153);
                  result4928 := \$19135_binop_int6434374_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                end case;
              when PAUSE_GET5612 =>
                \$19169_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$19171_compare6444358_id\ := "000010000111";
                \$19171_compare6444358_arg\ := \$19166_binop_compare6454377_arg\(0 to 31) & \$19166_binop_compare6454377_arg\(48 to 78) & \$19169_v\(0 to 30);
                state_var5920 := \$19171_COMPARE6444358\;
              when PAUSE_GET5616 =>
                \$19177_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$19179_compare6444358_id\ := "000010001001";
                \$19179_compare6444358_arg\ := \$19174_binop_compare6454378_arg\(0 to 31) & \$19174_binop_compare6454378_arg\(48 to 78) & \$19177_v\(0 to 30);
                state_var5920 := \$19179_COMPARE6444358\;
              when PAUSE_GET5620 =>
                \$19185_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$19187_compare6444358_id\ := "000010001011";
                \$19187_compare6444358_arg\ := \$19182_binop_compare6454379_arg\(0 to 31) & \$19182_binop_compare6454379_arg\(48 to 78) & \$19185_v\(0 to 30);
                state_var5920 := \$19187_COMPARE6444358\;
              when PAUSE_GET5624 =>
                \$19193_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$19195_compare6444358_id\ := "000010001101";
                \$19195_compare6444358_arg\ := \$19190_binop_compare6454380_arg\(0 to 31) & \$19190_binop_compare6454380_arg\(48 to 78) & \$19193_v\(0 to 30);
                state_var5920 := \$19195_COMPARE6444358\;
              when PAUSE_GET5628 =>
                \$19201_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$19203_compare6444358_id\ := "000010001111";
                \$19203_compare6444358_arg\ := \$19198_binop_compare6454381_arg\(0 to 31) & \$19198_binop_compare6454381_arg\(48 to 78) & \$19201_v\(0 to 30);
                state_var5920 := \$19203_COMPARE6444358\;
              when PAUSE_GET5632 =>
                \$19209_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$19211_compare6444358_id\ := "000010010001";
                \$19211_compare6444358_arg\ := \$19206_binop_compare6454382_arg\(0 to 31) & \$19206_binop_compare6454382_arg\(48 to 78) & \$19209_v\(0 to 30);
                state_var5920 := \$19211_COMPARE6444358\;
              when PAUSE_GET5635 =>
                \$19216_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$19216_v\ & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5638 =>
                \$19218_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"2") & \$19218_v\ & 
                work.Int.add(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5647 =>
                \$19220\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"2") & \$19220\ & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5650 =>
                \$19222\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"2") & \$19222\ & 
                work.Int.add(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5665 =>
                \$19226\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := eclat_resize(\$19226\(0 to 30),16) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(16 to 47) & 
                work.Int.sub(eclat_resize(\$19215_argument1\,8), "00000001") & \$18788\(104 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5668 =>
                \$19227\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := eclat_resize(\$19227\(0 to 30),16) & \$18788\(16 to 47) & 
                work.Int.sub(\$18788\(48 to 63), eclat_resize(\$19215_argument1\,16)) & \$18788\(16 to 47) & 
                work.Int.sub(\$18788\(96 to 103), "00000001") & \$18788\(104 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5671 =>
                \$19230_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := eclat_resize(\$19228_v\(0 to 30),16) & \$18788\(16 to 47) & 
                work.Int.sub(work.Int.sub(work.Int.sub(work.Int.sub(\$18788\(48 to 63), eclat_resize(\$19215_argument1\,16)), X"000" & X"1"), X"000" & X"1"), X"000" & X"1") & \$19229_v\ & eclat_resize(\$19230_v\(0 to 30),8) & \$18788\(104 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5674 =>
                \$19229_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5673\ := \$ram_lock\;
                if \$v5673\(0) = '1' then
                  state_var5920 := Q_WAIT5672;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$18788\(48 to 63), eclat_resize(\$19215_argument1\,16)), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5671;
                end if;
              when PAUSE_GET5677 =>
                \$19228_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5676\ := \$ram_lock\;
                if \$v5676\(0) = '1' then
                  state_var5920 := Q_WAIT5675;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$18788\(48 to 63), eclat_resize(\$19215_argument1\,16)), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5674;
                end if;
              when PAUSE_GET5681 =>
                \$19237_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := eclat_resize(\$19235_v\(0 to 30),16) & \$19231\(64 to 95) & 
                work.Int.sub(work.Int.sub(work.Int.sub(\$19234_sp\, X"000" & X"1"), X"000" & X"1"), X"000" & X"1") & \$19236_v\ & eclat_resize(\$19237_v\(0 to 30),8) & \$18788\(104 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5684 =>
                \$19236_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5683\ := \$ram_lock\;
                if \$v5683\(0) = '1' then
                  state_var5920 := Q_WAIT5682;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$19234_sp\, X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5681;
                end if;
              when PAUSE_GET5687 =>
                \$19235_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5686\ := \$ram_lock\;
                if \$v5686\(0) = '1' then
                  state_var5920 := Q_WAIT5685;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$19234_sp\, X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5684;
                end if;
              when PAUSE_GET5693 =>
                \$19241_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5692\ := \$ram_lock\;
                if \$v5692\(0) = '1' then
                  state_var5920 := Q_WAIT5691;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$19238_w6514383_arg\(32 to 62),16), eclat_resize(
                                                          work.Int.add(
                                                          \$19238_w6514383_arg\(0 to 7), "00000010"),16)), X"000" & X"1")));
                  \$ram_write\ <= \$19241_v\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5690;
                end if;
              when PAUSE_GET5707 =>
                \$19244_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"2") & \$19244_v\ & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5710 =>
                \$19246_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"2") & \$19246_v\ & 
                work.Int.add(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5722 =>
                \$19256_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"2") & \$19256_v\ & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5728 =>
                \$19257_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5727\ := \$ram_lock\;
                if \$v5727\(0) = '1' then
                  state_var5920 := Q_WAIT5726;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$18788\(16 to 46),16), eclat_resize(\$19215_argument1\,16)), X"000" & X"1")));
                  \$ram_write\ <= \$19257_v\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5725;
                end if;
              when PAUSE_GET5731 =>
                \$19266\ := \$code_value\;
                release(\$code_lock\);
                result4928 := work.Int.add(work.Int.add(\$18788\(0 to 15), X"000" & X"2"), eclat_resize(\$19266\,16)) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5734 =>
                \$19267_hd\ := \$ram_value\;
                release(\$ram_lock\);
                \$19265_ofs\ := work.Int.add(eclat_resize(\$19215_argument1\,16), 
                                             work.Int.lsr(eclat_resize(\$19267_hd\(0 to 30),16), X"000000" & X"18"));
                \$v5733\ := \$code_lock\;
                if \$v5733\(0) = '1' then
                  state_var5920 := Q_WAIT5732;
                else
                  acquire(\$code_lock\);
                  \$code_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                  \$18788\(0 to 15), X"000" & X"2"), \$19265_ofs\)));
                  state_var5920 := PAUSE_GET5731;
                end if;
              when PAUSE_GET5750 =>
                \$19274_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"2") & \$19273\(0 to 31) & 
                work.Int.sub(\$19273\(80 to 95), X"000" & X"1") & \$19274_v\ & \$19273\(128 to 135) & \$19273\(136 to 151) & \$19273\(152 to 153);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5757 =>
                \$19282_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"2") & \$19281\(0 to 31) & 
                work.Int.sub(\$19281\(80 to 95), X"000" & X"1") & \$19282_v\ & \$19281\(128 to 135) & \$19281\(136 to 151) & \$19281\(152 to 153);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5764 =>
                \$19279_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5763\ := \$ram_lock\;
                if \$v5763\(0) = '1' then
                  state_var5920 := Q_WAIT5762;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.sub(
                                                          \$18788\(48 to 63), X"000" & X"1")));
                  \$ram_write\ <= \$18788\(64 to 95); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5761;
                end if;
              when PAUSE_GET5767 =>
                \$19291_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"2") & \$19290\(0 to 31) & 
                work.Int.sub(\$19290\(80 to 95), X"000" & X"1") & \$19291_v\ & \$19290\(128 to 135) & \$19290\(136 to 151) & \$19290\(152 to 153);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5774 =>
                \$19288_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5773\ := \$ram_lock\;
                if \$v5773\(0) = '1' then
                  state_var5920 := Q_WAIT5772;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.sub(
                                                          work.Int.sub(
                                                          \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= \$18788\(64 to 95); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5771;
                end if;
              when PAUSE_GET5777 =>
                \$19287_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5776\ := \$ram_lock\;
                if \$v5776\(0) = '1' then
                  state_var5920 := Q_WAIT5775;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5774;
                end if;
              when PAUSE_GET5780 =>
                \$19301_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"2") & \$19300\(0 to 31) & 
                work.Int.sub(\$19300\(80 to 95), X"000" & X"1") & \$19301_v\ & \$19300\(128 to 135) & \$19300\(136 to 151) & \$19300\(152 to 153);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5787 =>
                \$19298_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5786\ := \$ram_lock\;
                if \$v5786\(0) = '1' then
                  state_var5920 := Q_WAIT5785;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.sub(
                                                          work.Int.sub(
                                                          work.Int.sub(
                                                          \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= \$18788\(64 to 95); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5784;
                end if;
              when PAUSE_GET5790 =>
                \$19297_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5789\ := \$ram_lock\;
                if \$v5789\(0) = '1' then
                  state_var5920 := Q_WAIT5788;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5787;
                end if;
              when PAUSE_GET5793 =>
                \$19296_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5792\ := \$ram_lock\;
                if \$v5792\(0) = '1' then
                  state_var5920 := Q_WAIT5791;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5790;
                end if;
              when PAUSE_GET5796 =>
                \$19312_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"2") & \$19311\(0 to 31) & 
                work.Int.sub(\$19311\(80 to 95), X"000" & X"1") & \$19312_v\ & \$19311\(128 to 135) & \$19311\(136 to 151) & \$19311\(152 to 153);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5803 =>
                \$19309_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5802\ := \$ram_lock\;
                if \$v5802\(0) = '1' then
                  state_var5920 := Q_WAIT5801;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.sub(
                                                          work.Int.sub(
                                                          work.Int.sub(
                                                          work.Int.sub(
                                                          \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= \$18788\(64 to 95); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5800;
                end if;
              when PAUSE_GET5806 =>
                \$19308_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5805\ := \$ram_lock\;
                if \$v5805\(0) = '1' then
                  state_var5920 := Q_WAIT5804;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5803;
                end if;
              when PAUSE_GET5809 =>
                \$19307_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5808\ := \$ram_lock\;
                if \$v5808\(0) = '1' then
                  state_var5920 := Q_WAIT5807;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5806;
                end if;
              when PAUSE_GET5812 =>
                \$19306_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5811\ := \$ram_lock\;
                if \$v5811\(0) = '1' then
                  state_var5920 := Q_WAIT5810;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5809;
                end if;
              when PAUSE_GET5821 =>
                \$19324_f0\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5820\ := \$ram_lock\;
                if \$v5820\(0) = '1' then
                  state_var5920 := Q_WAIT5819;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$18788\(16 to 46),16), X"000" & X"0"), X"000" & X"1")));
                  \$ram_write\ <= work.Int.add(\$19324_f0\(0 to 30), \$19215_argument1\) & eclat_true; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5818;
                end if;
              when PAUSE_GET5826 =>
                \$19342\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := eclat_resize(\$19342\(0 to 30),16) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(16 to 47) & 
                work.Int.sub(work.Int.add(\$18788\(96 to 103), eclat_resize(\$19215_argument1\,8)), "00000001") & \$18788\(104 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5832 =>
                \$19350_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5831\ := \$ram_lock\;
                if \$v5831\(0) = '1' then
                  state_var5920 := Q_WAIT5830;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$19347_fill6534389_arg\(48 to 78),16), \$19347_fill6534389_arg\(0 to 15)), X"000" & X"1")));
                  \$ram_write\ <= \$19350_v\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5829;
                end if;
              when PAUSE_GET5843 =>
                \$19354_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"3") & \$19354_v\ & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5846 =>
                \$19353\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5845\ := \$ram_lock\;
                if \$v5845\(0) = '1' then
                  state_var5920 := Q_WAIT5844;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$19353\(0 to 30),16), eclat_resize(\$19340_argument2\,16)), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5843;
                end if;
              when PAUSE_GET5849 =>
                \$19357_v\ := \$ram_value\;
                release(\$ram_lock\);
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"3") & \$19357_v\ & 
                work.Int.add(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5852 =>
                \$19356\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5851\ := \$ram_lock\;
                if \$v5851\(0) = '1' then
                  state_var5920 := Q_WAIT5850;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$19356\(0 to 30),16), eclat_resize(\$19340_argument2\,16)), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5849;
                end if;
              when PAUSE_GET5861 =>
                \$19364_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5860\ := \$ram_lock\;
                if \$v5860\(0) = '1' then
                  state_var5920 := Q_WAIT5859;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$19361_fill6544390_arg\(48 to 78),16), \$19361_fill6544390_arg\(0 to 15)), X"000" & X"1")));
                  \$ram_write\ <= \$19364_v\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5858;
                end if;
              when PAUSE_GET5884 =>
                \$19423_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v5883\ := \$ram_lock\;
                if \$v5883\(0) = '1' then
                  state_var5920 := Q_WAIT5882;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$19420_w06554397_arg\(64 to 94),16), 
                                                          work.Int.sub(
                                                          work.Int.add(
                                                          \$19420_w06554397_arg\(0 to 15), 
                                                          work.Int.mul(
                                                          X"000" & X"2", \$19420_w06554397_arg\(32 to 47))), X"000" & X"1")), X"000" & X"1")));
                  \$ram_write\ <= \$19423_v\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5881;
                end if;
              when PAUSE_GET5895 =>
                \$19427\ := \$code_value\;
                release(\$code_lock\);
                \$19428\ := work.Int.print(clk,\$19427\);
                \$19429\ := work.Print.print_newline(clk,eclat_unit);
                result4928 := \$18788\(0 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_GET5899 =>
                \$19408_argument3\ := \$code_value\;
                release(\$code_lock\);
                \$v5898\ := eclat_resize(\$18816\,8);
                case \$v5898\ is
                when "00101100" =>
                  \$v5894\ := work.Int.gt(eclat_resize(\$19340_argument2\,16), X"000" & X"0");
                  if \$v5894\(0) = '1' then
                    \$v5893\ := \$ram_lock\;
                    if \$v5893\(0) = '1' then
                      state_var5920 := Q_WAIT5892;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                      \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                      state_var5920 := PAUSE_SET5891;
                    end if;
                  else
                    \$19409_sp\ := \$18788\(48 to 63);
                    \$18793_make_block579_id\ := "000010111010";
                    \$18793_make_block579_arg\ := \$19409_sp\ & \$18788\(16 to 47) & \$18788\(64 to 95) & "11110111" & 
                    work.Int.add(work.Int.sub(work.Int.mul(X"000" & X"2", eclat_resize(\$19215_argument1\,16)), X"000" & X"1"), eclat_resize(\$19340_argument2\,16));
                    state_var5920 := \$18793_MAKE_BLOCK579\;
                  end if;
                when others =>
                  \$19426\ := work.Print.print_string(clk,of_string("unknown opcode : "));
                  \$v5897\ := \$code_lock\;
                  if \$v5897\(0) = '1' then
                    state_var5920 := Q_WAIT5896;
                  else
                    acquire(\$code_lock\);
                    \$code_ptr\ <= to_integer(unsigned(\$18788\(0 to 15)));
                    state_var5920 := PAUSE_GET5895;
                  end if;
                end case;
              when PAUSE_GET5903 =>
                \$19340_argument2\ := \$code_value\;
                release(\$code_lock\);
                \$v5902\ := eclat_resize(\$18816\,8);
                case \$v5902\ is
                when "00100100" =>
                  \$18798_w652_id\ := "000010100110";
                  \$18798_w652_arg\ := X"000" & X"1" & \$18788\(48 to 63) & eclat_resize(\$19215_argument1\,16) & eclat_resize(\$19340_argument2\,16);
                  state_var5920 := \$18798_W652\;
                when "00101011" =>
                  \$v5842\ := work.Int.gt(eclat_resize(\$19215_argument1\,16), X"000" & X"0");
                  if \$v5842\(0) = '1' then
                    \$v5841\ := \$ram_lock\;
                    if \$v5841\(0) = '1' then
                      state_var5920 := Q_WAIT5840;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                      \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                      state_var5920 := PAUSE_SET5839;
                    end if;
                  else
                    \$19343_sp\ := \$18788\(48 to 63);
                    \$18793_make_block579_id\ := "000010101000";
                    \$18793_make_block579_arg\ := \$19343_sp\ & \$18788\(16 to 47) & \$18788\(64 to 95) & "11110111" & 
                    work.Int.add(eclat_resize(\$19215_argument1\,16), X"000" & X"1");
                    state_var5920 := \$18793_MAKE_BLOCK579\;
                  end if;
                when "00110111" =>
                  \$v5848\ := \$ram_lock\;
                  if \$v5848\(0) = '1' then
                    state_var5920 := Q_WAIT5847;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(X"3e80", eclat_resize(\$19215_argument1\,16))));
                    state_var5920 := PAUSE_GET5846;
                  end if;
                when "00111000" =>
                  \$v5857\ := \$ram_lock\;
                  if \$v5857\(0) = '1' then
                    state_var5920 := Q_WAIT5856;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5855;
                  end if;
                when "00111110" =>
                  \$18793_make_block579_id\ := "000010101010";
                  \$18793_make_block579_arg\ := \$18788\(48 to 63) & \$18788\(16 to 47) & \$18788\(64 to 95) & eclat_resize(\$19340_argument2\,8) & eclat_resize(\$19215_argument1\,16);
                  state_var5920 := \$18793_MAKE_BLOCK579\;
                when "10000011" =>
                  \$19366_compbranch6504391_id\ := "000010101100";
                  \$19366_compbranch6504391_arg\ := X"0000000" & X"0" & \$19215_argument1\ & \$19340_argument2\ & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  state_var5920 := \$19366_COMPBRANCH6504391\;
                when "10000100" =>
                  \$19373_compbranch6504392_id\ := "000010101110";
                  \$19373_compbranch6504392_arg\ := X"0000000" & X"1" & \$19215_argument1\ & \$19340_argument2\ & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  state_var5920 := \$19373_COMPBRANCH6504392\;
                when "10000101" =>
                  \$19380_compbranch6504393_id\ := "000010110000";
                  \$19380_compbranch6504393_arg\ := X"0000000" & X"2" & \$19215_argument1\ & \$19340_argument2\ & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  state_var5920 := \$19380_COMPBRANCH6504393\;
                when "10000110" =>
                  \$19387_compbranch6504394_id\ := "000010110010";
                  \$19387_compbranch6504394_arg\ := X"0000000" & X"3" & \$19215_argument1\ & \$19340_argument2\ & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  state_var5920 := \$19387_COMPBRANCH6504394\;
                when "10000111" =>
                  \$19394_compbranch6504395_id\ := "000010110100";
                  \$19394_compbranch6504395_arg\ := X"0000000" & X"4" & \$19215_argument1\ & \$19340_argument2\ & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  state_var5920 := \$19394_COMPBRANCH6504395\;
                when "10001000" =>
                  \$19401_compbranch6504396_id\ := "000010110110";
                  \$19401_compbranch6504396_arg\ := X"0000000" & X"5" & \$19215_argument1\ & \$19340_argument2\ & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  state_var5920 := \$19401_COMPBRANCH6504396\;
                when others =>
                  \$v5901\ := \$code_lock\;
                  if \$v5901\(0) = '1' then
                    state_var5920 := Q_WAIT5900;
                  else
                    acquire(\$code_lock\);
                    \$code_ptr\ <= to_integer(unsigned(work.Int.add(\$18788\(0 to 15), X"000" & X"3")));
                    state_var5920 := PAUSE_GET5899;
                  end if;
                end case;
              when PAUSE_GET5907 =>
                \$19215_argument1\ := \$code_value\;
                release(\$code_lock\);
                \$v5906\ := eclat_resize(\$18816\,8);
                case \$v5906\ is
                when "00001000" =>
                  \$v5637\ := \$ram_lock\;
                  if \$v5637\(0) = '1' then
                    state_var5920 := Q_WAIT5636;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                   \$18788\(48 to 63), eclat_resize(\$19215_argument1\,16)), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5635;
                  end if;
                when "00010010" =>
                  \$v5643\ := \$ram_lock\;
                  if \$v5643\(0) = '1' then
                    state_var5920 := Q_WAIT5642;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5641;
                  end if;
                when "00010011" =>
                  result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"2") & \$18788\(16 to 47) & 
                  work.Int.sub(\$18788\(48 to 63), eclat_resize(\$19215_argument1\,16)) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when "00010100" =>
                  \$v5646\ := \$ram_lock\;
                  if \$v5646\(0) = '1' then
                    state_var5920 := Q_WAIT5645;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.sub(
                                                            work.Int.sub(
                                                            \$18788\(48 to 63), X"000" & X"1"), eclat_resize(\$19215_argument1\,16))));
                    \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5644;
                  end if;
                when "00011001" =>
                  \$v5649\ := \$ram_lock\;
                  if \$v5649\(0) = '1' then
                    state_var5920 := Q_WAIT5648;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$18788\(64 to 94),16), 
                                                                   work.Int.sub(
                                                                   eclat_resize(\$19215_argument1\,16), X"000" & X"1")), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5647;
                  end if;
                when "00011110" =>
                  \$v5655\ := \$ram_lock\;
                  if \$v5655\(0) = '1' then
                    state_var5920 := Q_WAIT5654;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5653;
                  end if;
                when "00011111" =>
                  \$v5664\ := \$ram_lock\;
                  if \$v5664\(0) = '1' then
                    state_var5920 := Q_WAIT5663;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= eclat_resize(\$18788\(96 to 103),31) & eclat_true; \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5662;
                  end if;
                when "00100000" =>
                  \$v5667\ := \$ram_lock\;
                  if \$v5667\(0) = '1' then
                    state_var5920 := Q_WAIT5666;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$18788\(16 to 46),16), X"000" & X"0"), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5665;
                  end if;
                when "00100101" =>
                  \$18794_apply638_id\ := "000010010011";
                  \$18794_apply638_arg\ := eclat_true & eclat_false & eclat_false & \$18788\(96 to 103) & eclat_true & eclat_resize(\$19215_argument1\,16) & X"000" & X"1" & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(120 to 121) & \$18788\(64 to 95) & \$18788\(96 to 103) & \$18788\(104 to 119);
                  state_var5920 := \$18794_APPLY638\;
                when "00100110" =>
                  \$18794_apply638_id\ := "000010010100";
                  \$18794_apply638_arg\ := eclat_true & eclat_true & eclat_false & 
                  work.Int.add(\$18788\(96 to 103), "00000001") & eclat_true & eclat_resize(\$19215_argument1\,16) & X"000" & X"2" & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(120 to 121) & \$18788\(64 to 95) & \$18788\(96 to 103) & \$18788\(104 to 119);
                  state_var5920 := \$18794_APPLY638\;
                when "00100111" =>
                  \$18794_apply638_id\ := "000010010101";
                  \$18794_apply638_arg\ := eclat_true & eclat_true & eclat_true & 
                  work.Int.add(\$18788\(96 to 103), "00000010") & eclat_true & eclat_resize(\$19215_argument1\,16) & X"000" & X"3" & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(120 to 121) & \$18788\(64 to 95) & \$18788\(96 to 103) & \$18788\(104 to 119);
                  state_var5920 := \$18794_APPLY638\;
                when "00101000" =>
                  \$v5680\ := work.Int.gt(\$18788\(96 to 103), "00000000");
                  if \$v5680\(0) = '1' then
                    \$v5670\ := \$ram_lock\;
                    if \$v5670\(0) = '1' then
                      state_var5920 := Q_WAIT5669;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                        work.Int.add(
                                                        eclat_resize(\$18788\(16 to 46),16), X"000" & X"0"), X"000" & X"1")));
                      state_var5920 := PAUSE_GET5668;
                    end if;
                  else
                    \$v5679\ := \$ram_lock\;
                    if \$v5679\(0) = '1' then
                      state_var5920 := Q_WAIT5678;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(
                                                        work.Int.sub(
                                                        \$18788\(48 to 63), eclat_resize(\$19215_argument1\,16)), X"000" & X"1")));
                      state_var5920 := PAUSE_GET5677;
                    end if;
                  end if;
                when "00101010" =>
                  \$v5703\ := work.Int.ge(\$18788\(96 to 103), eclat_resize(\$19215_argument1\,8));
                  if \$v5703\(0) = '1' then
                    result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"2") & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 95) & 
                    work.Int.sub(\$18788\(96 to 103), eclat_resize(\$19215_argument1\,8)) & \$18788\(104 to 119) & \$18788\(120 to 121);
                    rdy4929 := eclat_true;
                    state_var5920 := IDLE4930;
                  else
                    \$18793_make_block579_id\ := "000010010111";
                    \$18793_make_block579_arg\ := \$18788\(48 to 63) & \$18788\(16 to 47) & \$18788\(64 to 95) & "11110111" & eclat_resize(
                    work.Int.add(\$18788\(96 to 103), "00000011"),16);
                    state_var5920 := \$18793_MAKE_BLOCK579\;
                  end if;
                when "00110000" =>
                  \$18795_offsetclosure_n639_id\ := "000010011000";
                  \$18795_offsetclosure_n639_arg\ := work.Int.add(\$18788\(0 to 15), X"000" & X"2") & \$18788\(48 to 63) & eclat_resize(\$19215_argument1\,16) & \$18788\(64 to 119) & \$18788\(120 to 121) & \$18788\(64 to 95);
                  state_var5920 := \$18795_OFFSETCLOSURE_N639\;
                when "00110100" =>
                  \$v5706\ := \$ram_lock\;
                  if \$v5706\(0) = '1' then
                    state_var5920 := Q_WAIT5705;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5704;
                  end if;
                when "00110101" =>
                  \$v5709\ := \$ram_lock\;
                  if \$v5709\(0) = '1' then
                    state_var5920 := Q_WAIT5708;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(X"3e80", eclat_resize(\$19215_argument1\,16))));
                    state_var5920 := PAUSE_GET5707;
                  end if;
                when "00110110" =>
                  \$v5715\ := \$ram_lock\;
                  if \$v5715\(0) = '1' then
                    state_var5920 := Q_WAIT5714;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5713;
                  end if;
                when "00111001" =>
                  \$v5718\ := \$ram_lock\;
                  if \$v5718\(0) = '1' then
                    state_var5920 := Q_WAIT5717;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            X"3e80", eclat_resize(\$19215_argument1\,16))));
                    \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5716;
                  end if;
                when "00111011" =>
                  \$18796_make_block_n646_id\ := "000010011010";
                  \$18796_make_block_n646_arg\ := work.Int.add(\$18788\(0 to 15), X"000" & X"2") & \$18788\(48 to 63) & eclat_false & eclat_false & eclat_false & \$19215_argument1\ & X"000" & X"0" & \$18788\(16 to 47) & \$18788\(120 to 121) & \$18788\(64 to 95) & \$18788\(96 to 103) & \$18788\(104 to 119);
                  state_var5920 := \$18796_MAKE_BLOCK_N646\;
                when "00111101" =>
                  \$v5721\ := \$ram_lock\;
                  if \$v5721\(0) = '1' then
                    state_var5920 := Q_WAIT5720;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5719;
                  end if;
                when "00111111" =>
                  \$18796_make_block_n646_id\ := "000010011100";
                  \$18796_make_block_n646_arg\ := work.Int.add(\$18788\(0 to 15), X"000" & X"2") & \$18788\(48 to 63) & eclat_true & eclat_false & eclat_false & \$19215_argument1\ & X"000" & X"1" & \$18788\(16 to 47) & \$18788\(120 to 121) & \$18788\(64 to 95) & \$18788\(96 to 103) & \$18788\(104 to 119);
                  state_var5920 := \$18796_MAKE_BLOCK_N646\;
                when "01000000" =>
                  \$18796_make_block_n646_id\ := "000010011101";
                  \$18796_make_block_n646_arg\ := work.Int.add(\$18788\(0 to 15), X"000" & X"2") & \$18788\(48 to 63) & eclat_true & eclat_true & eclat_false & \$19215_argument1\ & X"000" & X"2" & \$18788\(16 to 47) & \$18788\(120 to 121) & \$18788\(64 to 95) & \$18788\(96 to 103) & \$18788\(104 to 119);
                  state_var5920 := \$18796_MAKE_BLOCK_N646\;
                when "01000001" =>
                  \$18796_make_block_n646_id\ := "000010011110";
                  \$18796_make_block_n646_arg\ := work.Int.add(\$18788\(0 to 15), X"000" & X"2") & \$18788\(48 to 63) & eclat_true & eclat_true & eclat_true & \$19215_argument1\ & X"000" & X"3" & \$18788\(16 to 47) & \$18788\(120 to 121) & \$18788\(64 to 95) & \$18788\(96 to 103) & \$18788\(104 to 119);
                  state_var5920 := \$18796_MAKE_BLOCK_N646\;
                when "01000010" =>
                  \$19249\ := work.Print.print_string(clk,of_string("fatal error: "));
                  \$19250\ := work.Print.print_string(clk,of_string("unsupported instruction SETFLOATFIELD"));
                  \$19251\ := work.Print.print_newline(clk,eclat_unit);
                  \$19252_forever6704384_id\ := "000010011111";
                  \$19252_forever6704384_arg\ := eclat_unit;
                  state_var5920 := \$19252_FOREVER6704384\;
                when "01000111" =>
                  \$19255\ := work.Assertion.ok(work.Bool.lnot(""&\$18788\(47)));
                  \$v5724\ := \$ram_lock\;
                  if \$v5724\(0) = '1' then
                    state_var5920 := Q_WAIT5723;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$18788\(16 to 46),16), eclat_resize(\$19215_argument1\,16)), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5722;
                  end if;
                when "01001101" =>
                  \$v5730\ := \$ram_lock\;
                  if \$v5730\(0) = '1' then
                    state_var5920 := Q_WAIT5729;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18788\(48 to 63), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5728;
                  end if;
                when "01001110" =>
                  \$19259\ := work.Print.print_string(clk,of_string("fatal error: "));
                  \$19260\ := work.Print.print_string(clk,of_string("unsupported instruction SETFLOATFIELD"));
                  \$19261\ := work.Print.print_newline(clk,eclat_unit);
                  \$19262_forever6704385_id\ := "000010100000";
                  \$19262_forever6704385_arg\ := eclat_unit;
                  state_var5920 := \$19262_FOREVER6704385\;
                when "01010111" =>
                  \$v5737\ := ""&\$18788\(47);
                  if \$v5737\(0) = '1' then
                    \$19265_ofs\ := eclat_resize(\$18788\(16 to 46),16);
                    \$v5733\ := \$code_lock\;
                    if \$v5733\(0) = '1' then
                      state_var5920 := Q_WAIT5732;
                    else
                      acquire(\$code_lock\);
                      \$code_ptr\ <= to_integer(unsigned(work.Int.add(
                                                         work.Int.add(
                                                         \$18788\(0 to 15), X"000" & X"2"), \$19265_ofs\)));
                      state_var5920 := PAUSE_GET5731;
                    end if;
                  else
                    \$v5736\ := \$ram_lock\;
                    if \$v5736\(0) = '1' then
                      state_var5920 := Q_WAIT5735;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18788\(16 to 46),16)));
                      state_var5920 := PAUSE_GET5734;
                    end if;
                  end if;
                when "01010100" =>
                  result4928 := work.Int.add(work.Int.add(\$18788\(0 to 15), X"000" & X"1"), eclat_resize(\$19215_argument1\,16)) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when "01011001" =>
                  \$v5749\ := \$ram_lock\;
                  if \$v5749\(0) = '1' then
                    state_var5920 := Q_WAIT5748;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= eclat_resize(\$18788\(96 to 103),31) & eclat_true; \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5747;
                  end if;
                when "01011100" =>
                  result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 95) & \$18788\(96 to 103) & \$18788\(104 to 119) & \$18788\(120 to 121);
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when "01011101" =>
                  \$v5756\ := \$ram_lock\;
                  if \$v5756\(0) = '1' then
                    state_var5920 := Q_WAIT5755;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= \$18788\(64 to 95); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5754;
                  end if;
                when "01011110" =>
                  \$v5766\ := \$ram_lock\;
                  if \$v5766\(0) = '1' then
                    state_var5920 := Q_WAIT5765;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18788\(48 to 63), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5764;
                  end if;
                when "01011111" =>
                  \$v5779\ := \$ram_lock\;
                  if \$v5779\(0) = '1' then
                    state_var5920 := Q_WAIT5778;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18788\(48 to 63), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5777;
                  end if;
                when "01100000" =>
                  \$v5795\ := \$ram_lock\;
                  if \$v5795\(0) = '1' then
                    state_var5920 := Q_WAIT5794;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18788\(48 to 63), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5793;
                  end if;
                when "01100001" =>
                  \$v5814\ := \$ram_lock\;
                  if \$v5814\(0) = '1' then
                    state_var5920 := Q_WAIT5813;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18788\(48 to 63), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5812;
                  end if;
                when "01100010" =>
                  \$19317\ := work.Print.print_string(clk,of_string("fatal error: "));
                  \$19318\ := work.Print.print_string(clk,of_string("unsupported instruction CALLN"));
                  \$19319\ := work.Print.print_newline(clk,eclat_unit);
                  \$19320_forever6704386_id\ := "000010100001";
                  \$19320_forever6704386_arg\ := eclat_unit;
                  state_var5920 := \$19320_FOREVER6704386\;
                when "01100111" =>
                  result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"2") & \$19215_argument1\ & eclat_true & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when "01101100" =>
                  \$v5817\ := \$ram_lock\;
                  if \$v5817\(0) = '1' then
                    state_var5920 := Q_WAIT5816;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5815;
                  end if;
                when "01111111" =>
                  result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"2") & 
                  work.Int.add(\$18788\(16 to 46), \$19215_argument1\) & eclat_true & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when "10000000" =>
                  \$v5823\ := \$ram_lock\;
                  if \$v5823\(0) = '1' then
                    state_var5920 := Q_WAIT5822;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$18788\(16 to 46),16), X"000" & X"0"), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5821;
                  end if;
                when "10001011" =>
                  \$19326_compbranch6504387_id\ := "000010100011";
                  \$19326_compbranch6504387_arg\ := X"0000000" & X"2" & \$19215_argument1\ & \$18788\(16 to 46) & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  state_var5920 := \$19326_COMPBRANCH6504387\;
                when "10001100" =>
                  \$19333_compbranch6504388_id\ := "000010100101";
                  \$19333_compbranch6504388_arg\ := X"0000000" & X"5" & \$19215_argument1\ & \$18788\(16 to 46) & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  state_var5920 := \$19333_COMPBRANCH6504388\;
                when others =>
                  \$v5905\ := \$code_lock\;
                  if \$v5905\(0) = '1' then
                    state_var5920 := Q_WAIT5904;
                  else
                    acquire(\$code_lock\);
                    \$code_ptr\ <= to_integer(unsigned(work.Int.add(\$18788\(0 to 15), X"000" & X"2")));
                    state_var5920 := PAUSE_GET5903;
                  end if;
                end case;
              when PAUSE_GET5911 =>
                \$18816\ := \$code_value\;
                release(\$code_lock\);
                \$v5910\ := eclat_resize(\$18816\,8);
                case \$v5910\ is
                when "00000000" =>
                  \$v5254\ := \$ram_lock\;
                  if \$v5254\(0) = '1' then
                    state_var5920 := Q_WAIT5253;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                   \$18788\(48 to 63), X"000" & X"0"), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5252;
                  end if;
                when "00000001" =>
                  \$v5257\ := \$ram_lock\;
                  if \$v5257\(0) = '1' then
                    state_var5920 := Q_WAIT5256;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                   \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5255;
                  end if;
                when "00000010" =>
                  \$v5260\ := \$ram_lock\;
                  if \$v5260\(0) = '1' then
                    state_var5920 := Q_WAIT5259;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                   \$18788\(48 to 63), X"000" & X"2"), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5258;
                  end if;
                when "00000011" =>
                  \$v5263\ := \$ram_lock\;
                  if \$v5263\(0) = '1' then
                    state_var5920 := Q_WAIT5262;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                   \$18788\(48 to 63), X"000" & X"3"), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5261;
                  end if;
                when "00000100" =>
                  \$v5266\ := \$ram_lock\;
                  if \$v5266\(0) = '1' then
                    state_var5920 := Q_WAIT5265;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                   \$18788\(48 to 63), X"000" & X"4"), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5264;
                  end if;
                when "00000101" =>
                  \$v5269\ := \$ram_lock\;
                  if \$v5269\(0) = '1' then
                    state_var5920 := Q_WAIT5268;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                   \$18788\(48 to 63), X"000" & X"5"), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5267;
                  end if;
                when "00000110" =>
                  \$v5272\ := \$ram_lock\;
                  if \$v5272\(0) = '1' then
                    state_var5920 := Q_WAIT5271;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                   \$18788\(48 to 63), X"000" & X"6"), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5270;
                  end if;
                when "00000111" =>
                  \$v5275\ := \$ram_lock\;
                  if \$v5275\(0) = '1' then
                    state_var5920 := Q_WAIT5274;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                   \$18788\(48 to 63), X"000" & X"7"), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5273;
                  end if;
                when "00001001" =>
                  \$v5278\ := \$ram_lock\;
                  if \$v5278\(0) = '1' then
                    state_var5920 := Q_WAIT5277;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5276;
                  end if;
                when "00001010" =>
                  \$v5281\ := \$ram_lock\;
                  if \$v5281\(0) = '1' then
                    state_var5920 := Q_WAIT5280;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5279;
                  end if;
                when "00001011" =>
                  \$v5287\ := \$ram_lock\;
                  if \$v5287\(0) = '1' then
                    state_var5920 := Q_WAIT5286;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5285;
                  end if;
                when "00001100" =>
                  \$v5293\ := \$ram_lock\;
                  if \$v5293\(0) = '1' then
                    state_var5920 := Q_WAIT5292;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5291;
                  end if;
                when "00001101" =>
                  \$v5299\ := \$ram_lock\;
                  if \$v5299\(0) = '1' then
                    state_var5920 := Q_WAIT5298;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5297;
                  end if;
                when "00001110" =>
                  \$v5305\ := \$ram_lock\;
                  if \$v5305\(0) = '1' then
                    state_var5920 := Q_WAIT5304;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5303;
                  end if;
                when "00001111" =>
                  \$v5311\ := \$ram_lock\;
                  if \$v5311\(0) = '1' then
                    state_var5920 := Q_WAIT5310;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5309;
                  end if;
                when "00010000" =>
                  \$v5317\ := \$ram_lock\;
                  if \$v5317\(0) = '1' then
                    state_var5920 := Q_WAIT5316;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5315;
                  end if;
                when "00010001" =>
                  \$v5323\ := \$ram_lock\;
                  if \$v5323\(0) = '1' then
                    state_var5920 := Q_WAIT5322;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5321;
                  end if;
                when "00010101" =>
                  \$v5326\ := \$ram_lock\;
                  if \$v5326\(0) = '1' then
                    state_var5920 := Q_WAIT5325;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$18788\(64 to 94),16), 
                                                                   work.Int.sub(
                                                                   X"000" & X"1", X"000" & X"1")), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5324;
                  end if;
                when "00010110" =>
                  \$v5329\ := \$ram_lock\;
                  if \$v5329\(0) = '1' then
                    state_var5920 := Q_WAIT5328;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$18788\(64 to 94),16), 
                                                                   work.Int.sub(
                                                                   X"000" & X"2", X"000" & X"1")), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5327;
                  end if;
                when "00010111" =>
                  \$v5332\ := \$ram_lock\;
                  if \$v5332\(0) = '1' then
                    state_var5920 := Q_WAIT5331;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$18788\(64 to 94),16), 
                                                                   work.Int.sub(
                                                                   X"000" & X"3", X"000" & X"1")), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5330;
                  end if;
                when "00011000" =>
                  \$v5335\ := \$ram_lock\;
                  if \$v5335\(0) = '1' then
                    state_var5920 := Q_WAIT5334;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$18788\(64 to 94),16), 
                                                                   work.Int.sub(
                                                                   X"000" & X"4", X"000" & X"1")), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5333;
                  end if;
                when "00011010" =>
                  \$v5341\ := \$ram_lock\;
                  if \$v5341\(0) = '1' then
                    state_var5920 := Q_WAIT5340;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5339;
                  end if;
                when "00011011" =>
                  \$v5347\ := \$ram_lock\;
                  if \$v5347\(0) = '1' then
                    state_var5920 := Q_WAIT5346;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5345;
                  end if;
                when "00011100" =>
                  \$v5353\ := \$ram_lock\;
                  if \$v5353\(0) = '1' then
                    state_var5920 := Q_WAIT5352;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5351;
                  end if;
                when "00011101" =>
                  \$v5359\ := \$ram_lock\;
                  if \$v5359\(0) = '1' then
                    state_var5920 := Q_WAIT5358;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5357;
                  end if;
                when "00100001" =>
                  \$18794_apply638_id\ := "000000110101";
                  \$18794_apply638_arg\ := eclat_true & eclat_false & eclat_false & "00000000" & eclat_false & X"000" & X"0" & X"000" & X"0" & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(120 to 121) & \$18788\(64 to 95) & \$18788\(96 to 103) & \$18788\(104 to 119);
                  state_var5920 := \$18794_APPLY638\;
                when "00100010" =>
                  \$18794_apply638_id\ := "000000110110";
                  \$18794_apply638_arg\ := eclat_true & eclat_true & eclat_false & "00000001" & eclat_false & X"000" & X"0" & X"000" & X"0" & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(120 to 121) & \$18788\(64 to 95) & \$18788\(96 to 103) & \$18788\(104 to 119);
                  state_var5920 := \$18794_APPLY638\;
                when "00100011" =>
                  \$18794_apply638_id\ := "000000110111";
                  \$18794_apply638_arg\ := eclat_true & eclat_true & eclat_true & "00000010" & eclat_false & X"000" & X"0" & X"000" & X"0" & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(120 to 121) & \$18788\(64 to 95) & \$18788\(96 to 103) & \$18788\(104 to 119);
                  state_var5920 := \$18794_APPLY638\;
                when "00101001" =>
                  \$v5372\ := \$ram_lock\;
                  if \$v5372\(0) = '1' then
                    state_var5920 := Q_WAIT5371;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18788\(64 to 94),16)));
                    state_var5920 := PAUSE_GET5370;
                  end if;
                when "00101101" =>
                  \$18795_offsetclosure_n639_id\ := "000000111001";
                  \$18795_offsetclosure_n639_arg\ := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18788\(48 to 63) & 
                  work.Int.neg(X"000" & X"2") & \$18788\(64 to 119) & \$18788\(120 to 121) & \$18788\(64 to 95);
                  state_var5920 := \$18795_OFFSETCLOSURE_N639\;
                when "00101110" =>
                  \$18795_offsetclosure_n639_id\ := "000000111010";
                  \$18795_offsetclosure_n639_arg\ := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18788\(48 to 63) & X"000" & X"0" & \$18788\(64 to 119) & \$18788\(120 to 121) & \$18788\(64 to 95);
                  state_var5920 := \$18795_OFFSETCLOSURE_N639\;
                when "00101111" =>
                  \$18795_offsetclosure_n639_id\ := "000000111011";
                  \$18795_offsetclosure_n639_arg\ := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18788\(48 to 63) & X"000" & X"2" & \$18788\(64 to 119) & \$18788\(120 to 121) & \$18788\(64 to 95);
                  state_var5920 := \$18795_OFFSETCLOSURE_N639\;
                when "00110001" =>
                  \$v5375\ := \$ram_lock\;
                  if \$v5375\(0) = '1' then
                    state_var5920 := Q_WAIT5374;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5373;
                  end if;
                when "00110010" =>
                  \$v5378\ := \$ram_lock\;
                  if \$v5378\(0) = '1' then
                    state_var5920 := Q_WAIT5377;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5376;
                  end if;
                when "00110011" =>
                  \$v5381\ := \$ram_lock\;
                  if \$v5381\(0) = '1' then
                    state_var5920 := Q_WAIT5380;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5379;
                  end if;
                when "00111010" =>
                  \$18796_make_block_n646_id\ := "000000111111";
                  \$18796_make_block_n646_arg\ := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18788\(48 to 63) & eclat_false & eclat_false & eclat_false & "000"& X"000000" & X"0" & X"000" & X"0" & \$18788\(16 to 47) & \$18788\(120 to 121) & \$18788\(64 to 95) & \$18788\(96 to 103) & \$18788\(104 to 119);
                  state_var5920 := \$18796_MAKE_BLOCK_N646\;
                when "00111100" =>
                  \$v5384\ := \$ram_lock\;
                  if \$v5384\(0) = '1' then
                    state_var5920 := Q_WAIT5383;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5382;
                  end if;
                when "01000011" =>
                  \$18865\ := work.Assertion.ok(work.Bool.lnot(""&\$18788\(47)));
                  \$v5387\ := \$ram_lock\;
                  if \$v5387\(0) = '1' then
                    state_var5920 := Q_WAIT5386;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$18788\(16 to 46),16), X"000" & X"0"), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5385;
                  end if;
                when "01000100" =>
                  \$18867\ := work.Assertion.ok(work.Bool.lnot(""&\$18788\(47)));
                  \$v5390\ := \$ram_lock\;
                  if \$v5390\(0) = '1' then
                    state_var5920 := Q_WAIT5389;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$18788\(16 to 46),16), X"000" & X"1"), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5388;
                  end if;
                when "01000101" =>
                  \$18869\ := work.Assertion.ok(work.Bool.lnot(""&\$18788\(47)));
                  \$v5393\ := \$ram_lock\;
                  if \$v5393\(0) = '1' then
                    state_var5920 := Q_WAIT5392;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$18788\(16 to 46),16), X"000" & X"2"), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5391;
                  end if;
                when "01000110" =>
                  \$18871\ := work.Assertion.ok(work.Bool.lnot(""&\$18788\(47)));
                  \$v5396\ := \$ram_lock\;
                  if \$v5396\(0) = '1' then
                    state_var5920 := Q_WAIT5395;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$18788\(16 to 46),16), X"000" & X"3"), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5394;
                  end if;
                when "01001001" =>
                  \$v5402\ := \$ram_lock\;
                  if \$v5402\(0) = '1' then
                    state_var5920 := Q_WAIT5401;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18788\(48 to 63), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5400;
                  end if;
                when "01001010" =>
                  \$v5408\ := \$ram_lock\;
                  if \$v5408\(0) = '1' then
                    state_var5920 := Q_WAIT5407;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18788\(48 to 63), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5406;
                  end if;
                when "01001011" =>
                  \$v5414\ := \$ram_lock\;
                  if \$v5414\(0) = '1' then
                    state_var5920 := Q_WAIT5413;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18788\(48 to 63), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5412;
                  end if;
                when "01001100" =>
                  \$v5420\ := \$ram_lock\;
                  if \$v5420\(0) = '1' then
                    state_var5920 := Q_WAIT5419;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18788\(48 to 63), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5418;
                  end if;
                when "01001111" =>
                  \$v5423\ := \$ram_lock\;
                  if \$v5423\(0) = '1' then
                    state_var5920 := Q_WAIT5422;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18788\(16 to 46),16)));
                    state_var5920 := PAUSE_GET5421;
                  end if;
                when "01010000" =>
                  \$v5429\ := \$ram_lock\;
                  if \$v5429\(0) = '1' then
                    state_var5920 := Q_WAIT5428;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18788\(48 to 63), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5427;
                  end if;
                when "01010001" =>
                  \$v5438\ := \$ram_lock\;
                  if \$v5438\(0) = '1' then
                    state_var5920 := Q_WAIT5437;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18788\(48 to 63), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5436;
                  end if;
                when "01010010" =>
                  \$v5444\ := \$ram_lock\;
                  if \$v5444\(0) = '1' then
                    state_var5920 := Q_WAIT5443;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18788\(48 to 63), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5442;
                  end if;
                when "01010011" =>
                  \$v5453\ := \$ram_lock\;
                  if \$v5453\(0) = '1' then
                    state_var5920 := Q_WAIT5452;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18788\(48 to 63), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5451;
                  end if;
                when "01010101" =>
                  \$18797_branch_if648_id\ := "000001000001";
                  \$18797_branch_if648_arg\ := eclat_false & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  state_var5920 := \$18797_BRANCH_IF648\;
                when "01010110" =>
                  \$18797_branch_if648_id\ := "000001000010";
                  \$18797_branch_if648_arg\ := eclat_true & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  state_var5920 := \$18797_BRANCH_IF648\;
                when "01011000" =>
                  result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & 
                  eclat_if(work.Int.eq(\$18788\(16 to 46), "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when "01011010" =>
                  \$v5456\ := \$ram_lock\;
                  if \$v5456\(0) = '1' then
                    state_var5920 := Q_WAIT5455;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                   \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5454;
                  end if;
                when "01011011" =>
                  \$v5468\ := \$ram_lock\;
                  if \$v5468\(0) = '1' then
                    state_var5920 := Q_WAIT5467;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18788\(104 to 119), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5466;
                  end if;
                when "01100011" =>
                  result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & "000"& X"000000" & X"0" & eclat_true & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when "01100100" =>
                  result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when "01100101" =>
                  result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & "000"& X"000000" & X"2" & eclat_true & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when "01100110" =>
                  result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & "000"& X"000000" & X"3" & eclat_true & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when "01101000" =>
                  \$v5471\ := \$ram_lock\;
                  if \$v5471\(0) = '1' then
                    state_var5920 := Q_WAIT5470;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5469;
                  end if;
                when "01101001" =>
                  \$v5474\ := \$ram_lock\;
                  if \$v5474\(0) = '1' then
                    state_var5920 := Q_WAIT5473;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5472;
                  end if;
                when "01101010" =>
                  \$v5477\ := \$ram_lock\;
                  if \$v5477\(0) = '1' then
                    state_var5920 := Q_WAIT5476;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5475;
                  end if;
                when "01101011" =>
                  \$v5480\ := \$ram_lock\;
                  if \$v5480\(0) = '1' then
                    state_var5920 := Q_WAIT5479;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                    \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5478;
                  end if;
                when "01101110" =>
                  \$18901_binop_int6434361_id\ := "000001000111";
                  \$18901_binop_int6434361_arg\ := X"0000000" & X"0" & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  state_var5920 := \$18901_BINOP_INT6434361\;
                when "01101111" =>
                  \$18920_binop_int6434362_id\ := "000001001100";
                  \$18920_binop_int6434362_arg\ := X"0000000" & X"1" & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  state_var5920 := \$18920_BINOP_INT6434362\;
                when "01110000" =>
                  \$18939_binop_int6434363_id\ := "000001010001";
                  \$18939_binop_int6434363_arg\ := X"0000000" & X"2" & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  state_var5920 := \$18939_BINOP_INT6434363\;
                when "01110001" =>
                  \$18958_binop_int6434364_id\ := "000001010110";
                  \$18958_binop_int6434364_arg\ := X"0000000" & X"3" & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  state_var5920 := \$18958_BINOP_INT6434364\;
                when "01110010" =>
                  \$18977_binop_int6434365_id\ := "000001011011";
                  \$18977_binop_int6434365_arg\ := X"0000000" & X"4" & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  state_var5920 := \$18977_BINOP_INT6434365\;
                when "01110011" =>
                  \$18996_binop_int6434366_id\ := "000001100000";
                  \$18996_binop_int6434366_arg\ := X"0000000" & X"5" & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  state_var5920 := \$18996_BINOP_INT6434366\;
                when "01110100" =>
                  \$19015_binop_int6434367_id\ := "000001100101";
                  \$19015_binop_int6434367_arg\ := X"0000000" & X"6" & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  state_var5920 := \$19015_BINOP_INT6434367\;
                when "01110101" =>
                  \$19034_binop_int6434368_id\ := "000001101010";
                  \$19034_binop_int6434368_arg\ := X"0000000" & X"7" & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  state_var5920 := \$19034_BINOP_INT6434368\;
                when "01110110" =>
                  \$19053_binop_int6434369_id\ := "000001101111";
                  \$19053_binop_int6434369_arg\ := X"0000000" & X"8" & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  state_var5920 := \$19053_BINOP_INT6434369\;
                when "01110111" =>
                  \$19072_binop_int6434370_id\ := "000001110100";
                  \$19072_binop_int6434370_arg\ := X"0000000" & X"9" & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  state_var5920 := \$19072_BINOP_INT6434370\;
                when "01111000" =>
                  \$19091_binop_int6434371_id\ := "000001111001";
                  \$19091_binop_int6434371_arg\ := X"0000000" & X"a" & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  state_var5920 := \$19091_BINOP_INT6434371\;
                when "10000010" =>
                  \$19110\ := work.Print.print_string(clk,of_string("fatal error: "));
                  \$19111\ := work.Print.print_string(clk,of_string("unsupported instruction GETMETHOD"));
                  \$19112\ := work.Print.print_newline(clk,eclat_unit);
                  \$19113_forever6704372_id\ := "000001111010";
                  \$19113_forever6704372_arg\ := eclat_unit;
                  state_var5920 := \$19113_FOREVER6704372\;
                when "10001001" =>
                  \$19116_binop_int6434373_id\ := "000001111111";
                  \$19116_binop_int6434373_arg\ := X"0000000" & X"b" & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  state_var5920 := \$19116_BINOP_INT6434373\;
                when "10001010" =>
                  \$19135_binop_int6434374_id\ := "000010000100";
                  \$19135_binop_int6434374_arg\ := X"0000000" & X"c" & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  state_var5920 := \$19135_BINOP_INT6434374\;
                when "10001101" =>
                  \$19154\ := work.Print.print_string(clk,of_string("fatal error: "));
                  \$19155\ := work.Print.print_string(clk,of_string("unsupported instruction GETPUBMET"));
                  \$19156\ := work.Print.print_newline(clk,eclat_unit);
                  \$19157_forever6704375_id\ := "000010000101";
                  \$19157_forever6704375_arg\ := eclat_unit;
                  state_var5920 := \$19157_FOREVER6704375\;
                when "10001110" =>
                  \$19160\ := work.Print.print_string(clk,of_string("fatal error: "));
                  \$19161\ := work.Print.print_string(clk,of_string("unsupported instruction GETDYNMET"));
                  \$19162\ := work.Print.print_newline(clk,eclat_unit);
                  \$19163_forever6704376_id\ := "000010000110";
                  \$19163_forever6704376_arg\ := eclat_unit;
                  state_var5920 := \$19163_FOREVER6704376\;
                when "01111001" =>
                  \$19166_binop_compare6454377_id\ := "000010001000";
                  \$19166_binop_compare6454377_arg\ := X"0000000" & X"0" & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  state_var5920 := \$19166_BINOP_COMPARE6454377\;
                when "01111010" =>
                  \$19174_binop_compare6454378_id\ := "000010001010";
                  \$19174_binop_compare6454378_arg\ := X"0000000" & X"1" & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  state_var5920 := \$19174_BINOP_COMPARE6454378\;
                when "01111011" =>
                  \$19182_binop_compare6454379_id\ := "000010001100";
                  \$19182_binop_compare6454379_arg\ := X"0000000" & X"2" & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  state_var5920 := \$19182_BINOP_COMPARE6454379\;
                when "01111100" =>
                  \$19190_binop_compare6454380_id\ := "000010001110";
                  \$19190_binop_compare6454380_arg\ := X"0000000" & X"3" & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  state_var5920 := \$19190_BINOP_COMPARE6454380\;
                when "01111101" =>
                  \$19198_binop_compare6454381_id\ := "000010010000";
                  \$19198_binop_compare6454381_arg\ := X"0000000" & X"4" & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  state_var5920 := \$19198_BINOP_COMPARE6454381\;
                when "01111110" =>
                  \$19206_binop_compare6454382_id\ := "000010010010";
                  \$19206_binop_compare6454382_arg\ := X"0000000" & X"5" & \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  state_var5920 := \$19206_BINOP_COMPARE6454382\;
                when "10000001" =>
                  result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & 
                  eclat_if(""&\$18788\(47) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when "10001111" =>
                  \$19214\ := work.Print.print_string(clk,of_string("STOP : "));
                  result4928 := \$18788\(0 to 15) & \$18788\(16 to 47) & \$18788\(48 to 63) & \$18788\(64 to 119) & eclat_true & ""&\$18788\(121);
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                when others =>
                  \$v5909\ := \$code_lock\;
                  if \$v5909\(0) = '1' then
                    state_var5920 := Q_WAIT5908;
                  else
                    acquire(\$code_lock\);
                    \$code_ptr\ <= to_integer(unsigned(work.Int.add(\$18788\(0 to 15), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5907;
                  end if;
                end case;
              when PAUSE_SET4931 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19762\ := eclat_unit;
                \$18790_loop666_arg\ := work.Int.add(\$18790_loop666_arg\(0 to 15), X"000" & X"1") & \$18790_loop666_arg\(16 to 31) & \$18790_loop666_arg\(32 to 47) & \$18790_loop666_arg\(48 to 63);
                state_var5920 := \$18790_LOOP666\;
              when PAUSE_SET4938 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19743\ := eclat_unit;
                \$18791_loop665_arg\ := work.Int.add(\$18791_loop665_arg\(0 to 15), X"000" & X"1") & \$19742\(32 to 47) & \$18791_loop665_arg\(32 to 47) & \$18791_loop665_arg\(48 to 63) & \$18791_loop665_arg\(64 to 79) & \$18791_loop665_arg\(80 to 95);
                state_var5920 := \$18791_LOOP665\;
              when PAUSE_SET4941 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19758\ := eclat_unit;
                \$19742\ := eclat_resize(\$18791_loop665_arg\(16 to 31),31) & eclat_false & 
                work.Int.add(\$18791_loop665_arg\(16 to 31), work.Int.add(
                                                             eclat_resize(
                                                             work.Int.lsr(
                                                             \$19745_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$v4940\ := \$ram_lock\;
                if \$v4940\(0) = '1' then
                  state_var5920 := Q_WAIT4939;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$18791_loop665_arg\(64 to 79), \$18791_loop665_arg\(0 to 15))));
                  \$ram_write\ <= \$19742\(0 to 31); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET4938;
                end if;
              when PAUSE_SET4944 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19757\ := eclat_unit;
                \$v4943\ := \$ram_lock\;
                if \$v4943\(0) = '1' then
                  state_var5920 := Q_WAIT4942;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$19741\(0 to 30),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$18791_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET4941;
                end if;
              when PAUSE_SET4947 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19755\ := eclat_unit;
                \$18790_loop666_id\ := "000000100000";
                \$18790_loop666_arg\ := X"000" & X"1" & \$18791_loop665_arg\(16 to 31) & eclat_resize(\$19741\(0 to 30),16) & eclat_resize(
                work.Int.lsr(\$19745_hd\(0 to 30), X"0000000" & X"2"),16);
                state_var5920 := \$18790_LOOP666\;
              when PAUSE_SET5172 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19489\ := eclat_unit;
                \$18793_make_block579_result\ := \$19485\(0 to 31) & \$19485\(32 to 63) & eclat_resize(\$19485\(64 to 79),31) & eclat_false;
                case \$18793_make_block579_id\ is
                when "000000110100" =>
                  \$19444\ := \$18793_make_block579_result\;
                  \$v5230\ := ""&\$18796_make_block_n646_arg\(32);
                  if \$v5230\(0) = '1' then
                    \$v5229\ := \$ram_lock\;
                    if \$v5229\(0) = '1' then
                      state_var5920 := Q_WAIT5228;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                              work.Int.add(
                                                              eclat_resize(\$19444\(64 to 94),16), X"000" & X"0"), X"000" & X"1")));
                      \$ram_write\ <= \$19444\(0 to 31); \$ram_write_request\ <= '1';
                      state_var5920 := PAUSE_SET5227;
                    end if;
                  else
                    \$19445\ := eclat_unit;
                    \$v5226\ := ""&\$18796_make_block_n646_arg\(33);
                    if \$v5226\(0) = '1' then
                      \$v5225\ := \$ram_lock\;
                      if \$v5225\(0) = '1' then
                        state_var5920 := Q_WAIT5224;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(
                                                          \$18796_make_block_n646_arg\(16 to 31), X"000" & X"1")));
                        state_var5920 := PAUSE_GET5223;
                      end if;
                    else
                      \$19446_sp\ := \$18796_make_block_n646_arg\(16 to 31);
                      \$v5219\ := ""&\$18796_make_block_n646_arg\(34);
                      if \$v5219\(0) = '1' then
                        \$v5218\ := \$ram_lock\;
                        if \$v5218\(0) = '1' then
                          state_var5920 := Q_WAIT5217;
                        else
                          acquire(\$ram_lock\);
                          \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(
                                                            \$19446_sp\, X"000" & X"1")));
                          state_var5920 := PAUSE_GET5216;
                        end if;
                      else
                        \$19447_sp\ := \$19446_sp\;
                        \$18796_make_block_n646_result\ := \$18796_make_block_n646_arg\(0 to 15) & \$19444\(64 to 95) & \$19447_sp\ & \$19444\(32 to 63) & \$18796_make_block_n646_arg\(148 to 155) & \$18796_make_block_n646_arg\(156 to 171) & \$18796_make_block_n646_arg\(114 to 115);
                        result4928 := \$18796_make_block_n646_result\;
                        rdy4929 := eclat_true;
                        state_var5920 := IDLE4930;
                      end if;
                    end if;
                  end if;
                when "000010010111" =>
                  \$19231\ := \$18793_make_block579_result\;
                  \$v5702\ := \$ram_lock\;
                  if \$v5702\(0) = '1' then
                    state_var5920 := Q_WAIT5701;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            work.Int.add(
                                                            eclat_resize(\$19231\(64 to 94),16), X"000" & X"0"), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(work.Int.sub(work.Int.add(
                                                              \$18788\(0 to 15), X"000" & X"2"), X"000" & X"3"),31) & eclat_true; \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5700;
                  end if;
                when "000010101000" =>
                  \$19344\ := \$18793_make_block579_result\;
                  \$v5838\ := \$ram_lock\;
                  if \$v5838\(0) = '1' then
                    state_var5920 := Q_WAIT5837;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            work.Int.add(
                                                            eclat_resize(\$19344\(64 to 94),16), X"000" & X"0"), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(work.Int.add(work.Int.add(
                                                              \$18788\(0 to 15), X"000" & X"2"), eclat_resize(\$19340_argument2\,16)),31) & eclat_true; \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5836;
                  end if;
                when "000010101010" =>
                  \$19358\ := \$18793_make_block579_result\;
                  \$v5867\ := \$ram_lock\;
                  if \$v5867\(0) = '1' then
                    state_var5920 := Q_WAIT5866;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            work.Int.add(
                                                            eclat_resize(\$19358\(64 to 94),16), X"000" & X"0"), X"000" & X"1")));
                    \$ram_write\ <= \$19358\(0 to 31); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5865;
                  end if;
                when "000010111010" =>
                  \$19410\ := \$18793_make_block579_result\;
                  \$v5890\ := \$ram_lock\;
                  if \$v5890\(0) = '1' then
                    state_var5920 := Q_WAIT5889;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            work.Int.add(
                                                            eclat_resize(\$19410\(64 to 94),16), X"000" & X"0"), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(work.Int.add(work.Int.add(
                                                              \$18788\(0 to 15), X"000" & X"3"), eclat_resize(\$19408_argument3\,16)),31) & eclat_true; \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5888;
                  end if;
                when others =>
                  
                end case;
              when PAUSE_SET5178 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19470\ := eclat_unit;
                \$19468_sp\ := work.Int.add(\$19467_sp\, X"000" & X"1");
                \$v5177\ := \$ram_lock\;
                if \$v5177\(0) = '1' then
                  state_var5920 := Q_WAIT5176;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18794_apply638_arg\(60 to 90),16), X"000" & X"0"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5175;
                end if;
              when PAUSE_SET5182 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19471\ := eclat_unit;
                \$19467_sp\ := work.Int.add(\$19466_sp\, X"000" & X"1");
                \$v5181\ := ""&\$18794_apply638_arg\(0);
                if \$v5181\(0) = '1' then
                  \$v5180\ := \$ram_lock\;
                  if \$v5180\(0) = '1' then
                    state_var5920 := Q_WAIT5179;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19467_sp\));
                    \$ram_write\ <= \$19462\(0 to 31); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5178;
                  end if;
                else
                  \$19468_sp\ := \$19467_sp\;
                  \$v5177\ := \$ram_lock\;
                  if \$v5177\(0) = '1' then
                    state_var5920 := Q_WAIT5176;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$18794_apply638_arg\(60 to 90),16), X"000" & X"0"), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5175;
                  end if;
                end if;
              when PAUSE_SET5186 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19472\ := eclat_unit;
                \$19466_sp\ := work.Int.add(\$19465_sp\, X"000" & X"1");
                \$v5185\ := ""&\$18794_apply638_arg\(1);
                if \$v5185\(0) = '1' then
                  \$v5184\ := \$ram_lock\;
                  if \$v5184\(0) = '1' then
                    state_var5920 := Q_WAIT5183;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19466_sp\));
                    \$ram_write\ <= \$19463\(0 to 31); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5182;
                  end if;
                else
                  \$19467_sp\ := \$19466_sp\;
                  \$v5181\ := ""&\$18794_apply638_arg\(0);
                  if \$v5181\(0) = '1' then
                    \$v5180\ := \$ram_lock\;
                    if \$v5180\(0) = '1' then
                      state_var5920 := Q_WAIT5179;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(\$19467_sp\));
                      \$ram_write\ <= \$19462\(0 to 31); \$ram_write_request\ <= '1';
                      state_var5920 := PAUSE_SET5178;
                    end if;
                  else
                    \$19468_sp\ := \$19467_sp\;
                    \$v5177\ := \$ram_lock\;
                    if \$v5177\(0) = '1' then
                      state_var5920 := Q_WAIT5176;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                        work.Int.add(
                                                        eclat_resize(\$18794_apply638_arg\(60 to 90),16), X"000" & X"0"), X"000" & X"1")));
                      state_var5920 := PAUSE_GET5175;
                    end if;
                  end if;
                end if;
              when PAUSE_SET5190 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19475\ := eclat_unit;
                \$19465_sp\ := work.Int.add(work.Int.add(work.Int.add(
                                                         \$19464\(32 to 47), X"000" & X"1"), X"000" & X"1"), X"000" & X"1");
                \$v5189\ := ""&\$18794_apply638_arg\(2);
                if \$v5189\(0) = '1' then
                  \$v5188\ := \$ram_lock\;
                  if \$v5188\(0) = '1' then
                    state_var5920 := Q_WAIT5187;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$19465_sp\));
                    \$ram_write\ <= \$19464\(0 to 31); \$ram_write_request\ <= '1';
                    state_var5920 := PAUSE_SET5186;
                  end if;
                else
                  \$19466_sp\ := \$19465_sp\;
                  \$v5185\ := ""&\$18794_apply638_arg\(1);
                  if \$v5185\(0) = '1' then
                    \$v5184\ := \$ram_lock\;
                    if \$v5184\(0) = '1' then
                      state_var5920 := Q_WAIT5183;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(\$19466_sp\));
                      \$ram_write\ <= \$19463\(0 to 31); \$ram_write_request\ <= '1';
                      state_var5920 := PAUSE_SET5182;
                    end if;
                  else
                    \$19467_sp\ := \$19466_sp\;
                    \$v5181\ := ""&\$18794_apply638_arg\(0);
                    if \$v5181\(0) = '1' then
                      \$v5180\ := \$ram_lock\;
                      if \$v5180\(0) = '1' then
                        state_var5920 := Q_WAIT5179;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr_write\ <= to_integer(unsigned(\$19467_sp\));
                        \$ram_write\ <= \$19462\(0 to 31); \$ram_write_request\ <= '1';
                        state_var5920 := PAUSE_SET5178;
                      end if;
                    else
                      \$19468_sp\ := \$19467_sp\;
                      \$v5177\ := \$ram_lock\;
                      if \$v5177\(0) = '1' then
                        state_var5920 := Q_WAIT5176;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$18794_apply638_arg\(60 to 90),16), X"000" & X"0"), X"000" & X"1")));
                        state_var5920 := PAUSE_GET5175;
                      end if;
                    end if;
                  end if;
                end if;
              when PAUSE_SET5193 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19474\ := eclat_unit;
                \$v5192\ := \$ram_lock\;
                if \$v5192\(0) = '1' then
                  state_var5920 := Q_WAIT5191;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          \$19464\(32 to 47), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(work.Int.add(\$18794_apply638_arg\(44 to 59), X"000" & X"1"),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5190;
                end if;
              when PAUSE_SET5196 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19473\ := eclat_unit;
                \$v5195\ := \$ram_lock\;
                if \$v5195\(0) = '1' then
                  state_var5920 := Q_WAIT5194;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$19464\(32 to 47), X"000" & X"1")));
                  \$ram_write\ <= \$18794_apply638_arg\(110 to 141); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5193;
                end if;
              when PAUSE_SET5213 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19449\ := eclat_unit;
                \$19447_sp\ := work.Int.sub(\$19446_sp\, X"000" & X"1");
                \$18796_make_block_n646_result\ := \$18796_make_block_n646_arg\(0 to 15) & \$19444\(64 to 95) & \$19447_sp\ & \$19444\(32 to 63) & \$18796_make_block_n646_arg\(148 to 155) & \$18796_make_block_n646_arg\(156 to 171) & \$18796_make_block_n646_arg\(114 to 115);
                result4928 := \$18796_make_block_n646_result\;
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_SET5220 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19451\ := eclat_unit;
                \$19446_sp\ := work.Int.sub(\$18796_make_block_n646_arg\(16 to 31), X"000" & X"1");
                \$v5219\ := ""&\$18796_make_block_n646_arg\(34);
                if \$v5219\(0) = '1' then
                  \$v5218\ := \$ram_lock\;
                  if \$v5218\(0) = '1' then
                    state_var5920 := Q_WAIT5217;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19446_sp\, X"000" & X"1")));
                    state_var5920 := PAUSE_GET5216;
                  end if;
                else
                  \$19447_sp\ := \$19446_sp\;
                  \$18796_make_block_n646_result\ := \$18796_make_block_n646_arg\(0 to 15) & \$19444\(64 to 95) & \$19447_sp\ & \$19444\(32 to 63) & \$18796_make_block_n646_arg\(148 to 155) & \$18796_make_block_n646_arg\(156 to 171) & \$18796_make_block_n646_arg\(114 to 115);
                  result4928 := \$18796_make_block_n646_result\;
                  rdy4929 := eclat_true;
                  state_var5920 := IDLE4930;
                end if;
              when PAUSE_SET5227 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19445\ := eclat_unit;
                \$v5226\ := ""&\$18796_make_block_n646_arg\(33);
                if \$v5226\(0) = '1' then
                  \$v5225\ := \$ram_lock\;
                  if \$v5225\(0) = '1' then
                    state_var5920 := Q_WAIT5224;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18796_make_block_n646_arg\(16 to 31), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5223;
                  end if;
                else
                  \$19446_sp\ := \$18796_make_block_n646_arg\(16 to 31);
                  \$v5219\ := ""&\$18796_make_block_n646_arg\(34);
                  if \$v5219\(0) = '1' then
                    \$v5218\ := \$ram_lock\;
                    if \$v5218\(0) = '1' then
                      state_var5920 := Q_WAIT5217;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(
                                                        \$19446_sp\, X"000" & X"1")));
                      state_var5920 := PAUSE_GET5216;
                    end if;
                  else
                    \$19447_sp\ := \$19446_sp\;
                    \$18796_make_block_n646_result\ := \$18796_make_block_n646_arg\(0 to 15) & \$19444\(64 to 95) & \$19447_sp\ & \$19444\(32 to 63) & \$18796_make_block_n646_arg\(148 to 155) & \$18796_make_block_n646_arg\(156 to 171) & \$18796_make_block_n646_arg\(114 to 115);
                    result4928 := \$18796_make_block_n646_result\;
                    rdy4929 := eclat_true;
                    state_var5920 := IDLE4930;
                  end if;
                end if;
              when PAUSE_SET5235 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19438\ := eclat_unit;
                \$18798_w652_arg\ := work.Int.add(\$18798_w652_arg\(0 to 15), X"000" & X"1") & \$18798_w652_arg\(16 to 31) & \$18798_w652_arg\(32 to 47) & \$18798_w652_arg\(48 to 63);
                state_var5920 := \$18798_W652\;
              when PAUSE_SET5242 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19434\ := eclat_unit;
                \$18799_w1656_arg\ := work.Int.add(\$18799_w1656_arg\(0 to 15), X"000" & X"1") & \$18799_w1656_arg\(16 to 31) & \$18799_w1656_arg\(32 to 47) & \$18799_w1656_arg\(48 to 79);
                state_var5920 := \$18799_W1656\;
              when PAUSE_SET5248 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19432\ := eclat_unit;
                \$v5247\ := \$code_lock\;
                if \$v5247\(0) = '1' then
                  state_var5920 := Q_WAIT5246;
                else
                  acquire(\$code_lock\);
                  \$code_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                  \$18799_w1656_arg\(16 to 31), X"000" & X"3"), \$18799_w1656_arg\(0 to 15))));
                  state_var5920 := PAUSE_GET5245;
                end if;
              when PAUSE_SET5276 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18825\ := eclat_unit;
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18788\(16 to 47) & 
                work.Int.add(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_SET5279 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18826\ := eclat_unit;
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & \$18788\(16 to 47) & 
                work.Int.add(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_SET5285 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18827\ := eclat_unit;
                \$v5284\ := \$ram_lock\;
                if \$v5284\(0) = '1' then
                  state_var5920 := Q_WAIT5283;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5282;
                end if;
              when PAUSE_SET5291 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18829\ := eclat_unit;
                \$v5290\ := \$ram_lock\;
                if \$v5290\(0) = '1' then
                  state_var5920 := Q_WAIT5289;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"2"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5288;
                end if;
              when PAUSE_SET5297 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18831\ := eclat_unit;
                \$v5296\ := \$ram_lock\;
                if \$v5296\(0) = '1' then
                  state_var5920 := Q_WAIT5295;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"3"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5294;
                end if;
              when PAUSE_SET5303 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18833\ := eclat_unit;
                \$v5302\ := \$ram_lock\;
                if \$v5302\(0) = '1' then
                  state_var5920 := Q_WAIT5301;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"4"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5300;
                end if;
              when PAUSE_SET5309 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18835\ := eclat_unit;
                \$v5308\ := \$ram_lock\;
                if \$v5308\(0) = '1' then
                  state_var5920 := Q_WAIT5307;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"5"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5306;
                end if;
              when PAUSE_SET5315 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18837\ := eclat_unit;
                \$v5314\ := \$ram_lock\;
                if \$v5314\(0) = '1' then
                  state_var5920 := Q_WAIT5313;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"6"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5312;
                end if;
              when PAUSE_SET5321 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18839\ := eclat_unit;
                \$v5320\ := \$ram_lock\;
                if \$v5320\(0) = '1' then
                  state_var5920 := Q_WAIT5319;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"7"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5318;
                end if;
              when PAUSE_SET5339 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18845\ := eclat_unit;
                \$v5338\ := \$ram_lock\;
                if \$v5338\(0) = '1' then
                  state_var5920 := Q_WAIT5337;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18788\(64 to 94),16), 
                                                                 work.Int.sub(
                                                                 X"000" & X"1", X"000" & X"1")), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5336;
                end if;
              when PAUSE_SET5345 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18847\ := eclat_unit;
                \$v5344\ := \$ram_lock\;
                if \$v5344\(0) = '1' then
                  state_var5920 := Q_WAIT5343;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18788\(64 to 94),16), 
                                                                 work.Int.sub(
                                                                 X"000" & X"2", X"000" & X"1")), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5342;
                end if;
              when PAUSE_SET5351 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18849\ := eclat_unit;
                \$v5350\ := \$ram_lock\;
                if \$v5350\(0) = '1' then
                  state_var5920 := Q_WAIT5349;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18788\(64 to 94),16), 
                                                                 work.Int.sub(
                                                                 X"000" & X"3", X"000" & X"1")), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5348;
                end if;
              when PAUSE_SET5357 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18851\ := eclat_unit;
                \$v5356\ := \$ram_lock\;
                if \$v5356\(0) = '1' then
                  state_var5920 := Q_WAIT5355;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18788\(64 to 94),16), 
                                                                 work.Int.sub(
                                                                 X"000" & X"4", X"000" & X"1")), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5354;
                end if;
              when PAUSE_SET5363 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18860\ := eclat_unit;
                \$18856_loop_push6494360_arg\ := work.Int.add(\$18856_loop_push6494360_arg\(0 to 15), X"000" & X"1") & 
                work.Int.add(\$18856_loop_push6494360_arg\(16 to 23), "00000001") & \$18856_loop_push6494360_arg\(24 to 55) & \$18856_loop_push6494360_arg\(56 to 63);
                state_var5920 := \$18856_LOOP_PUSH6494360\;
              when PAUSE_SET5373 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18861\ := eclat_unit;
                \$18795_offsetclosure_n639_id\ := "000000111100";
                \$18795_offsetclosure_n639_arg\ := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & 
                work.Int.add(\$18788\(48 to 63), X"000" & X"1") & work.Int.neg(
                                                                  X"000" & X"2") & \$18788\(64 to 119) & \$18788\(120 to 121) & \$18788\(64 to 95);
                state_var5920 := \$18795_OFFSETCLOSURE_N639\;
              when PAUSE_SET5376 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18862\ := eclat_unit;
                \$18795_offsetclosure_n639_id\ := "000000111101";
                \$18795_offsetclosure_n639_arg\ := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & 
                work.Int.add(\$18788\(48 to 63), X"000" & X"1") & X"000" & X"0" & \$18788\(64 to 119) & \$18788\(120 to 121) & \$18788\(64 to 95);
                state_var5920 := \$18795_OFFSETCLOSURE_N639\;
              when PAUSE_SET5379 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18863\ := eclat_unit;
                \$18795_offsetclosure_n639_id\ := "000000111110";
                \$18795_offsetclosure_n639_arg\ := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & 
                work.Int.add(\$18788\(48 to 63), X"000" & X"1") & X"000" & X"2" & \$18788\(64 to 119) & \$18788\(120 to 121) & \$18788\(64 to 95);
                state_var5920 := \$18795_OFFSETCLOSURE_N639\;
              when PAUSE_SET5382 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18864\ := eclat_unit;
                \$18796_make_block_n646_id\ := "000001000000";
                \$18796_make_block_n646_arg\ := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & 
                work.Int.add(\$18788\(48 to 63), X"000" & X"1") & eclat_false & eclat_false & eclat_false & "000"& X"000000" & X"0" & X"000" & X"0" & \$18788\(16 to 47) & \$18788\(120 to 121) & \$18788\(64 to 95) & \$18788\(96 to 103) & \$18788\(104 to 119);
                state_var5920 := \$18796_MAKE_BLOCK_N646\;
              when PAUSE_SET5397 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18874\ := eclat_unit;
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & 
                work.Int.sub(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_SET5403 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18876\ := eclat_unit;
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & 
                work.Int.sub(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_SET5409 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18878\ := eclat_unit;
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & 
                work.Int.sub(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_SET5415 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18880\ := eclat_unit;
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & 
                work.Int.sub(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_SET5430 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18886\ := eclat_unit;
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & 
                work.Int.sub(work.Int.sub(\$18788\(48 to 63), X"000" & X"1"), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_SET5445 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18891\ := eclat_unit;
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & 
                work.Int.sub(work.Int.sub(\$18788\(48 to 63), X"000" & X"1"), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_SET5469 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18897\ := eclat_unit;
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & "000"& X"000000" & X"0" & eclat_true & 
                work.Int.add(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_SET5472 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18898\ := eclat_unit;
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & 
                work.Int.add(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_SET5475 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18899\ := eclat_unit;
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & "000"& X"000000" & X"2" & eclat_true & 
                work.Int.add(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_SET5478 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18900\ := eclat_unit;
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"1") & "000"& X"000000" & X"3" & eclat_true & 
                work.Int.add(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_SET5641 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19217\ := eclat_unit;
                \$v5640\ := \$ram_lock\;
                if \$v5640\(0) = '1' then
                  state_var5920 := Q_WAIT5639;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$18788\(48 to 63), X"000" & X"1"), eclat_resize(\$19215_argument1\,16)), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5638;
                end if;
              when PAUSE_SET5644 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19219\ := eclat_unit;
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"2") & "000"& X"000000" & X"1" & eclat_true & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_SET5653 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19221\ := eclat_unit;
                \$v5652\ := \$ram_lock\;
                if \$v5652\(0) = '1' then
                  state_var5920 := Q_WAIT5651;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18788\(64 to 94),16), 
                                                                 work.Int.sub(
                                                                 eclat_resize(\$19215_argument1\,16), X"000" & X"1")), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5650;
                end if;
              when PAUSE_SET5656 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19225\ := eclat_unit;
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"2") & \$18788\(16 to 47) & 
                work.Int.add(work.Int.add(work.Int.add(\$18788\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_SET5659 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19224\ := eclat_unit;
                \$v5658\ := \$ram_lock\;
                if \$v5658\(0) = '1' then
                  state_var5920 := Q_WAIT5657;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(work.Int.add(work.Int.add(
                                                            \$18788\(0 to 15), X"000" & X"1"), eclat_resize(\$19215_argument1\,16)),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5656;
                end if;
              when PAUSE_SET5662 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19223\ := eclat_unit;
                \$v5661\ := \$ram_lock\;
                if \$v5661\(0) = '1' then
                  state_var5920 := Q_WAIT5660;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$18788\(48 to 63), X"000" & X"1")));
                  \$ram_write\ <= \$18788\(64 to 95); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5659;
                end if;
              when PAUSE_SET5690 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19242\ := eclat_unit;
                \$19238_w6514383_arg\ := work.Int.add(\$19238_w6514383_arg\(0 to 7), "00000001") & 
                work.Int.sub(\$19238_w6514383_arg\(8 to 23), X"000" & X"1") & \$19238_w6514383_arg\(24 to 31) & \$19238_w6514383_arg\(32 to 63);
                state_var5920 := \$19238_W6514383\;
              when PAUSE_SET5697 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19233\ := eclat_unit;
                \$19238_w6514383_id\ := "000010010110";
                \$19238_w6514383_arg\ := "00000000" & \$18788\(48 to 63) & \$18788\(96 to 103) & \$19231\(64 to 95);
                state_var5920 := \$19238_W6514383\;
              when PAUSE_SET5700 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19232\ := eclat_unit;
                \$v5699\ := \$ram_lock\;
                if \$v5699\(0) = '1' then
                  state_var5920 := Q_WAIT5698;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$19231\(64 to 94),16), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= \$19231\(32 to 63); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5697;
                end if;
              when PAUSE_SET5704 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19243\ := eclat_unit;
                \$18795_offsetclosure_n639_id\ := "000010011001";
                \$18795_offsetclosure_n639_arg\ := work.Int.add(\$18788\(0 to 15), X"000" & X"2") & 
                work.Int.add(\$18788\(48 to 63), X"000" & X"1") & eclat_resize(\$19215_argument1\,16) & \$18788\(64 to 119) & \$18788\(120 to 121) & \$18788\(64 to 95);
                state_var5920 := \$18795_OFFSETCLOSURE_N639\;
              when PAUSE_SET5713 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19245\ := eclat_unit;
                \$v5712\ := \$ram_lock\;
                if \$v5712\(0) = '1' then
                  state_var5920 := Q_WAIT5711;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(X"3e80", eclat_resize(\$19215_argument1\,16))));
                  state_var5920 := PAUSE_GET5710;
                end if;
              when PAUSE_SET5716 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19247\ := eclat_unit;
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"2") & "000"& X"000000" & X"1" & eclat_true & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_SET5719 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19248\ := eclat_unit;
                \$18796_make_block_n646_id\ := "000010011011";
                \$18796_make_block_n646_arg\ := work.Int.add(\$18788\(0 to 15), X"000" & X"2") & 
                work.Int.add(\$18788\(48 to 63), X"000" & X"1") & eclat_false & eclat_false & eclat_false & \$19215_argument1\ & X"000" & X"0" & \$18788\(16 to 47) & \$18788\(120 to 121) & \$18788\(64 to 95) & \$18788\(96 to 103) & \$18788\(104 to 119);
                state_var5920 := \$18796_MAKE_BLOCK_N646\;
              when PAUSE_SET5725 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19258\ := eclat_unit;
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"2") & "000"& X"000000" & X"1" & eclat_true & 
                work.Int.sub(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_SET5738 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19271\ := eclat_unit;
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"2") & \$18788\(16 to 47) & 
                work.Int.add(work.Int.add(work.Int.add(work.Int.add(\$18788\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1"), X"000" & X"1") & \$18788\(64 to 95) & \$18788\(96 to 103) & 
                work.Int.add(work.Int.add(work.Int.add(work.Int.add(\$18788\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1"), X"000" & X"1") & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_SET5741 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19270\ := eclat_unit;
                \$v5740\ := \$ram_lock\;
                if \$v5740\(0) = '1' then
                  state_var5920 := Q_WAIT5739;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          work.Int.add(
                                                          \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(work.Int.add(work.Int.add(
                                                            \$18788\(0 to 15), X"000" & X"1"), eclat_resize(\$19215_argument1\,16)),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5738;
                end if;
              when PAUSE_SET5744 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19269\ := eclat_unit;
                \$v5743\ := \$ram_lock\;
                if \$v5743\(0) = '1' then
                  state_var5920 := Q_WAIT5742;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$18788\(104 to 119),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5741;
                end if;
              when PAUSE_SET5747 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19268\ := eclat_unit;
                \$v5746\ := \$ram_lock\;
                if \$v5746\(0) = '1' then
                  state_var5920 := Q_WAIT5745;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$18788\(48 to 63), X"000" & X"1")));
                  \$ram_write\ <= \$18788\(64 to 95); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5744;
                end if;
              when PAUSE_SET5754 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19272\ := eclat_unit;
                \$v5753\ := \$19215_argument1\;
                case \$v5753\ is
                when "000"& X"000000" & X"0" =>
                  \$19275\ := work.Print.print_string(clk,of_string("======> "));
                  \$19276\ := work.Int.print(clk,\$18788\(16 to 46));
                  \$19277\ := work.Print.print_newline(clk,eclat_unit);
                  \$19273\ := "000"& X"000000" & X"1" & eclat_true & \$18788\(0 to 15) & \$18788\(16 to 47) & 
                  work.Int.add(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 95) & \$18788\(96 to 103) & \$18788\(104 to 119) & \$18788\(120 to 121);
                  \$v5752\ := \$ram_lock\;
                  if \$v5752\(0) = '1' then
                    state_var5920 := Q_WAIT5751;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19273\(80 to 95), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5750;
                  end if;
                when others =>
                  \$19278\ := work.Print.print_string(clk,of_string("unknown primitive"));
                  \$19273\ := "000"& X"000000" & X"1" & eclat_true & \$18788\(0 to 15) & \$18788\(16 to 47) & 
                  work.Int.add(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 95) & \$18788\(96 to 103) & \$18788\(104 to 119) & \$18788\(120 to 121);
                  \$v5752\ := \$ram_lock\;
                  if \$v5752\(0) = '1' then
                    state_var5920 := Q_WAIT5751;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19273\(80 to 95), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5750;
                  end if;
                end case;
              when PAUSE_SET5761 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19280\ := eclat_unit;
                \$v5760\ := \$19215_argument1\;
                case \$v5760\ is
                when "000"& X"000000" & X"0" =>
                  \$19283\ := work.Print.print_string(clk,of_string("======> "));
                  \$19284\ := work.Int.print(clk,\$18788\(16 to 46));
                  \$19285\ := work.Print.print_newline(clk,eclat_unit);
                  \$19281\ := "000"& X"000000" & X"1" & eclat_true & \$18788\(0 to 15) & \$18788\(16 to 47) & 
                  work.Int.add(work.Int.sub(\$18788\(48 to 63), X"000" & X"1"), X"000" & X"1") & \$18788\(64 to 95) & \$18788\(96 to 103) & \$18788\(104 to 119) & \$18788\(120 to 121);
                  \$v5759\ := \$ram_lock\;
                  if \$v5759\(0) = '1' then
                    state_var5920 := Q_WAIT5758;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19281\(80 to 95), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5757;
                  end if;
                when others =>
                  \$19286\ := work.Print.print_string(clk,of_string("unknown primitive"));
                  \$19281\ := "000"& X"000000" & X"1" & eclat_true & \$18788\(0 to 15) & \$18788\(16 to 47) & 
                  work.Int.add(work.Int.sub(\$18788\(48 to 63), X"000" & X"1"), X"000" & X"1") & \$18788\(64 to 95) & \$18788\(96 to 103) & \$18788\(104 to 119) & \$18788\(120 to 121);
                  \$v5759\ := \$ram_lock\;
                  if \$v5759\(0) = '1' then
                    state_var5920 := Q_WAIT5758;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19281\(80 to 95), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5757;
                  end if;
                end case;
              when PAUSE_SET5771 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19289\ := eclat_unit;
                \$v5770\ := \$19215_argument1\;
                case \$v5770\ is
                when "000"& X"000000" & X"0" =>
                  \$19292\ := work.Print.print_string(clk,of_string("======> "));
                  \$19293\ := work.Int.print(clk,\$18788\(16 to 46));
                  \$19294\ := work.Print.print_newline(clk,eclat_unit);
                  \$19290\ := "000"& X"000000" & X"1" & eclat_true & \$18788\(0 to 15) & \$18788\(16 to 47) & 
                  work.Int.add(work.Int.sub(work.Int.sub(\$18788\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1") & \$18788\(64 to 95) & \$18788\(96 to 103) & \$18788\(104 to 119) & \$18788\(120 to 121);
                  \$v5769\ := \$ram_lock\;
                  if \$v5769\(0) = '1' then
                    state_var5920 := Q_WAIT5768;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19290\(80 to 95), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5767;
                  end if;
                when others =>
                  \$19295\ := work.Print.print_string(clk,of_string("unknown primitive"));
                  \$19290\ := "000"& X"000000" & X"1" & eclat_true & \$18788\(0 to 15) & \$18788\(16 to 47) & 
                  work.Int.add(work.Int.sub(work.Int.sub(\$18788\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1") & \$18788\(64 to 95) & \$18788\(96 to 103) & \$18788\(104 to 119) & \$18788\(120 to 121);
                  \$v5769\ := \$ram_lock\;
                  if \$v5769\(0) = '1' then
                    state_var5920 := Q_WAIT5768;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19290\(80 to 95), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5767;
                  end if;
                end case;
              when PAUSE_SET5784 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19299\ := eclat_unit;
                \$v5783\ := \$19215_argument1\;
                case \$v5783\ is
                when "000"& X"000000" & X"0" =>
                  \$19302\ := work.Print.print_string(clk,of_string("======> "));
                  \$19303\ := work.Int.print(clk,\$18788\(16 to 46));
                  \$19304\ := work.Print.print_newline(clk,eclat_unit);
                  \$19300\ := "000"& X"000000" & X"1" & eclat_true & \$18788\(0 to 15) & \$18788\(16 to 47) & 
                  work.Int.add(work.Int.sub(work.Int.sub(work.Int.sub(
                                                         \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1"), X"000" & X"1") & \$18788\(64 to 95) & \$18788\(96 to 103) & \$18788\(104 to 119) & \$18788\(120 to 121);
                  \$v5782\ := \$ram_lock\;
                  if \$v5782\(0) = '1' then
                    state_var5920 := Q_WAIT5781;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19300\(80 to 95), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5780;
                  end if;
                when others =>
                  \$19305\ := work.Print.print_string(clk,of_string("unknown primitive"));
                  \$19300\ := "000"& X"000000" & X"1" & eclat_true & \$18788\(0 to 15) & \$18788\(16 to 47) & 
                  work.Int.add(work.Int.sub(work.Int.sub(work.Int.sub(
                                                         \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1"), X"000" & X"1") & \$18788\(64 to 95) & \$18788\(96 to 103) & \$18788\(104 to 119) & \$18788\(120 to 121);
                  \$v5782\ := \$ram_lock\;
                  if \$v5782\(0) = '1' then
                    state_var5920 := Q_WAIT5781;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19300\(80 to 95), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5780;
                  end if;
                end case;
              when PAUSE_SET5800 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19310\ := eclat_unit;
                \$v5799\ := \$19215_argument1\;
                case \$v5799\ is
                when "000"& X"000000" & X"0" =>
                  \$19313\ := work.Print.print_string(clk,of_string("======> "));
                  \$19314\ := work.Int.print(clk,\$18788\(16 to 46));
                  \$19315\ := work.Print.print_newline(clk,eclat_unit);
                  \$19311\ := "000"& X"000000" & X"1" & eclat_true & \$18788\(0 to 15) & \$18788\(16 to 47) & 
                  work.Int.add(work.Int.sub(work.Int.sub(work.Int.sub(
                                                         work.Int.sub(
                                                         \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1"), X"000" & X"1"), X"000" & X"1") & \$18788\(64 to 95) & \$18788\(96 to 103) & \$18788\(104 to 119) & \$18788\(120 to 121);
                  \$v5798\ := \$ram_lock\;
                  if \$v5798\(0) = '1' then
                    state_var5920 := Q_WAIT5797;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19311\(80 to 95), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5796;
                  end if;
                when others =>
                  \$19316\ := work.Print.print_string(clk,of_string("unknown primitive"));
                  \$19311\ := "000"& X"000000" & X"1" & eclat_true & \$18788\(0 to 15) & \$18788\(16 to 47) & 
                  work.Int.add(work.Int.sub(work.Int.sub(work.Int.sub(
                                                         work.Int.sub(
                                                         \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1"), X"000" & X"1"), X"000" & X"1") & \$18788\(64 to 95) & \$18788\(96 to 103) & \$18788\(104 to 119) & \$18788\(120 to 121);
                  \$v5798\ := \$ram_lock\;
                  if \$v5798\(0) = '1' then
                    state_var5920 := Q_WAIT5797;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19311\(80 to 95), X"000" & X"1")));
                    state_var5920 := PAUSE_GET5796;
                  end if;
                end case;
              when PAUSE_SET5815 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19323\ := eclat_unit;
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"2") & \$19215_argument1\ & eclat_true & 
                work.Int.add(\$18788\(48 to 63), X"000" & X"1") & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_SET5818 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19325\ := eclat_unit;
                result4928 := work.Int.add(\$18788\(0 to 15), X"000" & X"2") & "000"& X"000000" & X"1" & eclat_true & \$18788\(48 to 63) & \$18788\(64 to 119) & \$18788\(120 to 121);
                rdy4929 := eclat_true;
                state_var5920 := IDLE4930;
              when PAUSE_SET5829 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19351\ := eclat_unit;
                \$19347_fill6534389_arg\ := work.Int.add(\$19347_fill6534389_arg\(0 to 15), X"000" & X"1") & 
                work.Int.sub(\$19347_fill6534389_arg\(16 to 31), X"000" & X"1") & \$19347_fill6534389_arg\(32 to 47) & \$19347_fill6534389_arg\(48 to 79);
                state_var5920 := \$19347_FILL6534389\;
              when PAUSE_SET5836 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19345\ := eclat_unit;
                \$19347_fill6534389_id\ := "000010100111";
                \$19347_fill6534389_arg\ := X"000" & X"1" & \$19343_sp\ & eclat_resize(\$19215_argument1\,16) & \$19344\(64 to 95);
                state_var5920 := \$19347_FILL6534389\;
              when PAUSE_SET5839 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19352\ := eclat_unit;
                \$19343_sp\ := work.Int.add(\$18788\(48 to 63), X"000" & X"1");
                \$18793_make_block579_id\ := "000010101000";
                \$18793_make_block579_arg\ := \$19343_sp\ & \$18788\(16 to 47) & \$18788\(64 to 95) & "11110111" & 
                work.Int.add(eclat_resize(\$19215_argument1\,16), X"000" & X"1");
                state_var5920 := \$18793_MAKE_BLOCK579\;
              when PAUSE_SET5855 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19355\ := eclat_unit;
                \$v5854\ := \$ram_lock\;
                if \$v5854\(0) = '1' then
                  state_var5920 := Q_WAIT5853;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(X"3e80", eclat_resize(\$19215_argument1\,16))));
                  state_var5920 := PAUSE_GET5852;
                end if;
              when PAUSE_SET5858 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19365\ := eclat_unit;
                \$19361_fill6544390_arg\ := work.Int.add(\$19361_fill6544390_arg\(0 to 15), X"000" & X"1") & 
                work.Int.sub(\$19361_fill6544390_arg\(16 to 31), X"000" & X"1") & \$19361_fill6544390_arg\(32 to 47) & \$19361_fill6544390_arg\(48 to 79);
                state_var5920 := \$19361_FILL6544390\;
              when PAUSE_SET5865 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19359\ := eclat_unit;
                \$19361_fill6544390_id\ := "000010101001";
                \$19361_fill6544390_arg\ := X"000" & X"1" & \$18788\(48 to 63) & eclat_resize(\$19215_argument1\,16) & \$19358\(64 to 95);
                state_var5920 := \$19361_FILL6544390\;
              when PAUSE_SET5874 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19419\ := eclat_unit;
                \$19416_w36574398_arg\ := work.Int.add(\$19416_w36574398_arg\(0 to 15), X"000" & X"1") & 
                work.Int.add(\$19416_w36574398_arg\(16 to 31), X"000" & X"1") & \$19416_w36574398_arg\(32 to 47) & \$19416_w36574398_arg\(48 to 79);
                state_var5920 := \$19416_W36574398\;
              when PAUSE_SET5878 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19414\ := eclat_unit;
                \$19416_w36574398_id\ := "000010110111";
                \$19416_w36574398_arg\ := X"000" & X"1" & work.Int.add(
                                                          \$19412_sp\, X"000" & X"1") & eclat_resize(\$19215_argument1\,16) & \$19410\(64 to 95);
                state_var5920 := \$19416_W36574398\;
              when PAUSE_SET5881 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19424\ := eclat_unit;
                \$19420_w06554397_arg\ := work.Int.add(\$19420_w06554397_arg\(0 to 15), X"000" & X"1") & 
                work.Int.sub(\$19420_w06554397_arg\(16 to 31), X"000" & X"1") & \$19420_w06554397_arg\(32 to 47) & \$19420_w06554397_arg\(48 to 63) & \$19420_w06554397_arg\(64 to 95);
                state_var5920 := \$19420_W06554397\;
              when PAUSE_SET5888 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19411\ := eclat_unit;
                \$19420_w06554397_id\ := "000010111001";
                \$19420_w06554397_arg\ := X"000" & X"0" & \$19409_sp\ & eclat_resize(\$19215_argument1\,16) & eclat_resize(\$19340_argument2\,16) & \$19410\(64 to 95);
                state_var5920 := \$19420_W06554397\;
              when PAUSE_SET5891 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$19425\ := eclat_unit;
                \$19409_sp\ := work.Int.add(\$18788\(48 to 63), X"000" & X"1");
                \$18793_make_block579_id\ := "000010111010";
                \$18793_make_block579_arg\ := \$19409_sp\ & \$18788\(16 to 47) & \$18788\(64 to 95) & "11110111" & 
                work.Int.add(work.Int.sub(work.Int.mul(X"000" & X"2", eclat_resize(\$19215_argument1\,16)), X"000" & X"1"), eclat_resize(\$19340_argument2\,16));
                state_var5920 := \$18793_MAKE_BLOCK579\;
              when Q_WAIT4932 =>
                \$v4933\ := \$ram_lock\;
                if \$v4933\(0) = '1' then
                  state_var5920 := Q_WAIT4932;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$18790_loop666_arg\(16 to 31), \$18790_loop666_arg\(0 to 15))));
                  \$ram_write\ <= \$19761\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET4931;
                end if;
              when Q_WAIT4935 =>
                \$v4936\ := \$ram_lock\;
                if \$v4936\(0) = '1' then
                  state_var5920 := Q_WAIT4935;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$18790_loop666_arg\(32 to 47), \$18790_loop666_arg\(0 to 15))));
                  state_var5920 := PAUSE_GET4934;
                end if;
              when Q_WAIT4939 =>
                \$v4940\ := \$ram_lock\;
                if \$v4940\(0) = '1' then
                  state_var5920 := Q_WAIT4939;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$18791_loop665_arg\(64 to 79), \$18791_loop665_arg\(0 to 15))));
                  \$ram_write\ <= \$19742\(0 to 31); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET4938;
                end if;
              when Q_WAIT4942 =>
                \$v4943\ := \$ram_lock\;
                if \$v4943\(0) = '1' then
                  state_var5920 := Q_WAIT4942;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$19741\(0 to 30),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$18791_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET4941;
                end if;
              when Q_WAIT4945 =>
                \$v4946\ := \$ram_lock\;
                if \$v4946\(0) = '1' then
                  state_var5920 := Q_WAIT4945;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$19741\(0 to 30),16)));
                  \$ram_write\ <= eclat_resize(\$18791_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET4944;
                end if;
              when Q_WAIT4948 =>
                \$v4949\ := \$ram_lock\;
                if \$v4949\(0) = '1' then
                  state_var5920 := Q_WAIT4948;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18791_loop665_arg\(16 to 31)));
                  \$ram_write\ <= \$19745_hd\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET4947;
                end if;
              when Q_WAIT4951 =>
                \$v4952\ := \$ram_lock\;
                if \$v4952\(0) = '1' then
                  state_var5920 := Q_WAIT4951;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$19741\(0 to 30),16)));
                  state_var5920 := PAUSE_GET4950;
                end if;
              when Q_WAIT4955 =>
                \$v4956\ := \$ram_lock\;
                if \$v4956\(0) = '1' then
                  state_var5920 := Q_WAIT4955;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19741\(0 to 30),16), X"000" & X"1")));
                  state_var5920 := PAUSE_GET4954;
                end if;
              when Q_WAIT4959 =>
                \$v4960\ := \$ram_lock\;
                if \$v4960\(0) = '1' then
                  state_var5920 := Q_WAIT4959;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$18791_loop665_arg\(64 to 79), \$18791_loop665_arg\(0 to 15))));
                  state_var5920 := PAUSE_GET4958;
                end if;
              when Q_WAIT5173 =>
                \$v5174\ := \$ram_lock\;
                if \$v5174\(0) = '1' then
                  state_var5920 := Q_WAIT5173;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$19485\(64 to 79)));
                  \$ram_write\ <= work.Int.lor(work.Int.lsl(eclat_resize(\$18793_make_block579_arg\(80 to 87),31), X"000000" & X"18"), 
                                               work.Int.lsl(eclat_resize(
                                                            eclat_if(
                                                            work.Int.eq(
                                                            \$18793_make_block579_arg\(88 to 103), X"000" & X"0") & X"000" & X"1" & \$18793_make_block579_arg\(88 to 103)),31), X"0000000" & X"2")) & eclat_true; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5172;
                end if;
              when Q_WAIT5176 =>
                \$v5177\ := \$ram_lock\;
                if \$v5177\(0) = '1' then
                  state_var5920 := Q_WAIT5176;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18794_apply638_arg\(60 to 90),16), X"000" & X"0"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5175;
                end if;
              when Q_WAIT5179 =>
                \$v5180\ := \$ram_lock\;
                if \$v5180\(0) = '1' then
                  state_var5920 := Q_WAIT5179;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$19467_sp\));
                  \$ram_write\ <= \$19462\(0 to 31); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5178;
                end if;
              when Q_WAIT5183 =>
                \$v5184\ := \$ram_lock\;
                if \$v5184\(0) = '1' then
                  state_var5920 := Q_WAIT5183;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$19466_sp\));
                  \$ram_write\ <= \$19463\(0 to 31); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5182;
                end if;
              when Q_WAIT5187 =>
                \$v5188\ := \$ram_lock\;
                if \$v5188\(0) = '1' then
                  state_var5920 := Q_WAIT5187;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$19465_sp\));
                  \$ram_write\ <= \$19464\(0 to 31); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5186;
                end if;
              when Q_WAIT5191 =>
                \$v5192\ := \$ram_lock\;
                if \$v5192\(0) = '1' then
                  state_var5920 := Q_WAIT5191;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          \$19464\(32 to 47), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(work.Int.add(\$18794_apply638_arg\(44 to 59), X"000" & X"1"),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5190;
                end if;
              when Q_WAIT5194 =>
                \$v5195\ := \$ram_lock\;
                if \$v5195\(0) = '1' then
                  state_var5920 := Q_WAIT5194;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$19464\(32 to 47), X"000" & X"1")));
                  \$ram_write\ <= \$18794_apply638_arg\(110 to 141); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5193;
                end if;
              when Q_WAIT5197 =>
                \$v5198\ := \$ram_lock\;
                if \$v5198\(0) = '1' then
                  state_var5920 := Q_WAIT5197;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$19464\(32 to 47)));
                  \$ram_write\ <= eclat_resize(\$18794_apply638_arg\(142 to 149),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5196;
                end if;
              when Q_WAIT5201 =>
                \$v5202\ := \$ram_lock\;
                if \$v5202\(0) = '1' then
                  state_var5920 := Q_WAIT5201;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19463\(32 to 47), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5200;
                end if;
              when Q_WAIT5205 =>
                \$v5206\ := \$ram_lock\;
                if \$v5206\(0) = '1' then
                  state_var5920 := Q_WAIT5205;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19462\(32 to 47), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5204;
                end if;
              when Q_WAIT5209 =>
                \$v5210\ := \$ram_lock\;
                if \$v5210\(0) = '1' then
                  state_var5920 := Q_WAIT5209;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18794_apply638_arg\(92 to 107), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5208;
                end if;
              when Q_WAIT5214 =>
                \$v5215\ := \$ram_lock\;
                if \$v5215\(0) = '1' then
                  state_var5920 := Q_WAIT5214;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$19444\(64 to 94),16), X"000" & X"2"), X"000" & X"1")));
                  \$ram_write\ <= \$19448_v\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5213;
                end if;
              when Q_WAIT5217 =>
                \$v5218\ := \$ram_lock\;
                if \$v5218\(0) = '1' then
                  state_var5920 := Q_WAIT5217;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19446_sp\, X"000" & X"1")));
                  state_var5920 := PAUSE_GET5216;
                end if;
              when Q_WAIT5221 =>
                \$v5222\ := \$ram_lock\;
                if \$v5222\(0) = '1' then
                  state_var5920 := Q_WAIT5221;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$19444\(64 to 94),16), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= \$19450_v\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5220;
                end if;
              when Q_WAIT5224 =>
                \$v5225\ := \$ram_lock\;
                if \$v5225\(0) = '1' then
                  state_var5920 := Q_WAIT5224;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18796_make_block_n646_arg\(16 to 31), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5223;
                end if;
              when Q_WAIT5228 =>
                \$v5229\ := \$ram_lock\;
                if \$v5229\(0) = '1' then
                  state_var5920 := Q_WAIT5228;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$19444\(64 to 94),16), X"000" & X"0"), X"000" & X"1")));
                  \$ram_write\ <= \$19444\(0 to 31); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5227;
                end if;
              when Q_WAIT5232 =>
                \$v5233\ := \$code_lock\;
                if \$v5233\(0) = '1' then
                  state_var5920 := Q_WAIT5232;
                else
                  acquire(\$code_lock\);
                  \$code_ptr\ <= to_integer(unsigned(work.Int.add(\$18797_branch_if648_arg\(1 to 16), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5231;
                end if;
              when Q_WAIT5236 =>
                \$v5237\ := \$ram_lock\;
                if \$v5237\(0) = '1' then
                  state_var5920 := Q_WAIT5236;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.sub(
                                                          work.Int.sub(
                                                          work.Int.sub(
                                                          \$18798_w652_arg\(16 to 31), \$18798_w652_arg\(32 to 47)), \$18798_w652_arg\(48 to 63)), \$18798_w652_arg\(0 to 15))));
                  \$ram_write\ <= \$19437\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5235;
                end if;
              when Q_WAIT5239 =>
                \$v5240\ := \$ram_lock\;
                if \$v5240\(0) = '1' then
                  state_var5920 := Q_WAIT5239;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18798_w652_arg\(16 to 31), \$18798_w652_arg\(0 to 15))));
                  state_var5920 := PAUSE_GET5238;
                end if;
              when Q_WAIT5243 =>
                \$v5244\ := \$ram_lock\;
                if \$v5244\(0) = '1' then
                  state_var5920 := Q_WAIT5243;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$18799_w1656_arg\(48 to 78),16), 
                                                          work.Int.mul(
                                                          X"000" & X"2", \$18799_w1656_arg\(0 to 15))), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(work.Int.add(work.Int.add(
                                                            \$18799_w1656_arg\(16 to 31), X"000" & X"2"), eclat_resize(\$19433\,16)),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5242;
                end if;
              when Q_WAIT5246 =>
                \$v5247\ := \$code_lock\;
                if \$v5247\(0) = '1' then
                  state_var5920 := Q_WAIT5246;
                else
                  acquire(\$code_lock\);
                  \$code_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                  \$18799_w1656_arg\(16 to 31), X"000" & X"3"), \$18799_w1656_arg\(0 to 15))));
                  state_var5920 := PAUSE_GET5245;
                end if;
              when Q_WAIT5249 =>
                \$v5250\ := \$ram_lock\;
                if \$v5250\(0) = '1' then
                  state_var5920 := Q_WAIT5249;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$18799_w1656_arg\(48 to 78),16), 
                                                          work.Int.sub(
                                                          work.Int.mul(
                                                          X"000" & X"2", \$18799_w1656_arg\(0 to 15)), X"000" & X"1")), X"000" & X"1")));
                  \$ram_write\ <= work.Int.lor(work.Int.lsl(eclat_resize("11111001",31), X"000000" & X"18"), 
                                               work.Int.lsl(eclat_resize(
                                                            work.Int.mul(
                                                            X"000" & X"2", \$18799_w1656_arg\(0 to 15)),31), X"0000000" & X"2")) & eclat_true; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5248;
                end if;
              when Q_WAIT5253 =>
                \$v5254\ := \$ram_lock\;
                if \$v5254\(0) = '1' then
                  state_var5920 := Q_WAIT5253;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$18788\(48 to 63), X"000" & X"0"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5252;
                end if;
              when Q_WAIT5256 =>
                \$v5257\ := \$ram_lock\;
                if \$v5257\(0) = '1' then
                  state_var5920 := Q_WAIT5256;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5255;
                end if;
              when Q_WAIT5259 =>
                \$v5260\ := \$ram_lock\;
                if \$v5260\(0) = '1' then
                  state_var5920 := Q_WAIT5259;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$18788\(48 to 63), X"000" & X"2"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5258;
                end if;
              when Q_WAIT5262 =>
                \$v5263\ := \$ram_lock\;
                if \$v5263\(0) = '1' then
                  state_var5920 := Q_WAIT5262;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$18788\(48 to 63), X"000" & X"3"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5261;
                end if;
              when Q_WAIT5265 =>
                \$v5266\ := \$ram_lock\;
                if \$v5266\(0) = '1' then
                  state_var5920 := Q_WAIT5265;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$18788\(48 to 63), X"000" & X"4"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5264;
                end if;
              when Q_WAIT5268 =>
                \$v5269\ := \$ram_lock\;
                if \$v5269\(0) = '1' then
                  state_var5920 := Q_WAIT5268;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$18788\(48 to 63), X"000" & X"5"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5267;
                end if;
              when Q_WAIT5271 =>
                \$v5272\ := \$ram_lock\;
                if \$v5272\(0) = '1' then
                  state_var5920 := Q_WAIT5271;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$18788\(48 to 63), X"000" & X"6"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5270;
                end if;
              when Q_WAIT5274 =>
                \$v5275\ := \$ram_lock\;
                if \$v5275\(0) = '1' then
                  state_var5920 := Q_WAIT5274;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$18788\(48 to 63), X"000" & X"7"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5273;
                end if;
              when Q_WAIT5277 =>
                \$v5278\ := \$ram_lock\;
                if \$v5278\(0) = '1' then
                  state_var5920 := Q_WAIT5277;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5276;
                end if;
              when Q_WAIT5280 =>
                \$v5281\ := \$ram_lock\;
                if \$v5281\(0) = '1' then
                  state_var5920 := Q_WAIT5280;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5279;
                end if;
              when Q_WAIT5283 =>
                \$v5284\ := \$ram_lock\;
                if \$v5284\(0) = '1' then
                  state_var5920 := Q_WAIT5283;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5282;
                end if;
              when Q_WAIT5286 =>
                \$v5287\ := \$ram_lock\;
                if \$v5287\(0) = '1' then
                  state_var5920 := Q_WAIT5286;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5285;
                end if;
              when Q_WAIT5289 =>
                \$v5290\ := \$ram_lock\;
                if \$v5290\(0) = '1' then
                  state_var5920 := Q_WAIT5289;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"2"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5288;
                end if;
              when Q_WAIT5292 =>
                \$v5293\ := \$ram_lock\;
                if \$v5293\(0) = '1' then
                  state_var5920 := Q_WAIT5292;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5291;
                end if;
              when Q_WAIT5295 =>
                \$v5296\ := \$ram_lock\;
                if \$v5296\(0) = '1' then
                  state_var5920 := Q_WAIT5295;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"3"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5294;
                end if;
              when Q_WAIT5298 =>
                \$v5299\ := \$ram_lock\;
                if \$v5299\(0) = '1' then
                  state_var5920 := Q_WAIT5298;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5297;
                end if;
              when Q_WAIT5301 =>
                \$v5302\ := \$ram_lock\;
                if \$v5302\(0) = '1' then
                  state_var5920 := Q_WAIT5301;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"4"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5300;
                end if;
              when Q_WAIT5304 =>
                \$v5305\ := \$ram_lock\;
                if \$v5305\(0) = '1' then
                  state_var5920 := Q_WAIT5304;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5303;
                end if;
              when Q_WAIT5307 =>
                \$v5308\ := \$ram_lock\;
                if \$v5308\(0) = '1' then
                  state_var5920 := Q_WAIT5307;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"5"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5306;
                end if;
              when Q_WAIT5310 =>
                \$v5311\ := \$ram_lock\;
                if \$v5311\(0) = '1' then
                  state_var5920 := Q_WAIT5310;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5309;
                end if;
              when Q_WAIT5313 =>
                \$v5314\ := \$ram_lock\;
                if \$v5314\(0) = '1' then
                  state_var5920 := Q_WAIT5313;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"6"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5312;
                end if;
              when Q_WAIT5316 =>
                \$v5317\ := \$ram_lock\;
                if \$v5317\(0) = '1' then
                  state_var5920 := Q_WAIT5316;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5315;
                end if;
              when Q_WAIT5319 =>
                \$v5320\ := \$ram_lock\;
                if \$v5320\(0) = '1' then
                  state_var5920 := Q_WAIT5319;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"7"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5318;
                end if;
              when Q_WAIT5322 =>
                \$v5323\ := \$ram_lock\;
                if \$v5323\(0) = '1' then
                  state_var5920 := Q_WAIT5322;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5321;
                end if;
              when Q_WAIT5325 =>
                \$v5326\ := \$ram_lock\;
                if \$v5326\(0) = '1' then
                  state_var5920 := Q_WAIT5325;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18788\(64 to 94),16), 
                                                                 work.Int.sub(
                                                                 X"000" & X"1", X"000" & X"1")), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5324;
                end if;
              when Q_WAIT5328 =>
                \$v5329\ := \$ram_lock\;
                if \$v5329\(0) = '1' then
                  state_var5920 := Q_WAIT5328;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18788\(64 to 94),16), 
                                                                 work.Int.sub(
                                                                 X"000" & X"2", X"000" & X"1")), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5327;
                end if;
              when Q_WAIT5331 =>
                \$v5332\ := \$ram_lock\;
                if \$v5332\(0) = '1' then
                  state_var5920 := Q_WAIT5331;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18788\(64 to 94),16), 
                                                                 work.Int.sub(
                                                                 X"000" & X"3", X"000" & X"1")), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5330;
                end if;
              when Q_WAIT5334 =>
                \$v5335\ := \$ram_lock\;
                if \$v5335\(0) = '1' then
                  state_var5920 := Q_WAIT5334;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18788\(64 to 94),16), 
                                                                 work.Int.sub(
                                                                 X"000" & X"4", X"000" & X"1")), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5333;
                end if;
              when Q_WAIT5337 =>
                \$v5338\ := \$ram_lock\;
                if \$v5338\(0) = '1' then
                  state_var5920 := Q_WAIT5337;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18788\(64 to 94),16), 
                                                                 work.Int.sub(
                                                                 X"000" & X"1", X"000" & X"1")), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5336;
                end if;
              when Q_WAIT5340 =>
                \$v5341\ := \$ram_lock\;
                if \$v5341\(0) = '1' then
                  state_var5920 := Q_WAIT5340;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5339;
                end if;
              when Q_WAIT5343 =>
                \$v5344\ := \$ram_lock\;
                if \$v5344\(0) = '1' then
                  state_var5920 := Q_WAIT5343;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18788\(64 to 94),16), 
                                                                 work.Int.sub(
                                                                 X"000" & X"2", X"000" & X"1")), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5342;
                end if;
              when Q_WAIT5346 =>
                \$v5347\ := \$ram_lock\;
                if \$v5347\(0) = '1' then
                  state_var5920 := Q_WAIT5346;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5345;
                end if;
              when Q_WAIT5349 =>
                \$v5350\ := \$ram_lock\;
                if \$v5350\(0) = '1' then
                  state_var5920 := Q_WAIT5349;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18788\(64 to 94),16), 
                                                                 work.Int.sub(
                                                                 X"000" & X"3", X"000" & X"1")), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5348;
                end if;
              when Q_WAIT5352 =>
                \$v5353\ := \$ram_lock\;
                if \$v5353\(0) = '1' then
                  state_var5920 := Q_WAIT5352;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5351;
                end if;
              when Q_WAIT5355 =>
                \$v5356\ := \$ram_lock\;
                if \$v5356\(0) = '1' then
                  state_var5920 := Q_WAIT5355;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18788\(64 to 94),16), 
                                                                 work.Int.sub(
                                                                 X"000" & X"4", X"000" & X"1")), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5354;
                end if;
              when Q_WAIT5358 =>
                \$v5359\ := \$ram_lock\;
                if \$v5359\(0) = '1' then
                  state_var5920 := Q_WAIT5358;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5357;
                end if;
              when Q_WAIT5361 =>
                \$v5362\ := \$ram_lock\;
                if \$v5362\(0) = '1' then
                  state_var5920 := Q_WAIT5361;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18788\(64 to 94),16), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5360;
                end if;
              when Q_WAIT5364 =>
                \$v5365\ := \$ram_lock\;
                if \$v5365\(0) = '1' then
                  state_var5920 := Q_WAIT5364;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18856_loop_push6494360_arg\(0 to 15)));
                  \$ram_write\ <= \$18859\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5363;
                end if;
              when Q_WAIT5367 =>
                \$v5368\ := \$ram_lock\;
                if \$v5368\(0) = '1' then
                  state_var5920 := Q_WAIT5367;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18856_loop_push6494360_arg\(24 to 54),16), eclat_resize(
                                                                 work.Int.add(
                                                                 \$18856_loop_push6494360_arg\(16 to 23), "00000010"),16)), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5366;
                end if;
              when Q_WAIT5371 =>
                \$v5372\ := \$ram_lock\;
                if \$v5372\(0) = '1' then
                  state_var5920 := Q_WAIT5371;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18788\(64 to 94),16)));
                  state_var5920 := PAUSE_GET5370;
                end if;
              when Q_WAIT5374 =>
                \$v5375\ := \$ram_lock\;
                if \$v5375\(0) = '1' then
                  state_var5920 := Q_WAIT5374;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5373;
                end if;
              when Q_WAIT5377 =>
                \$v5378\ := \$ram_lock\;
                if \$v5378\(0) = '1' then
                  state_var5920 := Q_WAIT5377;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5376;
                end if;
              when Q_WAIT5380 =>
                \$v5381\ := \$ram_lock\;
                if \$v5381\(0) = '1' then
                  state_var5920 := Q_WAIT5380;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5379;
                end if;
              when Q_WAIT5383 =>
                \$v5384\ := \$ram_lock\;
                if \$v5384\(0) = '1' then
                  state_var5920 := Q_WAIT5383;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5382;
                end if;
              when Q_WAIT5386 =>
                \$v5387\ := \$ram_lock\;
                if \$v5387\(0) = '1' then
                  state_var5920 := Q_WAIT5386;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18788\(16 to 46),16), X"000" & X"0"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5385;
                end if;
              when Q_WAIT5389 =>
                \$v5390\ := \$ram_lock\;
                if \$v5390\(0) = '1' then
                  state_var5920 := Q_WAIT5389;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18788\(16 to 46),16), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5388;
                end if;
              when Q_WAIT5392 =>
                \$v5393\ := \$ram_lock\;
                if \$v5393\(0) = '1' then
                  state_var5920 := Q_WAIT5392;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18788\(16 to 46),16), X"000" & X"2"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5391;
                end if;
              when Q_WAIT5395 =>
                \$v5396\ := \$ram_lock\;
                if \$v5396\(0) = '1' then
                  state_var5920 := Q_WAIT5395;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18788\(16 to 46),16), X"000" & X"3"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5394;
                end if;
              when Q_WAIT5398 =>
                \$v5399\ := \$ram_lock\;
                if \$v5399\(0) = '1' then
                  state_var5920 := Q_WAIT5398;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$18788\(16 to 46),16), X"000" & X"0"), X"000" & X"1")));
                  \$ram_write\ <= \$18873_v\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5397;
                end if;
              when Q_WAIT5401 =>
                \$v5402\ := \$ram_lock\;
                if \$v5402\(0) = '1' then
                  state_var5920 := Q_WAIT5401;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18788\(48 to 63), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5400;
                end if;
              when Q_WAIT5404 =>
                \$v5405\ := \$ram_lock\;
                if \$v5405\(0) = '1' then
                  state_var5920 := Q_WAIT5404;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$18788\(16 to 46),16), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= \$18875_v\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5403;
                end if;
              when Q_WAIT5407 =>
                \$v5408\ := \$ram_lock\;
                if \$v5408\(0) = '1' then
                  state_var5920 := Q_WAIT5407;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18788\(48 to 63), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5406;
                end if;
              when Q_WAIT5410 =>
                \$v5411\ := \$ram_lock\;
                if \$v5411\(0) = '1' then
                  state_var5920 := Q_WAIT5410;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$18788\(16 to 46),16), X"000" & X"2"), X"000" & X"1")));
                  \$ram_write\ <= \$18877_v\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5409;
                end if;
              when Q_WAIT5413 =>
                \$v5414\ := \$ram_lock\;
                if \$v5414\(0) = '1' then
                  state_var5920 := Q_WAIT5413;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18788\(48 to 63), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5412;
                end if;
              when Q_WAIT5416 =>
                \$v5417\ := \$ram_lock\;
                if \$v5417\(0) = '1' then
                  state_var5920 := Q_WAIT5416;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$18788\(16 to 46),16), X"000" & X"3"), X"000" & X"1")));
                  \$ram_write\ <= \$18879_v\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5415;
                end if;
              when Q_WAIT5419 =>
                \$v5420\ := \$ram_lock\;
                if \$v5420\(0) = '1' then
                  state_var5920 := Q_WAIT5419;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18788\(48 to 63), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5418;
                end if;
              when Q_WAIT5422 =>
                \$v5423\ := \$ram_lock\;
                if \$v5423\(0) = '1' then
                  state_var5920 := Q_WAIT5422;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18788\(16 to 46),16)));
                  state_var5920 := PAUSE_GET5421;
                end if;
              when Q_WAIT5425 =>
                \$v5426\ := \$ram_lock\;
                if \$v5426\(0) = '1' then
                  state_var5920 := Q_WAIT5425;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18788\(16 to 46),16), eclat_resize(\$18882_v\(0 to 30),16)), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5424;
                end if;
              when Q_WAIT5428 =>
                \$v5429\ := \$ram_lock\;
                if \$v5429\(0) = '1' then
                  state_var5920 := Q_WAIT5428;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18788\(48 to 63), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5427;
                end if;
              when Q_WAIT5431 =>
                \$v5432\ := \$ram_lock\;
                if \$v5432\(0) = '1' then
                  state_var5920 := Q_WAIT5431;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$18788\(16 to 46),16), eclat_resize(\$18884_v\(0 to 30),16)), X"000" & X"1")));
                  \$ram_write\ <= \$18885_v\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5430;
                end if;
              when Q_WAIT5434 =>
                \$v5435\ := \$ram_lock\;
                if \$v5435\(0) = '1' then
                  state_var5920 := Q_WAIT5434;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5433;
                end if;
              when Q_WAIT5437 =>
                \$v5438\ := \$ram_lock\;
                if \$v5438\(0) = '1' then
                  state_var5920 := Q_WAIT5437;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18788\(48 to 63), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5436;
                end if;
              when Q_WAIT5440 =>
                \$v5441\ := \$ram_lock\;
                if \$v5441\(0) = '1' then
                  state_var5920 := Q_WAIT5440;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18788\(16 to 46),16), eclat_resize(\$18887_v\(0 to 30),16)), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5439;
                end if;
              when Q_WAIT5443 =>
                \$v5444\ := \$ram_lock\;
                if \$v5444\(0) = '1' then
                  state_var5920 := Q_WAIT5443;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18788\(48 to 63), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5442;
                end if;
              when Q_WAIT5446 =>
                \$v5447\ := \$ram_lock\;
                if \$v5447\(0) = '1' then
                  state_var5920 := Q_WAIT5446;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$18788\(16 to 46),16), eclat_resize(\$18889_v\(0 to 30),16)), X"000" & X"1")));
                  \$ram_write\ <= \$18890_v\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5445;
                end if;
              when Q_WAIT5449 =>
                \$v5450\ := \$ram_lock\;
                if \$v5450\(0) = '1' then
                  state_var5920 := Q_WAIT5449;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5448;
                end if;
              when Q_WAIT5452 =>
                \$v5453\ := \$ram_lock\;
                if \$v5453\(0) = '1' then
                  state_var5920 := Q_WAIT5452;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18788\(48 to 63), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5451;
                end if;
              when Q_WAIT5455 =>
                \$v5456\ := \$ram_lock\;
                if \$v5456\(0) = '1' then
                  state_var5920 := Q_WAIT5455;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5454;
                end if;
              when Q_WAIT5458 =>
                \$v5459\ := \$ram_lock\;
                if \$v5459\(0) = '1' then
                  state_var5920 := Q_WAIT5458;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$18788\(104 to 119), X"000" & X"1"), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5457;
                end if;
              when Q_WAIT5461 =>
                \$v5462\ := \$ram_lock\;
                if \$v5462\(0) = '1' then
                  state_var5920 := Q_WAIT5461;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$18788\(104 to 119), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5460;
                end if;
              when Q_WAIT5464 =>
                \$v5465\ := \$ram_lock\;
                if \$v5465\(0) = '1' then
                  state_var5920 := Q_WAIT5464;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$18788\(104 to 119), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5463;
                end if;
              when Q_WAIT5467 =>
                \$v5468\ := \$ram_lock\;
                if \$v5468\(0) = '1' then
                  state_var5920 := Q_WAIT5467;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18788\(104 to 119), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5466;
                end if;
              when Q_WAIT5470 =>
                \$v5471\ := \$ram_lock\;
                if \$v5471\(0) = '1' then
                  state_var5920 := Q_WAIT5470;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5469;
                end if;
              when Q_WAIT5473 =>
                \$v5474\ := \$ram_lock\;
                if \$v5474\(0) = '1' then
                  state_var5920 := Q_WAIT5473;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5472;
                end if;
              when Q_WAIT5476 =>
                \$v5477\ := \$ram_lock\;
                if \$v5477\(0) = '1' then
                  state_var5920 := Q_WAIT5476;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5475;
                end if;
              when Q_WAIT5479 =>
                \$v5480\ := \$ram_lock\;
                if \$v5480\(0) = '1' then
                  state_var5920 := Q_WAIT5479;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5478;
                end if;
              when Q_WAIT5489 =>
                \$v5490\ := \$ram_lock\;
                if \$v5490\(0) = '1' then
                  state_var5920 := Q_WAIT5489;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18901_binop_int6434361_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5488;
                end if;
              when Q_WAIT5499 =>
                \$v5500\ := \$ram_lock\;
                if \$v5500\(0) = '1' then
                  state_var5920 := Q_WAIT5499;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18920_binop_int6434362_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5498;
                end if;
              when Q_WAIT5509 =>
                \$v5510\ := \$ram_lock\;
                if \$v5510\(0) = '1' then
                  state_var5920 := Q_WAIT5509;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18939_binop_int6434363_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5508;
                end if;
              when Q_WAIT5519 =>
                \$v5520\ := \$ram_lock\;
                if \$v5520\(0) = '1' then
                  state_var5920 := Q_WAIT5519;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18958_binop_int6434364_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5518;
                end if;
              when Q_WAIT5529 =>
                \$v5530\ := \$ram_lock\;
                if \$v5530\(0) = '1' then
                  state_var5920 := Q_WAIT5529;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18977_binop_int6434365_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5528;
                end if;
              when Q_WAIT5539 =>
                \$v5540\ := \$ram_lock\;
                if \$v5540\(0) = '1' then
                  state_var5920 := Q_WAIT5539;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18996_binop_int6434366_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5538;
                end if;
              when Q_WAIT5549 =>
                \$v5550\ := \$ram_lock\;
                if \$v5550\(0) = '1' then
                  state_var5920 := Q_WAIT5549;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19015_binop_int6434367_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5548;
                end if;
              when Q_WAIT5559 =>
                \$v5560\ := \$ram_lock\;
                if \$v5560\(0) = '1' then
                  state_var5920 := Q_WAIT5559;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19034_binop_int6434368_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5558;
                end if;
              when Q_WAIT5569 =>
                \$v5570\ := \$ram_lock\;
                if \$v5570\(0) = '1' then
                  state_var5920 := Q_WAIT5569;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19053_binop_int6434369_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5568;
                end if;
              when Q_WAIT5579 =>
                \$v5580\ := \$ram_lock\;
                if \$v5580\(0) = '1' then
                  state_var5920 := Q_WAIT5579;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19072_binop_int6434370_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5578;
                end if;
              when Q_WAIT5589 =>
                \$v5590\ := \$ram_lock\;
                if \$v5590\(0) = '1' then
                  state_var5920 := Q_WAIT5589;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19091_binop_int6434371_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5588;
                end if;
              when Q_WAIT5599 =>
                \$v5600\ := \$ram_lock\;
                if \$v5600\(0) = '1' then
                  state_var5920 := Q_WAIT5599;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19116_binop_int6434373_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5598;
                end if;
              when Q_WAIT5609 =>
                \$v5610\ := \$ram_lock\;
                if \$v5610\(0) = '1' then
                  state_var5920 := Q_WAIT5609;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19135_binop_int6434374_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5608;
                end if;
              when Q_WAIT5613 =>
                \$v5614\ := \$ram_lock\;
                if \$v5614\(0) = '1' then
                  state_var5920 := Q_WAIT5613;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19166_binop_compare6454377_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5612;
                end if;
              when Q_WAIT5617 =>
                \$v5618\ := \$ram_lock\;
                if \$v5618\(0) = '1' then
                  state_var5920 := Q_WAIT5617;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19174_binop_compare6454378_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5616;
                end if;
              when Q_WAIT5621 =>
                \$v5622\ := \$ram_lock\;
                if \$v5622\(0) = '1' then
                  state_var5920 := Q_WAIT5621;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19182_binop_compare6454379_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5620;
                end if;
              when Q_WAIT5625 =>
                \$v5626\ := \$ram_lock\;
                if \$v5626\(0) = '1' then
                  state_var5920 := Q_WAIT5625;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19190_binop_compare6454380_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5624;
                end if;
              when Q_WAIT5629 =>
                \$v5630\ := \$ram_lock\;
                if \$v5630\(0) = '1' then
                  state_var5920 := Q_WAIT5629;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19198_binop_compare6454381_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5628;
                end if;
              when Q_WAIT5633 =>
                \$v5634\ := \$ram_lock\;
                if \$v5634\(0) = '1' then
                  state_var5920 := Q_WAIT5633;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19206_binop_compare6454382_arg\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5632;
                end if;
              when Q_WAIT5636 =>
                \$v5637\ := \$ram_lock\;
                if \$v5637\(0) = '1' then
                  state_var5920 := Q_WAIT5636;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$18788\(48 to 63), eclat_resize(\$19215_argument1\,16)), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5635;
                end if;
              when Q_WAIT5639 =>
                \$v5640\ := \$ram_lock\;
                if \$v5640\(0) = '1' then
                  state_var5920 := Q_WAIT5639;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$18788\(48 to 63), X"000" & X"1"), eclat_resize(\$19215_argument1\,16)), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5638;
                end if;
              when Q_WAIT5642 =>
                \$v5643\ := \$ram_lock\;
                if \$v5643\(0) = '1' then
                  state_var5920 := Q_WAIT5642;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5641;
                end if;
              when Q_WAIT5645 =>
                \$v5646\ := \$ram_lock\;
                if \$v5646\(0) = '1' then
                  state_var5920 := Q_WAIT5645;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.sub(
                                                          work.Int.sub(
                                                          \$18788\(48 to 63), X"000" & X"1"), eclat_resize(\$19215_argument1\,16))));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5644;
                end if;
              when Q_WAIT5648 =>
                \$v5649\ := \$ram_lock\;
                if \$v5649\(0) = '1' then
                  state_var5920 := Q_WAIT5648;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18788\(64 to 94),16), 
                                                                 work.Int.sub(
                                                                 eclat_resize(\$19215_argument1\,16), X"000" & X"1")), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5647;
                end if;
              when Q_WAIT5651 =>
                \$v5652\ := \$ram_lock\;
                if \$v5652\(0) = '1' then
                  state_var5920 := Q_WAIT5651;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18788\(64 to 94),16), 
                                                                 work.Int.sub(
                                                                 eclat_resize(\$19215_argument1\,16), X"000" & X"1")), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5650;
                end if;
              when Q_WAIT5654 =>
                \$v5655\ := \$ram_lock\;
                if \$v5655\(0) = '1' then
                  state_var5920 := Q_WAIT5654;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5653;
                end if;
              when Q_WAIT5657 =>
                \$v5658\ := \$ram_lock\;
                if \$v5658\(0) = '1' then
                  state_var5920 := Q_WAIT5657;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(work.Int.add(work.Int.add(
                                                            \$18788\(0 to 15), X"000" & X"1"), eclat_resize(\$19215_argument1\,16)),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5656;
                end if;
              when Q_WAIT5660 =>
                \$v5661\ := \$ram_lock\;
                if \$v5661\(0) = '1' then
                  state_var5920 := Q_WAIT5660;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$18788\(48 to 63), X"000" & X"1")));
                  \$ram_write\ <= \$18788\(64 to 95); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5659;
                end if;
              when Q_WAIT5663 =>
                \$v5664\ := \$ram_lock\;
                if \$v5664\(0) = '1' then
                  state_var5920 := Q_WAIT5663;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= eclat_resize(\$18788\(96 to 103),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5662;
                end if;
              when Q_WAIT5666 =>
                \$v5667\ := \$ram_lock\;
                if \$v5667\(0) = '1' then
                  state_var5920 := Q_WAIT5666;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18788\(16 to 46),16), X"000" & X"0"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5665;
                end if;
              when Q_WAIT5669 =>
                \$v5670\ := \$ram_lock\;
                if \$v5670\(0) = '1' then
                  state_var5920 := Q_WAIT5669;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18788\(16 to 46),16), X"000" & X"0"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5668;
                end if;
              when Q_WAIT5672 =>
                \$v5673\ := \$ram_lock\;
                if \$v5673\(0) = '1' then
                  state_var5920 := Q_WAIT5672;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$18788\(48 to 63), eclat_resize(\$19215_argument1\,16)), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5671;
                end if;
              when Q_WAIT5675 =>
                \$v5676\ := \$ram_lock\;
                if \$v5676\(0) = '1' then
                  state_var5920 := Q_WAIT5675;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$18788\(48 to 63), eclat_resize(\$19215_argument1\,16)), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5674;
                end if;
              when Q_WAIT5678 =>
                \$v5679\ := \$ram_lock\;
                if \$v5679\(0) = '1' then
                  state_var5920 := Q_WAIT5678;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$18788\(48 to 63), eclat_resize(\$19215_argument1\,16)), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5677;
                end if;
              when Q_WAIT5682 =>
                \$v5683\ := \$ram_lock\;
                if \$v5683\(0) = '1' then
                  state_var5920 := Q_WAIT5682;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$19234_sp\, X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5681;
                end if;
              when Q_WAIT5685 =>
                \$v5686\ := \$ram_lock\;
                if \$v5686\(0) = '1' then
                  state_var5920 := Q_WAIT5685;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$19234_sp\, X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5684;
                end if;
              when Q_WAIT5688 =>
                \$v5689\ := \$ram_lock\;
                if \$v5689\(0) = '1' then
                  state_var5920 := Q_WAIT5688;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19234_sp\, X"000" & X"1")));
                  state_var5920 := PAUSE_GET5687;
                end if;
              when Q_WAIT5691 =>
                \$v5692\ := \$ram_lock\;
                if \$v5692\(0) = '1' then
                  state_var5920 := Q_WAIT5691;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$19238_w6514383_arg\(32 to 62),16), eclat_resize(
                                                          work.Int.add(
                                                          \$19238_w6514383_arg\(0 to 7), "00000010"),16)), X"000" & X"1")));
                  \$ram_write\ <= \$19241_v\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5690;
                end if;
              when Q_WAIT5694 =>
                \$v5695\ := \$ram_lock\;
                if \$v5695\(0) = '1' then
                  state_var5920 := Q_WAIT5694;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19238_w6514383_arg\(8 to 23), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5693;
                end if;
              when Q_WAIT5698 =>
                \$v5699\ := \$ram_lock\;
                if \$v5699\(0) = '1' then
                  state_var5920 := Q_WAIT5698;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$19231\(64 to 94),16), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= \$19231\(32 to 63); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5697;
                end if;
              when Q_WAIT5701 =>
                \$v5702\ := \$ram_lock\;
                if \$v5702\(0) = '1' then
                  state_var5920 := Q_WAIT5701;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$19231\(64 to 94),16), X"000" & X"0"), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(work.Int.sub(work.Int.add(
                                                            \$18788\(0 to 15), X"000" & X"2"), X"000" & X"3"),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5700;
                end if;
              when Q_WAIT5705 =>
                \$v5706\ := \$ram_lock\;
                if \$v5706\(0) = '1' then
                  state_var5920 := Q_WAIT5705;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5704;
                end if;
              when Q_WAIT5708 =>
                \$v5709\ := \$ram_lock\;
                if \$v5709\(0) = '1' then
                  state_var5920 := Q_WAIT5708;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(X"3e80", eclat_resize(\$19215_argument1\,16))));
                  state_var5920 := PAUSE_GET5707;
                end if;
              when Q_WAIT5711 =>
                \$v5712\ := \$ram_lock\;
                if \$v5712\(0) = '1' then
                  state_var5920 := Q_WAIT5711;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(X"3e80", eclat_resize(\$19215_argument1\,16))));
                  state_var5920 := PAUSE_GET5710;
                end if;
              when Q_WAIT5714 =>
                \$v5715\ := \$ram_lock\;
                if \$v5715\(0) = '1' then
                  state_var5920 := Q_WAIT5714;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5713;
                end if;
              when Q_WAIT5717 =>
                \$v5718\ := \$ram_lock\;
                if \$v5718\(0) = '1' then
                  state_var5920 := Q_WAIT5717;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          X"3e80", eclat_resize(\$19215_argument1\,16))));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5716;
                end if;
              when Q_WAIT5720 =>
                \$v5721\ := \$ram_lock\;
                if \$v5721\(0) = '1' then
                  state_var5920 := Q_WAIT5720;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5719;
                end if;
              when Q_WAIT5723 =>
                \$v5724\ := \$ram_lock\;
                if \$v5724\(0) = '1' then
                  state_var5920 := Q_WAIT5723;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18788\(16 to 46),16), eclat_resize(\$19215_argument1\,16)), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5722;
                end if;
              when Q_WAIT5726 =>
                \$v5727\ := \$ram_lock\;
                if \$v5727\(0) = '1' then
                  state_var5920 := Q_WAIT5726;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$18788\(16 to 46),16), eclat_resize(\$19215_argument1\,16)), X"000" & X"1")));
                  \$ram_write\ <= \$19257_v\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5725;
                end if;
              when Q_WAIT5729 =>
                \$v5730\ := \$ram_lock\;
                if \$v5730\(0) = '1' then
                  state_var5920 := Q_WAIT5729;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18788\(48 to 63), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5728;
                end if;
              when Q_WAIT5732 =>
                \$v5733\ := \$code_lock\;
                if \$v5733\(0) = '1' then
                  state_var5920 := Q_WAIT5732;
                else
                  acquire(\$code_lock\);
                  \$code_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                  \$18788\(0 to 15), X"000" & X"2"), \$19265_ofs\)));
                  state_var5920 := PAUSE_GET5731;
                end if;
              when Q_WAIT5735 =>
                \$v5736\ := \$ram_lock\;
                if \$v5736\(0) = '1' then
                  state_var5920 := Q_WAIT5735;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18788\(16 to 46),16)));
                  state_var5920 := PAUSE_GET5734;
                end if;
              when Q_WAIT5739 =>
                \$v5740\ := \$ram_lock\;
                if \$v5740\(0) = '1' then
                  state_var5920 := Q_WAIT5739;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          work.Int.add(
                                                          \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(work.Int.add(work.Int.add(
                                                            \$18788\(0 to 15), X"000" & X"1"), eclat_resize(\$19215_argument1\,16)),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5738;
                end if;
              when Q_WAIT5742 =>
                \$v5743\ := \$ram_lock\;
                if \$v5743\(0) = '1' then
                  state_var5920 := Q_WAIT5742;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$18788\(104 to 119),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5741;
                end if;
              when Q_WAIT5745 =>
                \$v5746\ := \$ram_lock\;
                if \$v5746\(0) = '1' then
                  state_var5920 := Q_WAIT5745;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$18788\(48 to 63), X"000" & X"1")));
                  \$ram_write\ <= \$18788\(64 to 95); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5744;
                end if;
              when Q_WAIT5748 =>
                \$v5749\ := \$ram_lock\;
                if \$v5749\(0) = '1' then
                  state_var5920 := Q_WAIT5748;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= eclat_resize(\$18788\(96 to 103),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5747;
                end if;
              when Q_WAIT5751 =>
                \$v5752\ := \$ram_lock\;
                if \$v5752\(0) = '1' then
                  state_var5920 := Q_WAIT5751;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19273\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5750;
                end if;
              when Q_WAIT5755 =>
                \$v5756\ := \$ram_lock\;
                if \$v5756\(0) = '1' then
                  state_var5920 := Q_WAIT5755;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(64 to 95); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5754;
                end if;
              when Q_WAIT5758 =>
                \$v5759\ := \$ram_lock\;
                if \$v5759\(0) = '1' then
                  state_var5920 := Q_WAIT5758;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19281\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5757;
                end if;
              when Q_WAIT5762 =>
                \$v5763\ := \$ram_lock\;
                if \$v5763\(0) = '1' then
                  state_var5920 := Q_WAIT5762;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.sub(
                                                          \$18788\(48 to 63), X"000" & X"1")));
                  \$ram_write\ <= \$18788\(64 to 95); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5761;
                end if;
              when Q_WAIT5765 =>
                \$v5766\ := \$ram_lock\;
                if \$v5766\(0) = '1' then
                  state_var5920 := Q_WAIT5765;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18788\(48 to 63), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5764;
                end if;
              when Q_WAIT5768 =>
                \$v5769\ := \$ram_lock\;
                if \$v5769\(0) = '1' then
                  state_var5920 := Q_WAIT5768;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19290\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5767;
                end if;
              when Q_WAIT5772 =>
                \$v5773\ := \$ram_lock\;
                if \$v5773\(0) = '1' then
                  state_var5920 := Q_WAIT5772;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.sub(
                                                          work.Int.sub(
                                                          \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= \$18788\(64 to 95); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5771;
                end if;
              when Q_WAIT5775 =>
                \$v5776\ := \$ram_lock\;
                if \$v5776\(0) = '1' then
                  state_var5920 := Q_WAIT5775;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5774;
                end if;
              when Q_WAIT5778 =>
                \$v5779\ := \$ram_lock\;
                if \$v5779\(0) = '1' then
                  state_var5920 := Q_WAIT5778;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18788\(48 to 63), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5777;
                end if;
              when Q_WAIT5781 =>
                \$v5782\ := \$ram_lock\;
                if \$v5782\(0) = '1' then
                  state_var5920 := Q_WAIT5781;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19300\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5780;
                end if;
              when Q_WAIT5785 =>
                \$v5786\ := \$ram_lock\;
                if \$v5786\(0) = '1' then
                  state_var5920 := Q_WAIT5785;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.sub(
                                                          work.Int.sub(
                                                          work.Int.sub(
                                                          \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= \$18788\(64 to 95); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5784;
                end if;
              when Q_WAIT5788 =>
                \$v5789\ := \$ram_lock\;
                if \$v5789\(0) = '1' then
                  state_var5920 := Q_WAIT5788;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5787;
                end if;
              when Q_WAIT5791 =>
                \$v5792\ := \$ram_lock\;
                if \$v5792\(0) = '1' then
                  state_var5920 := Q_WAIT5791;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5790;
                end if;
              when Q_WAIT5794 =>
                \$v5795\ := \$ram_lock\;
                if \$v5795\(0) = '1' then
                  state_var5920 := Q_WAIT5794;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18788\(48 to 63), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5793;
                end if;
              when Q_WAIT5797 =>
                \$v5798\ := \$ram_lock\;
                if \$v5798\(0) = '1' then
                  state_var5920 := Q_WAIT5797;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19311\(80 to 95), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5796;
                end if;
              when Q_WAIT5801 =>
                \$v5802\ := \$ram_lock\;
                if \$v5802\(0) = '1' then
                  state_var5920 := Q_WAIT5801;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.sub(
                                                          work.Int.sub(
                                                          work.Int.sub(
                                                          work.Int.sub(
                                                          \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= \$18788\(64 to 95); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5800;
                end if;
              when Q_WAIT5804 =>
                \$v5805\ := \$ram_lock\;
                if \$v5805\(0) = '1' then
                  state_var5920 := Q_WAIT5804;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5803;
                end if;
              when Q_WAIT5807 =>
                \$v5808\ := \$ram_lock\;
                if \$v5808\(0) = '1' then
                  state_var5920 := Q_WAIT5807;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5806;
                end if;
              when Q_WAIT5810 =>
                \$v5811\ := \$ram_lock\;
                if \$v5811\(0) = '1' then
                  state_var5920 := Q_WAIT5810;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$18788\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5809;
                end if;
              when Q_WAIT5813 =>
                \$v5814\ := \$ram_lock\;
                if \$v5814\(0) = '1' then
                  state_var5920 := Q_WAIT5813;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$18788\(48 to 63), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5812;
                end if;
              when Q_WAIT5816 =>
                \$v5817\ := \$ram_lock\;
                if \$v5817\(0) = '1' then
                  state_var5920 := Q_WAIT5816;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5815;
                end if;
              when Q_WAIT5819 =>
                \$v5820\ := \$ram_lock\;
                if \$v5820\(0) = '1' then
                  state_var5920 := Q_WAIT5819;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$18788\(16 to 46),16), X"000" & X"0"), X"000" & X"1")));
                  \$ram_write\ <= work.Int.add(\$19324_f0\(0 to 30), \$19215_argument1\) & eclat_true; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5818;
                end if;
              when Q_WAIT5822 =>
                \$v5823\ := \$ram_lock\;
                if \$v5823\(0) = '1' then
                  state_var5920 := Q_WAIT5822;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18788\(16 to 46),16), X"000" & X"0"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5821;
                end if;
              when Q_WAIT5827 =>
                \$v5828\ := \$ram_lock\;
                if \$v5828\(0) = '1' then
                  state_var5920 := Q_WAIT5827;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$18788\(16 to 46),16), X"000" & X"0"), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5826;
                end if;
              when Q_WAIT5830 =>
                \$v5831\ := \$ram_lock\;
                if \$v5831\(0) = '1' then
                  state_var5920 := Q_WAIT5830;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$19347_fill6534389_arg\(48 to 78),16), \$19347_fill6534389_arg\(0 to 15)), X"000" & X"1")));
                  \$ram_write\ <= \$19350_v\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5829;
                end if;
              when Q_WAIT5833 =>
                \$v5834\ := \$ram_lock\;
                if \$v5834\(0) = '1' then
                  state_var5920 := Q_WAIT5833;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19347_fill6534389_arg\(16 to 31), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5832;
                end if;
              when Q_WAIT5837 =>
                \$v5838\ := \$ram_lock\;
                if \$v5838\(0) = '1' then
                  state_var5920 := Q_WAIT5837;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$19344\(64 to 94),16), X"000" & X"0"), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(work.Int.add(work.Int.add(
                                                            \$18788\(0 to 15), X"000" & X"2"), eclat_resize(\$19340_argument2\,16)),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5836;
                end if;
              when Q_WAIT5840 =>
                \$v5841\ := \$ram_lock\;
                if \$v5841\(0) = '1' then
                  state_var5920 := Q_WAIT5840;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5839;
                end if;
              when Q_WAIT5844 =>
                \$v5845\ := \$ram_lock\;
                if \$v5845\(0) = '1' then
                  state_var5920 := Q_WAIT5844;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$19353\(0 to 30),16), eclat_resize(\$19340_argument2\,16)), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5843;
                end if;
              when Q_WAIT5847 =>
                \$v5848\ := \$ram_lock\;
                if \$v5848\(0) = '1' then
                  state_var5920 := Q_WAIT5847;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(X"3e80", eclat_resize(\$19215_argument1\,16))));
                  state_var5920 := PAUSE_GET5846;
                end if;
              when Q_WAIT5850 =>
                \$v5851\ := \$ram_lock\;
                if \$v5851\(0) = '1' then
                  state_var5920 := Q_WAIT5850;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$19356\(0 to 30),16), eclat_resize(\$19340_argument2\,16)), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5849;
                end if;
              when Q_WAIT5853 =>
                \$v5854\ := \$ram_lock\;
                if \$v5854\(0) = '1' then
                  state_var5920 := Q_WAIT5853;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(X"3e80", eclat_resize(\$19215_argument1\,16))));
                  state_var5920 := PAUSE_GET5852;
                end if;
              when Q_WAIT5856 =>
                \$v5857\ := \$ram_lock\;
                if \$v5857\(0) = '1' then
                  state_var5920 := Q_WAIT5856;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5855;
                end if;
              when Q_WAIT5859 =>
                \$v5860\ := \$ram_lock\;
                if \$v5860\(0) = '1' then
                  state_var5920 := Q_WAIT5859;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$19361_fill6544390_arg\(48 to 78),16), \$19361_fill6544390_arg\(0 to 15)), X"000" & X"1")));
                  \$ram_write\ <= \$19364_v\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5858;
                end if;
              when Q_WAIT5862 =>
                \$v5863\ := \$ram_lock\;
                if \$v5863\(0) = '1' then
                  state_var5920 := Q_WAIT5862;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19361_fill6544390_arg\(16 to 31), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5861;
                end if;
              when Q_WAIT5866 =>
                \$v5867\ := \$ram_lock\;
                if \$v5867\(0) = '1' then
                  state_var5920 := Q_WAIT5866;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$19358\(64 to 94),16), X"000" & X"0"), X"000" & X"1")));
                  \$ram_write\ <= \$19358\(0 to 31); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5865;
                end if;
              when Q_WAIT5875 =>
                \$v5876\ := \$ram_lock\;
                if \$v5876\(0) = '1' then
                  state_var5920 := Q_WAIT5875;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$19416_w36574398_arg\(16 to 31)));
                  \$ram_write\ <= eclat_resize(work.Int.add(eclat_resize(\$19416_w36574398_arg\(48 to 78),16), 
                                                            work.Int.mul(
                                                            X"000" & X"2", \$19416_w36574398_arg\(0 to 15))),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5874;
                end if;
              when Q_WAIT5879 =>
                \$v5880\ := \$ram_lock\;
                if \$v5880\(0) = '1' then
                  state_var5920 := Q_WAIT5879;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$19412_sp\));
                  \$ram_write\ <= \$19410\(64 to 95); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5878;
                end if;
              when Q_WAIT5882 =>
                \$v5883\ := \$ram_lock\;
                if \$v5883\(0) = '1' then
                  state_var5920 := Q_WAIT5882;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$19420_w06554397_arg\(64 to 94),16), 
                                                          work.Int.sub(
                                                          work.Int.add(
                                                          \$19420_w06554397_arg\(0 to 15), 
                                                          work.Int.mul(
                                                          X"000" & X"2", \$19420_w06554397_arg\(32 to 47))), X"000" & X"1")), X"000" & X"1")));
                  \$ram_write\ <= \$19423_v\; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5881;
                end if;
              when Q_WAIT5885 =>
                \$v5886\ := \$ram_lock\;
                if \$v5886\(0) = '1' then
                  state_var5920 := Q_WAIT5885;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$19420_w06554397_arg\(16 to 31), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5884;
                end if;
              when Q_WAIT5889 =>
                \$v5890\ := \$ram_lock\;
                if \$v5890\(0) = '1' then
                  state_var5920 := Q_WAIT5889;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$19410\(64 to 94),16), X"000" & X"0"), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(work.Int.add(work.Int.add(
                                                            \$18788\(0 to 15), X"000" & X"3"), eclat_resize(\$19408_argument3\,16)),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5888;
                end if;
              when Q_WAIT5892 =>
                \$v5893\ := \$ram_lock\;
                if \$v5893\(0) = '1' then
                  state_var5920 := Q_WAIT5892;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$18788\(48 to 63)));
                  \$ram_write\ <= \$18788\(16 to 47); \$ram_write_request\ <= '1';
                  state_var5920 := PAUSE_SET5891;
                end if;
              when Q_WAIT5896 =>
                \$v5897\ := \$code_lock\;
                if \$v5897\(0) = '1' then
                  state_var5920 := Q_WAIT5896;
                else
                  acquire(\$code_lock\);
                  \$code_ptr\ <= to_integer(unsigned(\$18788\(0 to 15)));
                  state_var5920 := PAUSE_GET5895;
                end if;
              when Q_WAIT5900 =>
                \$v5901\ := \$code_lock\;
                if \$v5901\(0) = '1' then
                  state_var5920 := Q_WAIT5900;
                else
                  acquire(\$code_lock\);
                  \$code_ptr\ <= to_integer(unsigned(work.Int.add(\$18788\(0 to 15), X"000" & X"3")));
                  state_var5920 := PAUSE_GET5899;
                end if;
              when Q_WAIT5904 =>
                \$v5905\ := \$code_lock\;
                if \$v5905\(0) = '1' then
                  state_var5920 := Q_WAIT5904;
                else
                  acquire(\$code_lock\);
                  \$code_ptr\ <= to_integer(unsigned(work.Int.add(\$18788\(0 to 15), X"000" & X"2")));
                  state_var5920 := PAUSE_GET5903;
                end if;
              when Q_WAIT5908 =>
                \$v5909\ := \$code_lock\;
                if \$v5909\(0) = '1' then
                  state_var5920 := Q_WAIT5908;
                else
                  acquire(\$code_lock\);
                  \$code_ptr\ <= to_integer(unsigned(work.Int.add(\$18788\(0 to 15), X"000" & X"1")));
                  state_var5920 := PAUSE_GET5907;
                end if;
              when Q_WAIT5912 =>
                \$v5913\ := \$code_lock\;
                if \$v5913\(0) = '1' then
                  state_var5920 := Q_WAIT5912;
                else
                  acquire(\$code_lock\);
                  \$code_ptr\ <= to_integer(unsigned(\$18788\(0 to 15)));
                  state_var5920 := PAUSE_GET5911;
                end if;
              when IDLE4930 =>
                rdy4929 := eclat_false;
                \$18800\ := work.Print.print_string(clk,of_string("pc:"));
                \$18801\ := work.Int.print(clk,\$18788\(0 to 15));
                \$18802\ := work.Print.print_string(clk,of_string("|acc:"));
                \$18803\ := work.Int.print(clk,\$18788\(16 to 46));
                \$18804\ := work.Print.print_string(clk,of_string("<"));
                \$v5915\ := ""&\$18788\(47);
                if \$v5915\(0) = '1' then
                  \$18805\ := work.Print.print_string(clk,of_string("int"));
                  \$18806\ := work.Print.print_string(clk,of_string(">"));
                  \$18807\ := work.Print.print_string(clk,of_string("|sp:"));
                  \$18808\ := work.Int.print(clk,\$18788\(48 to 63));
                  \$18809\ := work.Print.print_string(clk,of_string("|env:"));
                  \$18810\ := work.Int.print(clk,\$18788\(64 to 94));
                  \$18811\ := work.Print.print_string(clk,of_string("<"));
                  \$v5914\ := ""&\$18788\(95);
                  if \$v5914\(0) = '1' then
                    \$18812\ := work.Print.print_string(clk,of_string("int"));
                    \$18813\ := work.Print.print_string(clk,of_string(">"));
                    \$18814\ := work.Print.print_newline(clk,eclat_unit);
                    \$18815\ := work.Assertion.ok(work.Int.lt(\$18788\(0 to 15), std_logic_vector(to_unsigned(code'length,16))));
                    \$v5913\ := \$code_lock\;
                    if \$v5913\(0) = '1' then
                      state_var5920 := Q_WAIT5912;
                    else
                      acquire(\$code_lock\);
                      \$code_ptr\ <= to_integer(unsigned(\$18788\(0 to 15)));
                      state_var5920 := PAUSE_GET5911;
                    end if;
                  else
                    \$18812\ := work.Print.print_string(clk,of_string("ptr"));
                    \$18813\ := work.Print.print_string(clk,of_string(">"));
                    \$18814\ := work.Print.print_newline(clk,eclat_unit);
                    \$18815\ := work.Assertion.ok(work.Int.lt(\$18788\(0 to 15), std_logic_vector(to_unsigned(code'length,16))));
                    \$v5913\ := \$code_lock\;
                    if \$v5913\(0) = '1' then
                      state_var5920 := Q_WAIT5912;
                    else
                      acquire(\$code_lock\);
                      \$code_ptr\ <= to_integer(unsigned(\$18788\(0 to 15)));
                      state_var5920 := PAUSE_GET5911;
                    end if;
                  end if;
                else
                  \$18805\ := work.Print.print_string(clk,of_string("ptr"));
                  \$18806\ := work.Print.print_string(clk,of_string(">"));
                  \$18807\ := work.Print.print_string(clk,of_string("|sp:"));
                  \$18808\ := work.Int.print(clk,\$18788\(48 to 63));
                  \$18809\ := work.Print.print_string(clk,of_string("|env:"));
                  \$18810\ := work.Int.print(clk,\$18788\(64 to 94));
                  \$18811\ := work.Print.print_string(clk,of_string("<"));
                  \$v5914\ := ""&\$18788\(95);
                  if \$v5914\(0) = '1' then
                    \$18812\ := work.Print.print_string(clk,of_string("int"));
                    \$18813\ := work.Print.print_string(clk,of_string(">"));
                    \$18814\ := work.Print.print_newline(clk,eclat_unit);
                    \$18815\ := work.Assertion.ok(work.Int.lt(\$18788\(0 to 15), std_logic_vector(to_unsigned(code'length,16))));
                    \$v5913\ := \$code_lock\;
                    if \$v5913\(0) = '1' then
                      state_var5920 := Q_WAIT5912;
                    else
                      acquire(\$code_lock\);
                      \$code_ptr\ <= to_integer(unsigned(\$18788\(0 to 15)));
                      state_var5920 := PAUSE_GET5911;
                    end if;
                  else
                    \$18812\ := work.Print.print_string(clk,of_string("ptr"));
                    \$18813\ := work.Print.print_string(clk,of_string(">"));
                    \$18814\ := work.Print.print_newline(clk,eclat_unit);
                    \$18815\ := work.Assertion.ok(work.Int.lt(\$18788\(0 to 15), std_logic_vector(to_unsigned(code'length,16))));
                    \$v5913\ := \$code_lock\;
                    if \$v5913\(0) = '1' then
                      state_var5920 := Q_WAIT5912;
                    else
                      acquire(\$code_lock\);
                      \$code_ptr\ <= to_integer(unsigned(\$18788\(0 to 15)));
                      state_var5920 := PAUSE_GET5911;
                    end if;
                  end if;
                end if;
              end case;
              
              if rdy4929(0) = '1' then
                
              else
                result4928 := \$18788\(0 to 121);
              end if;
              \$18789\ := result4928 & rdy4929;
              \$18788\ := \$18789\(0 to 121) & ""&\$18789\(122);
            end if;
            \$18787\ := \$18788\;
            \$18462\ := ""&\$18787\(120) & ""&\$18787\(122) & ""&\$18462\(2) & ""&\$18787\(121);
          end if;
          \$18443\ := \$18462\;
          \$v4571\ := ""&\$18443\(0);
          if \$v4571\(0) = '1' then
            \$18459\ := work.Print.print_string(clk,of_string("(cy="));
            \$18460\ := work.Int.print(clk,\$18442_cy\);
            \$18461\ := work.Print.print_string(clk,of_string(")"));
            \$18444\ := work.Print.print_newline(clk,eclat_unit);
            if \$v4337\(0) = '1' then
              
            else
              \$v4337\ := eclat_true;
              \$18458\ := eclat_false;
            end if;
            \$18458\ := eclat_if(""&\$18443\(0) & eclat_true & \$18458\);
            \$18445_x\ := \$18458\;
            if \$v4338\(0) = '1' then
              
            else
              \$v4338\ := eclat_true;
              \$18457\ := X"0000000" & X"0";
            end if;
            \$18457\ := eclat_if(work.Bool.lnot(\$18445_x\) & work.Int.add(
                                                              \$18457\, X"0000000" & X"1") & \$18457\);
            \$18446_dur\ := \$18457\;
            \$v4570\ := \$18445_x\;
            if \$v4570\(0) = '1' then
              \$18447\ := work.Int.print(clk,\$18446_dur\);
              \$v4569\ := \$18445_x\;
              if \$v4569\(0) = '1' then
                \$v4568\ := eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"3") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"2") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"1") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"0");
                case \$v4568\ is
                when "0000" =>
                  \$18451\ := "00000011";
                when "0001" =>
                  \$18451\ := "10011111";
                when "0010" =>
                  \$18451\ := "00100101";
                when "0011" =>
                  \$18451\ := "00001101";
                when "0100" =>
                  \$18451\ := "10011001";
                when "0101" =>
                  \$18451\ := "01001001";
                when "0110" =>
                  \$18451\ := "01000001";
                when "0111" =>
                  \$18451\ := "00011111";
                when "1000" =>
                  \$18451\ := "00000001";
                when "1001" =>
                  \$18451\ := "00001001";
                when "1010" =>
                  \$18451\ := "00010001";
                when "1011" =>
                  \$18451\ := "11000001";
                when "1100" =>
                  \$18451\ := "01100011";
                when "1101" =>
                  \$18451\ := "10000101";
                when "1110" =>
                  \$18451\ := "01100001";
                when "1111" =>
                  \$18451\ := "01110001";
                when others =>
                  \$18451\ := "11100011";
                end case;
                \$v4567\ := eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"7") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"6") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"5") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"4");
                case \$v4567\ is
                when "0000" =>
                  \$18452\ := "00000011";
                when "0001" =>
                  \$18452\ := "10011111";
                when "0010" =>
                  \$18452\ := "00100101";
                when "0011" =>
                  \$18452\ := "00001101";
                when "0100" =>
                  \$18452\ := "10011001";
                when "0101" =>
                  \$18452\ := "01001001";
                when "0110" =>
                  \$18452\ := "01000001";
                when "0111" =>
                  \$18452\ := "00011111";
                when "1000" =>
                  \$18452\ := "00000001";
                when "1001" =>
                  \$18452\ := "00001001";
                when "1010" =>
                  \$18452\ := "00010001";
                when "1011" =>
                  \$18452\ := "11000001";
                when "1100" =>
                  \$18452\ := "01100011";
                when "1101" =>
                  \$18452\ := "10000101";
                when "1110" =>
                  \$18452\ := "01100001";
                when "1111" =>
                  \$18452\ := "01110001";
                when others =>
                  \$18452\ := "11100011";
                end case;
                \$v4566\ := eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"b") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"a") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"9") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"8");
                case \$v4566\ is
                when "0000" =>
                  \$18453\ := "00000011";
                when "0001" =>
                  \$18453\ := "10011111";
                when "0010" =>
                  \$18453\ := "00100101";
                when "0011" =>
                  \$18453\ := "00001101";
                when "0100" =>
                  \$18453\ := "10011001";
                when "0101" =>
                  \$18453\ := "01001001";
                when "0110" =>
                  \$18453\ := "01000001";
                when "0111" =>
                  \$18453\ := "00011111";
                when "1000" =>
                  \$18453\ := "00000001";
                when "1001" =>
                  \$18453\ := "00001001";
                when "1010" =>
                  \$18453\ := "00010001";
                when "1011" =>
                  \$18453\ := "11000001";
                when "1100" =>
                  \$18453\ := "01100011";
                when "1101" =>
                  \$18453\ := "10000101";
                when "1110" =>
                  \$18453\ := "01100001";
                when "1111" =>
                  \$18453\ := "01110001";
                when others =>
                  \$18453\ := "11100011";
                end case;
                \$v4565\ := eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"f") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"e") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"d") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"c");
                case \$v4565\ is
                when "0000" =>
                  \$18454\ := "00000011";
                when "0001" =>
                  \$18454\ := "10011111";
                when "0010" =>
                  \$18454\ := "00100101";
                when "0011" =>
                  \$18454\ := "00001101";
                when "0100" =>
                  \$18454\ := "10011001";
                when "0101" =>
                  \$18454\ := "01001001";
                when "0110" =>
                  \$18454\ := "01000001";
                when "0111" =>
                  \$18454\ := "00011111";
                when "1000" =>
                  \$18454\ := "00000001";
                when "1001" =>
                  \$18454\ := "00001001";
                when "1010" =>
                  \$18454\ := "00010001";
                when "1011" =>
                  \$18454\ := "11000001";
                when "1100" =>
                  \$18454\ := "01100011";
                when "1101" =>
                  \$18454\ := "10000101";
                when "1110" =>
                  \$18454\ := "01100001";
                when "1111" =>
                  \$18454\ := "01110001";
                when others =>
                  \$18454\ := "11100011";
                end case;
                \$v4564\ := eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"13") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"12") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"11") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"10");
                case \$v4564\ is
                when "0000" =>
                  \$18455\ := "00000011";
                when "0001" =>
                  \$18455\ := "10011111";
                when "0010" =>
                  \$18455\ := "00100101";
                when "0011" =>
                  \$18455\ := "00001101";
                when "0100" =>
                  \$18455\ := "10011001";
                when "0101" =>
                  \$18455\ := "01001001";
                when "0110" =>
                  \$18455\ := "01000001";
                when "0111" =>
                  \$18455\ := "00011111";
                when "1000" =>
                  \$18455\ := "00000001";
                when "1001" =>
                  \$18455\ := "00001001";
                when "1010" =>
                  \$18455\ := "00010001";
                when "1011" =>
                  \$18455\ := "11000001";
                when "1100" =>
                  \$18455\ := "01100011";
                when "1101" =>
                  \$18455\ := "10000101";
                when "1110" =>
                  \$18455\ := "01100001";
                when "1111" =>
                  \$18455\ := "01110001";
                when others =>
                  \$18455\ := "11100011";
                end case;
                \$v4563\ := eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"17") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"16") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"15") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"14");
                case \$v4563\ is
                when "0000" =>
                  \$18456\ := "00000011";
                when "0001" =>
                  \$18456\ := "10011111";
                when "0010" =>
                  \$18456\ := "00100101";
                when "0011" =>
                  \$18456\ := "00001101";
                when "0100" =>
                  \$18456\ := "10011001";
                when "0101" =>
                  \$18456\ := "01001001";
                when "0110" =>
                  \$18456\ := "01000001";
                when "0111" =>
                  \$18456\ := "00011111";
                when "1000" =>
                  \$18456\ := "00000001";
                when "1001" =>
                  \$18456\ := "00001001";
                when "1010" =>
                  \$18456\ := "00010001";
                when "1011" =>
                  \$18456\ := "11000001";
                when "1100" =>
                  \$18456\ := "01100011";
                when "1101" =>
                  \$18456\ := "10000101";
                when "1110" =>
                  \$18456\ := "01100001";
                when "1111" =>
                  \$18456\ := "01110001";
                when others =>
                  \$18456\ := "11100011";
                end case;
                \$18448_dis\ := \$18451\ & \$18452\ & \$18453\ & \$18454\ & \$18455\ & \$18456\;
              else
                \$18448_dis\ := "00000011" & "00000011" & "00000011" & "00000011" & "00000011" & "00000011";
              end if;
              if \$v4339\(0) = '1' then
                
              else
                \$v4339\ := eclat_true;
                \$18450\ := X"0000000" & X"0";
              end if;
              \$18450\ := eclat_if(work.Int.eq(\$18450\, work.Int.add(
                                                         X"00" & X"989680", X"00" & X"989680")) & X"0000000" & X"0" & 
                          work.Int.add(\$18450\, X"0000000" & X"1"));
              \$18449\ := \$18450\;
              result4399 := ""&\$18443\(0) & work.Bool.lnot(""&\$18443\(1)) & 
              work.Int.gt(\$18449\, X"00" & X"989680") & ""&\$18443\(3) & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & \$18448_dis\;
              rdy4400 := eclat_true;
              state := IDLE4401;
            else
              \$18447\ := eclat_unit;
              \$v4569\ := \$18445_x\;
              if \$v4569\(0) = '1' then
                \$v4568\ := eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"3") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"2") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"1") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"0");
                case \$v4568\ is
                when "0000" =>
                  \$18451\ := "00000011";
                when "0001" =>
                  \$18451\ := "10011111";
                when "0010" =>
                  \$18451\ := "00100101";
                when "0011" =>
                  \$18451\ := "00001101";
                when "0100" =>
                  \$18451\ := "10011001";
                when "0101" =>
                  \$18451\ := "01001001";
                when "0110" =>
                  \$18451\ := "01000001";
                when "0111" =>
                  \$18451\ := "00011111";
                when "1000" =>
                  \$18451\ := "00000001";
                when "1001" =>
                  \$18451\ := "00001001";
                when "1010" =>
                  \$18451\ := "00010001";
                when "1011" =>
                  \$18451\ := "11000001";
                when "1100" =>
                  \$18451\ := "01100011";
                when "1101" =>
                  \$18451\ := "10000101";
                when "1110" =>
                  \$18451\ := "01100001";
                when "1111" =>
                  \$18451\ := "01110001";
                when others =>
                  \$18451\ := "11100011";
                end case;
                \$v4567\ := eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"7") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"6") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"5") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"4");
                case \$v4567\ is
                when "0000" =>
                  \$18452\ := "00000011";
                when "0001" =>
                  \$18452\ := "10011111";
                when "0010" =>
                  \$18452\ := "00100101";
                when "0011" =>
                  \$18452\ := "00001101";
                when "0100" =>
                  \$18452\ := "10011001";
                when "0101" =>
                  \$18452\ := "01001001";
                when "0110" =>
                  \$18452\ := "01000001";
                when "0111" =>
                  \$18452\ := "00011111";
                when "1000" =>
                  \$18452\ := "00000001";
                when "1001" =>
                  \$18452\ := "00001001";
                when "1010" =>
                  \$18452\ := "00010001";
                when "1011" =>
                  \$18452\ := "11000001";
                when "1100" =>
                  \$18452\ := "01100011";
                when "1101" =>
                  \$18452\ := "10000101";
                when "1110" =>
                  \$18452\ := "01100001";
                when "1111" =>
                  \$18452\ := "01110001";
                when others =>
                  \$18452\ := "11100011";
                end case;
                \$v4566\ := eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"b") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"a") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"9") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"8");
                case \$v4566\ is
                when "0000" =>
                  \$18453\ := "00000011";
                when "0001" =>
                  \$18453\ := "10011111";
                when "0010" =>
                  \$18453\ := "00100101";
                when "0011" =>
                  \$18453\ := "00001101";
                when "0100" =>
                  \$18453\ := "10011001";
                when "0101" =>
                  \$18453\ := "01001001";
                when "0110" =>
                  \$18453\ := "01000001";
                when "0111" =>
                  \$18453\ := "00011111";
                when "1000" =>
                  \$18453\ := "00000001";
                when "1001" =>
                  \$18453\ := "00001001";
                when "1010" =>
                  \$18453\ := "00010001";
                when "1011" =>
                  \$18453\ := "11000001";
                when "1100" =>
                  \$18453\ := "01100011";
                when "1101" =>
                  \$18453\ := "10000101";
                when "1110" =>
                  \$18453\ := "01100001";
                when "1111" =>
                  \$18453\ := "01110001";
                when others =>
                  \$18453\ := "11100011";
                end case;
                \$v4565\ := eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"f") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"e") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"d") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"c");
                case \$v4565\ is
                when "0000" =>
                  \$18454\ := "00000011";
                when "0001" =>
                  \$18454\ := "10011111";
                when "0010" =>
                  \$18454\ := "00100101";
                when "0011" =>
                  \$18454\ := "00001101";
                when "0100" =>
                  \$18454\ := "10011001";
                when "0101" =>
                  \$18454\ := "01001001";
                when "0110" =>
                  \$18454\ := "01000001";
                when "0111" =>
                  \$18454\ := "00011111";
                when "1000" =>
                  \$18454\ := "00000001";
                when "1001" =>
                  \$18454\ := "00001001";
                when "1010" =>
                  \$18454\ := "00010001";
                when "1011" =>
                  \$18454\ := "11000001";
                when "1100" =>
                  \$18454\ := "01100011";
                when "1101" =>
                  \$18454\ := "10000101";
                when "1110" =>
                  \$18454\ := "01100001";
                when "1111" =>
                  \$18454\ := "01110001";
                when others =>
                  \$18454\ := "11100011";
                end case;
                \$v4564\ := eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"13") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"12") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"11") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"10");
                case \$v4564\ is
                when "0000" =>
                  \$18455\ := "00000011";
                when "0001" =>
                  \$18455\ := "10011111";
                when "0010" =>
                  \$18455\ := "00100101";
                when "0011" =>
                  \$18455\ := "00001101";
                when "0100" =>
                  \$18455\ := "10011001";
                when "0101" =>
                  \$18455\ := "01001001";
                when "0110" =>
                  \$18455\ := "01000001";
                when "0111" =>
                  \$18455\ := "00011111";
                when "1000" =>
                  \$18455\ := "00000001";
                when "1001" =>
                  \$18455\ := "00001001";
                when "1010" =>
                  \$18455\ := "00010001";
                when "1011" =>
                  \$18455\ := "11000001";
                when "1100" =>
                  \$18455\ := "01100011";
                when "1101" =>
                  \$18455\ := "10000101";
                when "1110" =>
                  \$18455\ := "01100001";
                when "1111" =>
                  \$18455\ := "01110001";
                when others =>
                  \$18455\ := "11100011";
                end case;
                \$v4563\ := eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"17") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"16") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"15") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"14");
                case \$v4563\ is
                when "0000" =>
                  \$18456\ := "00000011";
                when "0001" =>
                  \$18456\ := "10011111";
                when "0010" =>
                  \$18456\ := "00100101";
                when "0011" =>
                  \$18456\ := "00001101";
                when "0100" =>
                  \$18456\ := "10011001";
                when "0101" =>
                  \$18456\ := "01001001";
                when "0110" =>
                  \$18456\ := "01000001";
                when "0111" =>
                  \$18456\ := "00011111";
                when "1000" =>
                  \$18456\ := "00000001";
                when "1001" =>
                  \$18456\ := "00001001";
                when "1010" =>
                  \$18456\ := "00010001";
                when "1011" =>
                  \$18456\ := "11000001";
                when "1100" =>
                  \$18456\ := "01100011";
                when "1101" =>
                  \$18456\ := "10000101";
                when "1110" =>
                  \$18456\ := "01100001";
                when "1111" =>
                  \$18456\ := "01110001";
                when others =>
                  \$18456\ := "11100011";
                end case;
                \$18448_dis\ := \$18451\ & \$18452\ & \$18453\ & \$18454\ & \$18455\ & \$18456\;
              else
                \$18448_dis\ := "00000011" & "00000011" & "00000011" & "00000011" & "00000011" & "00000011";
              end if;
              if \$v4339\(0) = '1' then
                
              else
                \$v4339\ := eclat_true;
                \$18450\ := X"0000000" & X"0";
              end if;
              \$18450\ := eclat_if(work.Int.eq(\$18450\, work.Int.add(
                                                         X"00" & X"989680", X"00" & X"989680")) & X"0000000" & X"0" & 
                          work.Int.add(\$18450\, X"0000000" & X"1"));
              \$18449\ := \$18450\;
              result4399 := ""&\$18443\(0) & work.Bool.lnot(""&\$18443\(1)) & 
              work.Int.gt(\$18449\, X"00" & X"989680") & ""&\$18443\(3) & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & \$18448_dis\;
              rdy4400 := eclat_true;
              state := IDLE4401;
            end if;
          else
            \$18444\ := eclat_unit;
            if \$v4337\(0) = '1' then
              
            else
              \$v4337\ := eclat_true;
              \$18458\ := eclat_false;
            end if;
            \$18458\ := eclat_if(""&\$18443\(0) & eclat_true & \$18458\);
            \$18445_x\ := \$18458\;
            if \$v4338\(0) = '1' then
              
            else
              \$v4338\ := eclat_true;
              \$18457\ := X"0000000" & X"0";
            end if;
            \$18457\ := eclat_if(work.Bool.lnot(\$18445_x\) & work.Int.add(
                                                              \$18457\, X"0000000" & X"1") & \$18457\);
            \$18446_dur\ := \$18457\;
            \$v4570\ := \$18445_x\;
            if \$v4570\(0) = '1' then
              \$18447\ := work.Int.print(clk,\$18446_dur\);
              \$v4569\ := \$18445_x\;
              if \$v4569\(0) = '1' then
                \$v4568\ := eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"3") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"2") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"1") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"0");
                case \$v4568\ is
                when "0000" =>
                  \$18451\ := "00000011";
                when "0001" =>
                  \$18451\ := "10011111";
                when "0010" =>
                  \$18451\ := "00100101";
                when "0011" =>
                  \$18451\ := "00001101";
                when "0100" =>
                  \$18451\ := "10011001";
                when "0101" =>
                  \$18451\ := "01001001";
                when "0110" =>
                  \$18451\ := "01000001";
                when "0111" =>
                  \$18451\ := "00011111";
                when "1000" =>
                  \$18451\ := "00000001";
                when "1001" =>
                  \$18451\ := "00001001";
                when "1010" =>
                  \$18451\ := "00010001";
                when "1011" =>
                  \$18451\ := "11000001";
                when "1100" =>
                  \$18451\ := "01100011";
                when "1101" =>
                  \$18451\ := "10000101";
                when "1110" =>
                  \$18451\ := "01100001";
                when "1111" =>
                  \$18451\ := "01110001";
                when others =>
                  \$18451\ := "11100011";
                end case;
                \$v4567\ := eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"7") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"6") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"5") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"4");
                case \$v4567\ is
                when "0000" =>
                  \$18452\ := "00000011";
                when "0001" =>
                  \$18452\ := "10011111";
                when "0010" =>
                  \$18452\ := "00100101";
                when "0011" =>
                  \$18452\ := "00001101";
                when "0100" =>
                  \$18452\ := "10011001";
                when "0101" =>
                  \$18452\ := "01001001";
                when "0110" =>
                  \$18452\ := "01000001";
                when "0111" =>
                  \$18452\ := "00011111";
                when "1000" =>
                  \$18452\ := "00000001";
                when "1001" =>
                  \$18452\ := "00001001";
                when "1010" =>
                  \$18452\ := "00010001";
                when "1011" =>
                  \$18452\ := "11000001";
                when "1100" =>
                  \$18452\ := "01100011";
                when "1101" =>
                  \$18452\ := "10000101";
                when "1110" =>
                  \$18452\ := "01100001";
                when "1111" =>
                  \$18452\ := "01110001";
                when others =>
                  \$18452\ := "11100011";
                end case;
                \$v4566\ := eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"b") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"a") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"9") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"8");
                case \$v4566\ is
                when "0000" =>
                  \$18453\ := "00000011";
                when "0001" =>
                  \$18453\ := "10011111";
                when "0010" =>
                  \$18453\ := "00100101";
                when "0011" =>
                  \$18453\ := "00001101";
                when "0100" =>
                  \$18453\ := "10011001";
                when "0101" =>
                  \$18453\ := "01001001";
                when "0110" =>
                  \$18453\ := "01000001";
                when "0111" =>
                  \$18453\ := "00011111";
                when "1000" =>
                  \$18453\ := "00000001";
                when "1001" =>
                  \$18453\ := "00001001";
                when "1010" =>
                  \$18453\ := "00010001";
                when "1011" =>
                  \$18453\ := "11000001";
                when "1100" =>
                  \$18453\ := "01100011";
                when "1101" =>
                  \$18453\ := "10000101";
                when "1110" =>
                  \$18453\ := "01100001";
                when "1111" =>
                  \$18453\ := "01110001";
                when others =>
                  \$18453\ := "11100011";
                end case;
                \$v4565\ := eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"f") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"e") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"d") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"c");
                case \$v4565\ is
                when "0000" =>
                  \$18454\ := "00000011";
                when "0001" =>
                  \$18454\ := "10011111";
                when "0010" =>
                  \$18454\ := "00100101";
                when "0011" =>
                  \$18454\ := "00001101";
                when "0100" =>
                  \$18454\ := "10011001";
                when "0101" =>
                  \$18454\ := "01001001";
                when "0110" =>
                  \$18454\ := "01000001";
                when "0111" =>
                  \$18454\ := "00011111";
                when "1000" =>
                  \$18454\ := "00000001";
                when "1001" =>
                  \$18454\ := "00001001";
                when "1010" =>
                  \$18454\ := "00010001";
                when "1011" =>
                  \$18454\ := "11000001";
                when "1100" =>
                  \$18454\ := "01100011";
                when "1101" =>
                  \$18454\ := "10000101";
                when "1110" =>
                  \$18454\ := "01100001";
                when "1111" =>
                  \$18454\ := "01110001";
                when others =>
                  \$18454\ := "11100011";
                end case;
                \$v4564\ := eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"13") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"12") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"11") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"10");
                case \$v4564\ is
                when "0000" =>
                  \$18455\ := "00000011";
                when "0001" =>
                  \$18455\ := "10011111";
                when "0010" =>
                  \$18455\ := "00100101";
                when "0011" =>
                  \$18455\ := "00001101";
                when "0100" =>
                  \$18455\ := "10011001";
                when "0101" =>
                  \$18455\ := "01001001";
                when "0110" =>
                  \$18455\ := "01000001";
                when "0111" =>
                  \$18455\ := "00011111";
                when "1000" =>
                  \$18455\ := "00000001";
                when "1001" =>
                  \$18455\ := "00001001";
                when "1010" =>
                  \$18455\ := "00010001";
                when "1011" =>
                  \$18455\ := "11000001";
                when "1100" =>
                  \$18455\ := "01100011";
                when "1101" =>
                  \$18455\ := "10000101";
                when "1110" =>
                  \$18455\ := "01100001";
                when "1111" =>
                  \$18455\ := "01110001";
                when others =>
                  \$18455\ := "11100011";
                end case;
                \$v4563\ := eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"17") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"16") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"15") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"14");
                case \$v4563\ is
                when "0000" =>
                  \$18456\ := "00000011";
                when "0001" =>
                  \$18456\ := "10011111";
                when "0010" =>
                  \$18456\ := "00100101";
                when "0011" =>
                  \$18456\ := "00001101";
                when "0100" =>
                  \$18456\ := "10011001";
                when "0101" =>
                  \$18456\ := "01001001";
                when "0110" =>
                  \$18456\ := "01000001";
                when "0111" =>
                  \$18456\ := "00011111";
                when "1000" =>
                  \$18456\ := "00000001";
                when "1001" =>
                  \$18456\ := "00001001";
                when "1010" =>
                  \$18456\ := "00010001";
                when "1011" =>
                  \$18456\ := "11000001";
                when "1100" =>
                  \$18456\ := "01100011";
                when "1101" =>
                  \$18456\ := "10000101";
                when "1110" =>
                  \$18456\ := "01100001";
                when "1111" =>
                  \$18456\ := "01110001";
                when others =>
                  \$18456\ := "11100011";
                end case;
                \$18448_dis\ := \$18451\ & \$18452\ & \$18453\ & \$18454\ & \$18455\ & \$18456\;
              else
                \$18448_dis\ := "00000011" & "00000011" & "00000011" & "00000011" & "00000011" & "00000011";
              end if;
              if \$v4339\(0) = '1' then
                
              else
                \$v4339\ := eclat_true;
                \$18450\ := X"0000000" & X"0";
              end if;
              \$18450\ := eclat_if(work.Int.eq(\$18450\, work.Int.add(
                                                         X"00" & X"989680", X"00" & X"989680")) & X"0000000" & X"0" & 
                          work.Int.add(\$18450\, X"0000000" & X"1"));
              \$18449\ := \$18450\;
              result4399 := ""&\$18443\(0) & work.Bool.lnot(""&\$18443\(1)) & 
              work.Int.gt(\$18449\, X"00" & X"989680") & ""&\$18443\(3) & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & \$18448_dis\;
              rdy4400 := eclat_true;
              state := IDLE4401;
            else
              \$18447\ := eclat_unit;
              \$v4569\ := \$18445_x\;
              if \$v4569\(0) = '1' then
                \$v4568\ := eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"3") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"2") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"1") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"0");
                case \$v4568\ is
                when "0000" =>
                  \$18451\ := "00000011";
                when "0001" =>
                  \$18451\ := "10011111";
                when "0010" =>
                  \$18451\ := "00100101";
                when "0011" =>
                  \$18451\ := "00001101";
                when "0100" =>
                  \$18451\ := "10011001";
                when "0101" =>
                  \$18451\ := "01001001";
                when "0110" =>
                  \$18451\ := "01000001";
                when "0111" =>
                  \$18451\ := "00011111";
                when "1000" =>
                  \$18451\ := "00000001";
                when "1001" =>
                  \$18451\ := "00001001";
                when "1010" =>
                  \$18451\ := "00010001";
                when "1011" =>
                  \$18451\ := "11000001";
                when "1100" =>
                  \$18451\ := "01100011";
                when "1101" =>
                  \$18451\ := "10000101";
                when "1110" =>
                  \$18451\ := "01100001";
                when "1111" =>
                  \$18451\ := "01110001";
                when others =>
                  \$18451\ := "11100011";
                end case;
                \$v4567\ := eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"7") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"6") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"5") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"4");
                case \$v4567\ is
                when "0000" =>
                  \$18452\ := "00000011";
                when "0001" =>
                  \$18452\ := "10011111";
                when "0010" =>
                  \$18452\ := "00100101";
                when "0011" =>
                  \$18452\ := "00001101";
                when "0100" =>
                  \$18452\ := "10011001";
                when "0101" =>
                  \$18452\ := "01001001";
                when "0110" =>
                  \$18452\ := "01000001";
                when "0111" =>
                  \$18452\ := "00011111";
                when "1000" =>
                  \$18452\ := "00000001";
                when "1001" =>
                  \$18452\ := "00001001";
                when "1010" =>
                  \$18452\ := "00010001";
                when "1011" =>
                  \$18452\ := "11000001";
                when "1100" =>
                  \$18452\ := "01100011";
                when "1101" =>
                  \$18452\ := "10000101";
                when "1110" =>
                  \$18452\ := "01100001";
                when "1111" =>
                  \$18452\ := "01110001";
                when others =>
                  \$18452\ := "11100011";
                end case;
                \$v4566\ := eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"b") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"a") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"9") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"8");
                case \$v4566\ is
                when "0000" =>
                  \$18453\ := "00000011";
                when "0001" =>
                  \$18453\ := "10011111";
                when "0010" =>
                  \$18453\ := "00100101";
                when "0011" =>
                  \$18453\ := "00001101";
                when "0100" =>
                  \$18453\ := "10011001";
                when "0101" =>
                  \$18453\ := "01001001";
                when "0110" =>
                  \$18453\ := "01000001";
                when "0111" =>
                  \$18453\ := "00011111";
                when "1000" =>
                  \$18453\ := "00000001";
                when "1001" =>
                  \$18453\ := "00001001";
                when "1010" =>
                  \$18453\ := "00010001";
                when "1011" =>
                  \$18453\ := "11000001";
                when "1100" =>
                  \$18453\ := "01100011";
                when "1101" =>
                  \$18453\ := "10000101";
                when "1110" =>
                  \$18453\ := "01100001";
                when "1111" =>
                  \$18453\ := "01110001";
                when others =>
                  \$18453\ := "11100011";
                end case;
                \$v4565\ := eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"f") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"e") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"d") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"0000000" & X"c");
                case \$v4565\ is
                when "0000" =>
                  \$18454\ := "00000011";
                when "0001" =>
                  \$18454\ := "10011111";
                when "0010" =>
                  \$18454\ := "00100101";
                when "0011" =>
                  \$18454\ := "00001101";
                when "0100" =>
                  \$18454\ := "10011001";
                when "0101" =>
                  \$18454\ := "01001001";
                when "0110" =>
                  \$18454\ := "01000001";
                when "0111" =>
                  \$18454\ := "00011111";
                when "1000" =>
                  \$18454\ := "00000001";
                when "1001" =>
                  \$18454\ := "00001001";
                when "1010" =>
                  \$18454\ := "00010001";
                when "1011" =>
                  \$18454\ := "11000001";
                when "1100" =>
                  \$18454\ := "01100011";
                when "1101" =>
                  \$18454\ := "10000101";
                when "1110" =>
                  \$18454\ := "01100001";
                when "1111" =>
                  \$18454\ := "01110001";
                when others =>
                  \$18454\ := "11100011";
                end case;
                \$v4564\ := eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"13") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"12") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"11") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"10");
                case \$v4564\ is
                when "0000" =>
                  \$18455\ := "00000011";
                when "0001" =>
                  \$18455\ := "10011111";
                when "0010" =>
                  \$18455\ := "00100101";
                when "0011" =>
                  \$18455\ := "00001101";
                when "0100" =>
                  \$18455\ := "10011001";
                when "0101" =>
                  \$18455\ := "01001001";
                when "0110" =>
                  \$18455\ := "01000001";
                when "0111" =>
                  \$18455\ := "00011111";
                when "1000" =>
                  \$18455\ := "00000001";
                when "1001" =>
                  \$18455\ := "00001001";
                when "1010" =>
                  \$18455\ := "00010001";
                when "1011" =>
                  \$18455\ := "11000001";
                when "1100" =>
                  \$18455\ := "01100011";
                when "1101" =>
                  \$18455\ := "10000101";
                when "1110" =>
                  \$18455\ := "01100001";
                when "1111" =>
                  \$18455\ := "01110001";
                when others =>
                  \$18455\ := "11100011";
                end case;
                \$v4563\ := eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"17") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"16") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"15") & eclat_getBit(eclat_resize(\$18446_dur\,25) & X"000000" & X"14");
                case \$v4563\ is
                when "0000" =>
                  \$18456\ := "00000011";
                when "0001" =>
                  \$18456\ := "10011111";
                when "0010" =>
                  \$18456\ := "00100101";
                when "0011" =>
                  \$18456\ := "00001101";
                when "0100" =>
                  \$18456\ := "10011001";
                when "0101" =>
                  \$18456\ := "01001001";
                when "0110" =>
                  \$18456\ := "01000001";
                when "0111" =>
                  \$18456\ := "00011111";
                when "1000" =>
                  \$18456\ := "00000001";
                when "1001" =>
                  \$18456\ := "00001001";
                when "1010" =>
                  \$18456\ := "00010001";
                when "1011" =>
                  \$18456\ := "11000001";
                when "1100" =>
                  \$18456\ := "01100011";
                when "1101" =>
                  \$18456\ := "10000101";
                when "1110" =>
                  \$18456\ := "01100001";
                when "1111" =>
                  \$18456\ := "01110001";
                when others =>
                  \$18456\ := "11100011";
                end case;
                \$18448_dis\ := \$18451\ & \$18452\ & \$18453\ & \$18454\ & \$18455\ & \$18456\;
              else
                \$18448_dis\ := "00000011" & "00000011" & "00000011" & "00000011" & "00000011" & "00000011";
              end if;
              if \$v4339\(0) = '1' then
                
              else
                \$v4339\ := eclat_true;
                \$18450\ := X"0000000" & X"0";
              end if;
              \$18450\ := eclat_if(work.Int.eq(\$18450\, work.Int.add(
                                                         X"00" & X"989680", X"00" & X"989680")) & X"0000000" & X"0" & 
                          work.Int.add(\$18450\, X"0000000" & X"1"));
              \$18449\ := \$18450\;
              result4399 := ""&\$18443\(0) & work.Bool.lnot(""&\$18443\(1)) & 
              work.Int.gt(\$18449\, X"00" & X"989680") & ""&\$18443\(3) & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & \$18448_dis\;
              rdy4400 := eclat_true;
              state := IDLE4401;
            end if;
          end if;
        end if;
      end case;
      \state%next\ <= state;
      \state_var5924%next\ <= state_var5924;
      \state_var5923%next\ <= state_var5923;
      \state_var5922%next\ <= state_var5922;
      \state_var5921%next\ <= state_var5921;
      \state_var5920%next\ <= state_var5920;
      \$18606%next\ <= \$18606\;
      \$19190_binop_compare6454380_arg%next\ <= \$19190_binop_compare6454380_arg\;
      \$v4743%next\ <= \$v4743\;
      \$19072_binop_int6434370_arg%next\ <= \$19072_binop_int6434370_arg\;
      \$18910_modulo6684349_id%next\ <= \$18910_modulo6684349_id\;
      \$19299%next\ <= \$19299\;
      \$19069_modulo6684349_id%next\ <= \$19069_modulo6684349_id\;
      \$v5526%next\ <= \$v5526\;
      \$v4663%next\ <= \$v4663\;
      \$v5913%next\ <= \$v5913\;
      \$18602%next\ <= \$18602\;
      \$v5541%next\ <= \$v5541\;
      \$18809%next\ <= \$18809\;
      \$18751%next\ <= \$18751\;
      \$19272%next\ <= \$19272\;
      \$v5486%next\ <= \$v5486\;
      \$v5513%next\ <= \$v5513\;
      \$18729%next\ <= \$18729\;
      \$v5507%next\ <= \$v5507\;
      \$18801%next\ <= \$18801\;
      \$19779_loop666_id%next\ <= \$19779_loop666_id\;
      \$18775%next\ <= \$18775\;
      \$19874%next\ <= \$19874\;
      \$v5715%next\ <= \$v5715\;
      \$18974_modulo6684349_id%next\ <= \$18974_modulo6684349_id\;
      \$19828%next\ <= \$19828\;
      \$v4961%next\ <= \$v4961\;
      \$v4499%next\ <= \$v4499\;
      \$19326_compbranch6504387_result%next\ <= \$19326_compbranch6504387_result\;
      \$v5326%next\ <= \$v5326\;
      \$v5484%next\ <= \$v5484\;
      \$18504%next\ <= \$18504\;
      \$v5643%next\ <= \$v5643\;
      \$18945_modulo6684356_result%next\ <= \$18945_modulo6684356_result\;
      \$18933_modulo6684357_id%next\ <= \$18933_modulo6684357_id\;
      \$19250%next\ <= \$19250\;
      \$18624%next\ <= \$18624\;
      \$v4650%next\ <= \$v4650\;
      \$19553%next\ <= \$19553\;
      \$18637_w%next\ <= \$18637_w\;
      \$19380_compbranch6504393_id%next\ <= \$19380_compbranch6504393_id\;
      \$v5619%next\ <= \$v5619\;
      \$18835%next\ <= \$18835\;
      \$19579%next\ <= \$19579\;
      \$19758%next\ <= \$19758\;
      \$19085_modulo6684357_result%next\ <= \$19085_modulo6684357_result\;
      \$18776%next\ <= \$18776\;
      \$18875_v%next\ <= \$18875_v\;
      \$19132_modulo6684349_id%next\ <= \$19132_modulo6684349_id\;
      \$18619%next\ <= \$18619\;
      \$19163_forever6704376_arg%next\ <= \$19163_forever6704376_arg\;
      \$v4604%next\ <= \$v4604\;
      \$v5699%next\ <= \$v5699\;
      \$19292%next\ <= \$19292\;
      \$v5634%next\ <= \$v5634\;
      \$19416_w36574398_result%next\ <= \$19416_w36574398_result\;
      \$18993_modulo6684349_result%next\ <= \$18993_modulo6684349_result\;
      \$18581%next\ <= \$18581\;
      \$19866_hd%next\ <= \$19866_hd\;
      \$v5287%next\ <= \$v5287\;
      \$v4467%next\ <= \$v4467\;
      \$18900%next\ <= \$18900\;
      \$v4470%next\ <= \$v4470\;
      \$v4325%next\ <= \$v4325\;
      \$18696%next\ <= \$18696\;
      \$19245%next\ <= \$19245\;
      \$19024_modulo6684349_result%next\ <= \$19024_modulo6684349_result\;
      \$18945_modulo6684356_arg%next\ <= \$18945_modulo6684356_arg\;
      \$19689%next\ <= \$19689\;
      \$v4577%next\ <= \$v4577\;
      \$19140_r%next\ <= \$19140_r\;
      \$18802%next\ <= \$18802\;
      \$v5076%next\ <= \$v5076\;
      \$19001_r%next\ <= \$19001_r\;
      \$v5532%next\ <= \$v5532\;
      \$19501%next\ <= \$19501\;
      \$18769_hd%next\ <= \$18769_hd\;
      \$v5152%next\ <= \$v5152\;
      \$v4703%next\ <= \$v4703\;
      \$19122_modulo6684356_result%next\ <= \$19122_modulo6684356_result\;
      \$19499_aux664_id%next\ <= \$19499_aux664_id\;
      \$18483%next\ <= \$18483\;
      \$19290%next\ <= \$19290\;
      \$19273%next\ <= \$19273\;
      \$19104_modulo6684357_id%next\ <= \$19104_modulo6684357_id\;
      \$v4710%next\ <= \$v4710\;
      \$v4814%next\ <= \$v4814\;
      \$19170_res%next\ <= \$19170_res\;
      \$18924_res%next\ <= \$18924_res\;
      \$19863%next\ <= \$19863\;
      \$18821_v%next\ <= \$18821_v\;
      \$19827%next\ <= \$19827\;
      \$19432%next\ <= \$19432\;
      \$19448_v%next\ <= \$19448_v\;
      \$18630%next\ <= \$18630\;
      \$19094_v%next\ <= \$19094_v\;
      \$v4535%next\ <= \$v4535\;
      \$v5551%next\ <= \$v5551\;
      \$19028_modulo6684357_result%next\ <= \$19028_modulo6684357_result\;
      \$18939_binop_int6434363_result%next\ <= \$18939_binop_int6434363_result\;
      \$v5824%next\ <= \$v5824\;
      \$18788%next\ <= \$18788\;
      \$v5226%next\ <= \$v5226\;
      \$18582%next\ <= \$18582\;
      \$19081_modulo6684349_arg%next\ <= \$19081_modulo6684349_arg\;
      \$v5013%next\ <= \$v5013\;
      \$18881_hd%next\ <= \$18881_hd\;
      \$19525%next\ <= \$19525\;
      \$18509%next\ <= \$18509\;
      \$18793_make_block579_result%next\ <= \$18793_make_block579_result\;
      \$18974_modulo6684349_arg%next\ <= \$18974_modulo6684349_arg\;
      \$19235_v%next\ <= \$19235_v\;
      \$v4515%next\ <= \$v4515\;
      \$v5323%next\ <= \$v5323\;
      \$18655%next\ <= \$18655\;
      \$19906%next\ <= \$19906\;
      \$v5592%next\ <= \$v5592\;
      \$19194_res%next\ <= \$19194_res\;
      \$18990_modulo6684357_result%next\ <= \$18990_modulo6684357_result\;
      \$19947%next\ <= \$19947\;
      \$19672%next\ <= \$19672\;
      \$v5692%next\ <= \$v5692\;
      \$18474%next\ <= \$18474\;
      \$19641%next\ <= \$19641\;
      \$18855_next_env%next\ <= \$18855_next_env\;
      \$v5158%next\ <= \$v5158\;
      \$19040_modulo6684356_id%next\ <= \$19040_modulo6684356_id\;
      \$v5369%next\ <= \$v5369\;
      \$v5733%next\ <= \$v5733\;
      \$19661%next\ <= \$19661\;
      \$v5414%next\ <= \$v5414\;
      \$v4443%next\ <= \$v4443\;
      \$18876%next\ <= \$18876\;
      \$19653%next\ <= \$19653\;
      \$19508%next\ <= \$19508\;
      \$19358%next\ <= \$19358\;
      \$v5151%next\ <= \$v5151\;
      \$v5594%next\ <= \$v5594\;
      \$19043_modulo6684349_result%next\ <= \$19043_modulo6684349_result\;
      \$18859%next\ <= \$18859\;
      \$v4830%next\ <= \$v4830\;
      \$v5117%next\ <= \$v5117\;
      \$19445%next\ <= \$19445\;
      \$18867%next\ <= \$18867\;
      \$v5752%next\ <= \$v5752\;
      \$18865%next\ <= \$18865\;
      \$19890%next\ <= \$19890\;
      \$v4511%next\ <= \$v4511\;
      \$18455%next\ <= \$18455\;
      \$18512%next\ <= \$18512\;
      \$v4590%next\ <= \$v4590\;
      \$19427%next\ <= \$19427\;
      \$19934_hd%next\ <= \$19934_hd\;
      \$18846%next\ <= \$18846\;
      \$18524_loop666_result%next\ <= \$18524_loop666_result\;
      \$v4472%next\ <= \$v4472\;
      \$19723%next\ <= \$19723\;
      \$18778%next\ <= \$18778\;
      \$18694%next\ <= \$18694\;
      \$v5759%next\ <= \$v5759\;
      \$19066_modulo6684357_result%next\ <= \$19066_modulo6684357_result\;
      \$19850_w%next\ <= \$19850_w\;
      \$19419%next\ <= \$19419\;
      \$18961_v%next\ <= \$18961_v\;
      \$19201_v%next\ <= \$19201_v\;
      \$v5703%next\ <= \$v5703\;
      \$19274_v%next\ <= \$19274_v\;
      \$19394_compbranch6504395_arg%next\ <= \$19394_compbranch6504395_arg\;
      \$v5320%next\ <= \$v5320\;
      \$19166_binop_compare6454377_arg%next\ <= \$19166_binop_compare6454377_arg\;
      \$v5212%next\ <= \$v5212\;
      \$19704%next\ <= \$19704\;
      \$19930%next\ <= \$19930\;
      \$v5721%next\ <= \$v5721\;
      \$19458%next\ <= \$19458\;
      \$19185_v%next\ <= \$19185_v\;
      \$v5586%next\ <= \$v5586\;
      \$18738_next%next\ <= \$18738_next\;
      \$19364_v%next\ <= \$19364_v\;
      \$v5234%next\ <= \$v5234\;
      \$v5760%next\ <= \$v5760\;
      \$18974_modulo6684349_result%next\ <= \$18974_modulo6684349_result\;
      \$19797_next%next\ <= \$19797_next\;
      \$18745_hd%next\ <= \$18745_hd\;
      \$18797_branch_if648_result%next\ <= \$18797_branch_if648_result\;
      \$19589_copy_root_in_ram6634353_id%next\ <= \$19589_copy_root_in_ram6634353_id\;
      \$v5766%next\ <= \$v5766\;
      \$19478_v%next\ <= \$19478_v\;
      \$19752%next\ <= \$19752\;
      \$v4616%next\ <= \$v4616\;
      \$19894%next\ <= \$19894\;
      \$19819%next\ <= \$19819\;
      \$19489%next\ <= \$19489\;
      \$v5776%next\ <= \$v5776\;
      \$v5019%next\ <= \$v5019\;
      \$18807%next\ <= \$18807\;
      \$19504%next\ <= \$19504\;
      \$18650%next\ <= \$18650\;
      \$18837%next\ <= \$18837\;
      \$18569%next\ <= \$18569\;
      \$19129_modulo6684357_id%next\ <= \$19129_modulo6684357_id\;
      \$18805%next\ <= \$18805\;
      \$v5869%next\ <= \$v5869\;
      \$19112%next\ <= \$19112\;
      \$19135_binop_int6434374_arg%next\ <= \$19135_binop_int6434374_arg\;
      \$19002_modulo6684356_arg%next\ <= \$19002_modulo6684356_arg\;
      \$v5515%next\ <= \$v5515\;
      \$19319%next\ <= \$19319\;
      \$v5646%next\ <= \$v5646\;
      \$v4952%next\ <= \$v4952\;
      \$v5610%next\ <= \$v5610\;
      \$v5683%next\ <= \$v5683\;
      \$18958_binop_int6434364_result%next\ <= \$18958_binop_int6434364_result\;
      \$19342%next\ <= \$19342\;
      \$19657%next\ <= \$19657\;
      \$19777%next\ <= \$19777\;
      \$19620%next\ <= \$19620\;
      \$18793_make_block579_id%next\ <= \$18793_make_block579_id\;
      \$18521_loop666_arg%next\ <= \$18521_loop666_arg\;
      \$19803%next\ <= \$19803\;
      \$19217%next\ <= \$19217\;
      \$v4949%next\ <= \$v4949\;
      \$19486%next\ <= \$19486\;
      \$v5857%next\ <= \$v5857\;
      \$18482%next\ <= \$18482\;
      \$v4692%next\ <= \$v4692\;
      \$19309_v%next\ <= \$19309_v\;
      \$18529%next\ <= \$18529\;
      \$19916%next\ <= \$19916\;
      \$v5686%next\ <= \$v5686\;
      \$v4854%next\ <= \$v4854\;
      \$v4628%next\ <= \$v4628\;
      \$18703%next\ <= \$18703\;
      \$v5506%next\ <= \$v5506\;
      \$v4926%next\ <= \$v4926\;
      \$19829%next\ <= \$19829\;
      \$v4523%next\ <= \$v4523\;
      \$v4569%next\ <= \$v4569\;
      \$v5749%next\ <= \$v5749\;
      \$19209_v%next\ <= \$19209_v\;
      \$19482%next\ <= \$19482\;
      \$19611%next\ <= \$19611\;
      \$19811_copy_root_in_ram6634341_id%next\ <= \$19811_copy_root_in_ram6634341_id\;
      \$19784%next\ <= \$19784\;
      \$18502%next\ <= \$18502\;
      \$v4770%next\ <= \$v4770\;
      \$18667_w%next\ <= \$18667_w\;
      \$19434%next\ <= \$19434\;
      \$19333_compbranch6504388_arg%next\ <= \$19333_compbranch6504388_arg\;
      \$19732%next\ <= \$19732\;
      \$19609%next\ <= \$19609\;
      \$19714_next%next\ <= \$19714_next\;
      \$18815%next\ <= \$18815\;
      \$v5210%next\ <= \$v5210\;
      \$18565%next\ <= \$18565\;
      \$v4491%next\ <= \$v4491\;
      \$19076_res%next\ <= \$19076_res\;
      \$v4727%next\ <= \$v4727\;
      \$19015_binop_int6434367_id%next\ <= \$19015_binop_int6434367_id\;
      \$18986_modulo6684349_arg%next\ <= \$18986_modulo6684349_arg\;
      \$v4734%next\ <= \$v4734\;
      \$19656%next\ <= \$19656\;
      \$19496_aux664_arg%next\ <= \$19496_aux664_arg\;
      \$18480%next\ <= \$18480\;
      \$v5537%next\ <= \$v5537\;
      \$18458%next\ <= \$18458\;
      \$18993_modulo6684349_arg%next\ <= \$18993_modulo6684349_arg\;
      \$v5655%next\ <= \$v5655\;
      \$19294%next\ <= \$19294\;
      \$v5828%next\ <= \$v5828\;
      \$19583%next\ <= \$19583\;
      \$v5838%next\ <= \$v5838\;
      \$19163_forever6704376_id%next\ <= \$19163_forever6704376_id\;
      \$18723%next\ <= \$18723\;
      \$v4481%next\ <= \$v4481\;
      \$v5640%next\ <= \$v5640\;
      \$19314%next\ <= \$19314\;
      \$18762%next\ <= \$18762\;
      \$19034_binop_int6434368_arg%next\ <= \$19034_binop_int6434368_arg\;
      \$v4728%next\ <= \$v4728\;
      \$v4596%next\ <= \$v4596\;
      \$19062_modulo6684349_result%next\ <= \$19062_modulo6684349_result\;
      \$18914_modulo6684357_arg%next\ <= \$18914_modulo6684357_arg\;
      \$18590%next\ <= \$18590\;
      \$19902%next\ <= \$19902\;
      \$18670%next\ <= \$18670\;
      \$v5604%next\ <= \$v5604\;
      \$19248%next\ <= \$19248\;
      \$19088_modulo6684349_result%next\ <= \$19088_modulo6684349_result\;
      \$19464%next\ <= \$19464\;
      \$19072_binop_int6434370_result%next\ <= \$19072_binop_int6434370_result\;
      \$v4761%next\ <= \$v4761\;
      \$19816%next\ <= \$19816\;
      \$19081_modulo6684349_result%next\ <= \$19081_modulo6684349_result\;
      \$v4845%next\ <= \$v4845\;
      \$v4631%next\ <= \$v4631\;
      \$19326_compbranch6504387_arg%next\ <= \$19326_compbranch6504387_arg\;
      \$v5035%next\ <= \$v5035\;
      \$18685%next\ <= \$18685\;
      \$v5603%next\ <= \$v5603\;
      \$19628_w%next\ <= \$19628_w\;
      \$v5582%next\ <= \$v5582\;
      \$18948_modulo6684349_arg%next\ <= \$18948_modulo6684349_arg\;
      \$v5060%next\ <= \$v5060\;
      \$18668_hd%next\ <= \$18668_hd\;
      \$v4552%next\ <= \$v4552\;
      \$19187_compare6444358_result%next\ <= \$19187_compare6444358_result\;
      \$v5378%next\ <= \$v5378\;
      \$19623%next\ <= \$19623\;
      \$v5052%next\ <= \$v5052\;
      \$v4946%next\ <= \$v4946\;
      \$18664%next\ <= \$18664\;
      \$18646%next\ <= \$18646\;
      \$18852%next\ <= \$18852\;
      \$18485%next\ <= \$18485\;
      \$19190_binop_compare6454380_result%next\ <= \$19190_binop_compare6454380_result\;
      \$19043_modulo6684349_arg%next\ <= \$19043_modulo6684349_arg\;
      \$v4936%next\ <= \$v4936\;
      \$v4417%next\ <= \$v4417\;
      \$18447%next\ <= \$18447\;
      \$v4992%next\ <= \$v4992\;
      \$v5702%next\ <= \$v5702\;
      \$18967_modulo6684349_arg%next\ <= \$18967_modulo6684349_arg\;
      \$v5481%next\ <= \$v5481\;
      \$18952_modulo6684357_result%next\ <= \$18952_modulo6684357_result\;
      \$18662%next\ <= \$18662\;
      \$18600%next\ <= \$18600\;
      \$v5244%next\ <= \$v5244\;
      \$19600%next\ <= \$19600\;
      \$19838_copy_root_in_ram6634340_result%next\ <= \$19838_copy_root_in_ram6634340_result\;
      \$19885%next\ <= \$19885\;
      \$19685%next\ <= \$19685\;
      \$19187_compare6444358_id%next\ <= \$19187_compare6444358_id\;
      \$18926_modulo6684356_id%next\ <= \$18926_modulo6684356_id\;
      \$19720_w%next\ <= \$19720_w\;
      \$v5530%next\ <= \$v5530\;
      \$18644%next\ <= \$18644\;
      \$18466_loop666_id%next\ <= \$18466_loop666_id\;
      \$18638_hd%next\ <= \$18638_hd\;
      \$v4674%next\ <= \$v4674\;
      \$v5250%next\ <= \$v5250\;
      \$18563%next\ <= \$18563\;
      \$19062_modulo6684349_id%next\ <= \$19062_modulo6684349_id\;
      \$18645%next\ <= \$18645\;
      \$19897%next\ <= \$19897\;
      \$19139_res%next\ <= \$19139_res\;
      \$19347_fill6534389_arg%next\ <= \$19347_fill6534389_arg\;
      \$19495_loop665_arg%next\ <= \$19495_loop665_arg\;
      \$v4695%next\ <= \$v4695\;
      \$18576%next\ <= \$18576\;
      \$18578%next\ <= \$18578\;
      \$18440_make_block579_arg%next\ <= \$18440_make_block579_arg\;
      \$19157_forever6704375_id%next\ <= \$19157_forever6704375_id\;
      \$19246_v%next\ <= \$19246_v\;
      \$19495_loop665_id%next\ <= \$19495_loop665_id\;
      \$19515_next%next\ <= \$19515_next\;
      \$v4563%next\ <= \$v4563\;
      \$v4908%next\ <= \$v4908\;
      \$18635%next\ <= \$18635\;
      \$19251%next\ <= \$19251\;
      \$19648%next\ <= \$19648\;
      \$18613_copy_root_in_ram6634346_id%next\ <= \$18613_copy_root_in_ram6634346_id\;
      \$19780_loop665_arg%next\ <= \$19780_loop665_arg\;
      \$18571_copy_root_in_ram6634345_arg%next\ <= \$18571_copy_root_in_ram6634345_arg\;
      \$v5120%next\ <= \$v5120\;
      \$19854%next\ <= \$19854\;
      \$v4988%next\ <= \$v4988\;
      \$v5607%next\ <= \$v5607\;
      \$19848%next\ <= \$19848\;
      \$19232%next\ <= \$19232\;
      \$19814%next\ <= \$19814\;
      \$v4680%next\ <= \$v4680\;
      \$18906_r%next\ <= \$18906_r\;
      \$v5127%next\ <= \$v5127\;
      \$18620%next\ <= \$18620\;
      \$19887%next\ <= \$19887\;
      \$19296_v%next\ <= \$19296_v\;
      \$18709%next\ <= \$18709\;
      \$v4805%next\ <= \$v4805\;
      \$v5514%next\ <= \$v5514\;
      \$18913_r%next\ <= \$18913_r\;
      \$18457%next\ <= \$18457\;
      \$19269%next\ <= \$19269\;
      \$19569%next\ <= \$19569\;
      \$v5823%next\ <= \$v5823\;
      \$v5164%next\ <= \$v5164\;
      \$19721_hd%next\ <= \$19721_hd\;
      \$v5831%next\ <= \$v5831\;
      \$v4740%next\ <= \$v4740\;
      \$v5308%next\ <= \$v5308\;
      \$v4995%next\ <= \$v4995\;
      \$v4601%next\ <= \$v4601\;
      \$18484%next\ <= \$18484\;
      \$18733%next\ <= \$18733\;
      \$v4660%next\ <= \$v4660\;
      \$19408_argument3%next\ <= \$19408_argument3\;
      \$18828_v%next\ <= \$18828_v\;
      \$19390_b%next\ <= \$19390_b\;
      \$19727%next\ <= \$19727\;
      \$18510%next\ <= \$18510\;
      \$19662%next\ <= \$19662\;
      \$v5577%next\ <= \$v5577\;
      \$19015_binop_int6434367_arg%next\ <= \$19015_binop_int6434367_arg\;
      \$19413%next\ <= \$19413\;
      \$v4584%next\ <= \$v4584\;
      \$19845%next\ <= \$19845\;
      \$19337_compare6444359_id%next\ <= \$19337_compare6444359_id\;
      \$19698%next\ <= \$19698\;
      \$18566%next\ <= \$18566\;
      \$18767%next\ <= \$18767\;
      \$19359%next\ <= \$19359\;
      \$18977_binop_int6434365_arg%next\ <= \$18977_binop_int6434365_arg\;
      \$v4878%next\ <= \$v4878\;
      \$19267_hd%next\ <= \$19267_hd\;
      \$19679%next\ <= \$19679\;
      \$v5195%next\ <= \$v5195\;
      \$v4433%next\ <= \$v4433\;
      \$18864%next\ <= \$18864\;
      \$18996_binop_int6434366_arg%next\ <= \$18996_binop_int6434366_arg\;
      \$19599%next\ <= \$19599\;
      \$19526_forever6704355_arg%next\ <= \$19526_forever6704355_arg\;
      \$19578%next\ <= \$19578\;
      \$18605%next\ <= \$18605\;
      \$19558%next\ <= \$19558\;
      \$19280%next\ <= \$19280\;
      \$v5278%next\ <= \$v5278\;
      \$v5557%next\ <= \$v5557\;
      \$19817%next\ <= \$19817\;
      \$19238_w6514383_arg%next\ <= \$19238_w6514383_arg\;
      \$v5284%next\ <= \$v5284\;
      \$v5905%next\ <= \$v5905\;
      \$19488%next\ <= \$19488\;
      \$19474%next\ <= \$19474\;
      \$v5564%next\ <= \$v5564\;
      \$18591%next\ <= \$18591\;
      \$v4568%next\ <= \$v4568\;
      \$v5883%next\ <= \$v5883\;
      \$v5555%next\ <= \$v5555\;
      \$19726%next\ <= \$19726\;
      \$v4842%next\ <= \$v4842\;
      \$18834_v%next\ <= \$18834_v\;
      \$19401_compbranch6504396_result%next\ <= \$19401_compbranch6504396_result\;
      \$18699%next\ <= \$18699\;
      \$18680%next\ <= \$18680\;
      \$19751%next\ <= \$19751\;
      \$19157_forever6704375_arg%next\ <= \$19157_forever6704375_arg\;
      \$18584_hd%next\ <= \$18584_hd\;
      \$19867%next\ <= \$19867\;
      \$v5465%next\ <= \$v5465\;
      \$18999_v%next\ <= \$18999_v\;
      \$18623%next\ <= \$18623\;
      \$19754%next\ <= \$19754\;
      \$19825%next\ <= \$19825\;
      \$19312_v%next\ <= \$19312_v\;
      \$18936_modulo6684349_arg%next\ <= \$18936_modulo6684349_arg\;
      \$18460%next\ <= \$18460\;
      \$19596%next\ <= \$19596\;
      \$18795_offsetclosure_n639_result%next\ <= \$18795_offsetclosure_n639_result\;
      \$19918%next\ <= \$19918\;
      \$v4328%next\ <= \$v4328\;
      \$19373_compbranch6504392_result%next\ <= \$19373_compbranch6504392_result\;
      \$v5247%next\ <= \$v5247\;
      \$v4543%next\ <= \$v4543\;
      \$v5420%next\ <= \$v5420\;
      \$19505%next\ <= \$19505\;
      \$18570%next\ <= \$18570\;
      \$v5263%next\ <= \$v5263\;
      \$19391_compare6444359_id%next\ <= \$19391_compare6444359_id\;
      \$v5835%next\ <= \$v5835\;
      \$18962_res%next\ <= \$18962_res\;
      \$18822_v%next\ <= \$18822_v\;
      \$v5614%next\ <= \$v5614\;
      \$v5027%next\ <= \$v5027\;
      \$18610%next\ <= \$18610\;
      \$v5069%next\ <= \$v5069\;
      \$18684%next\ <= \$18684\;
      \$19535_copy_root_in_ram6634354_id%next\ <= \$19535_copy_root_in_ram6634354_id\;
      \$v5860%next\ <= \$v5860\;
      \$v4414%next\ <= \$v4414\;
      \$v5237%next\ <= \$v5237\;
      \$19066_modulo6684357_arg%next\ <= \$19066_modulo6684357_arg\;
      \$19852%next\ <= \$19852\;
      \$18577%next\ <= \$18577\;
      \$v5533%next\ <= \$v5533\;
      \$18553_forever6704348_arg%next\ <= \$18553_forever6704348_arg\;
      \$19387_compbranch6504394_id%next\ <= \$19387_compbranch6504394_id\;
      \$18643%next\ <= \$18643\;
      \$18754%next\ <= \$18754\;
      \$18933_modulo6684357_arg%next\ <= \$18933_modulo6684357_arg\;
      \$19397_b%next\ <= \$19397_b\;
      \$19279_v%next\ <= \$19279_v\;
      \$18933_modulo6684357_result%next\ <= \$18933_modulo6684357_result\;
      \$v5485%next\ <= \$v5485\;
      \$19550%next\ <= \$19550\;
      \$18816%next\ <= \$18816\;
      \$19495_loop665_result%next\ <= \$19495_loop665_result\;
      \$v5516%next\ <= \$v5516\;
      \$v5180%next\ <= \$v5180\;
      \$18952_modulo6684357_arg%next\ <= \$18952_modulo6684357_arg\;
      \$19855%next\ <= \$19855\;
      \$v5426%next\ <= \$v5426\;
      \$19313%next\ <= \$19313\;
      \$v5542%next\ <= \$v5542\;
      \$19565%next\ <= \$19565\;
      \$v4863%next\ <= \$v4863\;
      \$18980_v%next\ <= \$18980_v\;
      \$18521_loop666_id%next\ <= \$18521_loop666_id\;
      \$v5870%next\ <= \$v5870\;
      \$19800_next%next\ <= \$19800_next\;
      \$19746%next\ <= \$19746\;
      \$19851_hd%next\ <= \$19851_hd\;
      \$18488%next\ <= \$18488\;
      \$18746%next\ <= \$18746\;
      \$v5203%next\ <= \$v5203\;
      \$19222%next\ <= \$19222\;
      \$v5290%next\ <= \$v5290\;
      \$18796_make_block_n646_id%next\ <= \$18796_make_block_n646_id\;
      \$19096_r%next\ <= \$19096_r\;
      \$19450_v%next\ <= \$19450_v\;
      \$19651%next\ <= \$19651\;
      \$v5130%next\ <= \$v5130\;
      \$v5595%next\ <= \$v5595\;
      \$v4699%next\ <= \$v4699\;
      \$18559_copy_root_in_ram6634347_result%next\ <= \$18559_copy_root_in_ram6634347_result\;
      \$18831%next\ <= \$18831\;
      \$v5123%next\ <= \$v5123\;
      \$18829%next\ <= \$18829\;
      \$19761%next\ <= \$19761\;
      \$19547_copy_root_in_ram6634352_result%next\ <= \$19547_copy_root_in_ram6634352_result\;
      \$v5737%next\ <= \$v5737\;
      \$19676%next\ <= \$19676\;
      \$18450%next\ <= \$18450\;
      \$18982_r%next\ <= \$18982_r\;
      \$19179_compare6444358_arg%next\ <= \$19179_compare6444358_arg\;
      \$v4462%next\ <= \$v4462\;
      \$18717%next\ <= \$18717\;
      \$v5148%next\ <= \$v5148\;
      \$18571_copy_root_in_ram6634345_id%next\ <= \$18571_copy_root_in_ram6634345_id\;
      \$v5170%next\ <= \$v5170\;
      \$19438%next\ <= \$19438\;
      \$19647%next\ <= \$19647\;
      \$19483%next\ <= \$19483\;
      \$19361_fill6544390_arg%next\ <= \$19361_fill6544390_arg\;
      \$19861%next\ <= \$19861\;
      \$19211_compare6444358_id%next\ <= \$19211_compare6444358_id\;
      \$19786%next\ <= \$19786\;
      \$18725%next\ <= \$18725\;
      \$18459%next\ <= \$18459\;
      \$19135_binop_int6434374_result%next\ <= \$19135_binop_int6434374_result\;
      \$v5546%next\ <= \$v5546\;
      \$19724%next\ <= \$19724\;
      \$18711_w%next\ <= \$18711_w\;
      \$18948_modulo6684349_result%next\ <= \$18948_modulo6684349_result\;
      \$v5144%next\ <= \$v5144\;
      \$19908%next\ <= \$19908\;
      \$19858%next\ <= \$19858\;
      \$18779%next\ <= \$18779\;
      \$v5272%next\ <= \$v5272\;
      \$18612%next\ <= \$18612\;
      \$19303%next\ <= \$19303\;
      \$19551%next\ <= \$19551\;
      \$v5269%next\ <= \$v5269\;
      \$19186_res%next\ <= \$19186_res\;
      \$18689%next\ <= \$18689\;
      \$19631%next\ <= \$19631\;
      \$18791_loop665_arg%next\ <= \$18791_loop665_arg\;
      \$18905_res%next\ <= \$18905_res\;
      \$19694%next\ <= \$19694\;
      \$18755%next\ <= \$18755\;
      \$v5795%next\ <= \$v5795\;
      \$v5202%next\ <= \$v5202\;
      \$v5565%next\ <= \$v5565\;
      \$v4923%next\ <= \$v4923\;
      \$19835%next\ <= \$19835\;
      \$19588%next\ <= \$19588\;
      \$v4943%next\ <= \$v4943\;
      \$19078_modulo6684356_id%next\ <= \$19078_modulo6684356_id\;
      \$v5317%next\ <= \$v5317\;
      \result4434%next\ <= result4434;
      \$v5512%next\ <= \$v5512\;
      \$18465%next\ <= \$18465\;
      \$v4484%next\ <= \$v4484\;
      \$18830_v%next\ <= \$18830_v\;
      \$19779_loop666_arg%next\ <= \$19779_loop666_arg\;
      \$19616%next\ <= \$19616\;
      \$v4792%next\ <= \$v4792\;
      \$19088_modulo6684349_arg%next\ <= \$19088_modulo6684349_arg\;
      \$19666%next\ <= \$19666\;
      \$19179_compare6444358_id%next\ <= \$19179_compare6444358_id\;
      \$19681_next%next\ <= \$19681_next\;
      \$18742%next\ <= \$18742\;
      \$18795_offsetclosure_n639_arg%next\ <= \$18795_offsetclosure_n639_arg\;
      \$19384_compare6444359_id%next\ <= \$19384_compare6444359_id\;
      \$18993_modulo6684349_id%next\ <= \$18993_modulo6684349_id\;
      \$19610%next\ <= \$19610\;
      \$18856_loop_push6494360_arg%next\ <= \$18856_loop_push6494360_arg\;
      \$19909_w%next\ <= \$19909_w\;
      \$19686%next\ <= \$19686\;
      \$v4975%next\ <= \$v4975\;
      \$19019_res%next\ <= \$19019_res\;
      \$v5534%next\ <= \$v5534\;
      \$18479%next\ <= \$18479\;
      \$18525_loop665_result%next\ <= \$18525_loop665_result\;
      \$v5893%next\ <= \$v5893\;
      \$19671%next\ <= \$19671\;
      \$v4475%next\ <= \$v4475\;
      \$18734%next\ <= \$18734\;
      \$19128_r%next\ <= \$19128_r\;
      \$19750%next\ <= \$19750\;
      \$19499_aux664_arg%next\ <= \$19499_aux664_arg\;
      \$19826%next\ <= \$19826\;
      \$18799_w1656_result%next\ <= \$18799_w1656_result\;
      \$18798_w652_result%next\ <= \$18798_w652_result\;
      \$18467_loop665_arg%next\ <= \$18467_loop665_arg\;
      \$19021_modulo6684356_id%next\ <= \$19021_modulo6684356_id\;
      \$19088_modulo6684349_id%next\ <= \$19088_modulo6684349_id\;
      \$19162%next\ <= \$19162\;
      \$v4851%next\ <= \$v4851\;
      \$19357_v%next\ <= \$19357_v\;
      \$19097_modulo6684356_result%next\ <= \$19097_modulo6684356_result\;
      \$v5580%next\ <= \$v5580\;
      \$19012_modulo6684349_id%next\ <= \$19012_modulo6684349_id\;
      \$18765%next\ <= \$18765\;
      \$v4893%next\ <= \$v4893\;
      \$v5329%next\ <= \$v5329\;
      \$19936%next\ <= \$19936\;
      \$19020_r%next\ <= \$19020_r\;
      \$19238_w6514383_result%next\ <= \$19238_w6514383_result\;
      \$v5601%next\ <= \$v5601\;
      \$18996_binop_int6434366_id%next\ <= \$18996_binop_int6434366_id\;
      \$v5511%next\ <= \$v5511\;
      \$v4570%next\ <= \$v4570\;
      \$19675%next\ <= \$19675\;
      \$18601%next\ <= \$18601\;
      \$v4565%next\ <= \$v4565\;
      \$18552%next\ <= \$18552\;
      \$19077_r%next\ <= \$19077_r\;
      \$v5545%next\ <= \$v5545\;
      \$v5031%next\ <= \$v5031\;
      \$v5456%next\ <= \$v5456\;
      \$v5161%next\ <= \$v5161\;
      \$19075_v%next\ <= \$19075_v\;
      \$18791_loop665_result%next\ <= \$18791_loop665_result\;
      \$18750%next\ <= \$18750\;
      \$18718%next\ <= \$18718\;
      \$19849%next\ <= \$19849\;
      \$19059_modulo6684356_arg%next\ <= \$19059_modulo6684356_arg\;
      \$v4724%next\ <= \$v4724\;
      \$19423_v%next\ <= \$19423_v\;
      \$19352%next\ <= \$19352\;
      \$19601_copy_root_in_ram6634352_result%next\ <= \$19601_copy_root_in_ram6634352_result\;
      \$18789%next\ <= \$18789\;
      \$18977_binop_int6434365_id%next\ <= \$18977_binop_int6434365_id\;
      \$v5789%next\ <= \$v5789\;
      \$v5450%next\ <= \$v5450\;
      \$18681%next\ <= \$18681\;
      \$19206_binop_compare6454382_arg%next\ <= \$19206_binop_compare6454382_arg\;
      \$v5010%next\ <= \$v5010\;
      \$19523%next\ <= \$19523\;
      \$18964_modulo6684356_id%next\ <= \$18964_modulo6684356_id\;
      \$19923%next\ <= \$19923\;
      \$19361_fill6544390_result%next\ <= \$19361_fill6544390_result\;
      \$19535_copy_root_in_ram6634354_arg%next\ <= \$19535_copy_root_in_ram6634354_arg\;
      \$19564%next\ <= \$19564\;
      \$18770%next\ <= \$18770\;
      \$19790%next\ <= \$19790\;
      \$19509%next\ <= \$19509\;
      \$18598_w%next\ <= \$18598_w\;
      \$18462%next\ <= \$18462\;
      \$19873%next\ <= \$19873\;
      \$v5496%next\ <= \$v5496\;
      \$v5573%next\ <= \$v5573\;
      \$19177_v%next\ <= \$19177_v\;
      \$19320_forever6704386_arg%next\ <= \$19320_forever6704386_arg\;
      \$19069_modulo6684349_arg%next\ <= \$19069_modulo6684349_arg\;
      \$v5225%next\ <= \$v5225\;
      \$v5611%next\ <= \$v5611\;
      \$v5063%next\ <= \$v5063\;
      \$v5393%next\ <= \$v5393\;
      \$19778%next\ <= \$19778\;
      \$19821%next\ <= \$19821\;
      \$v5174%next\ <= \$v5174\;
      \$18494%next\ <= \$18494\;
      \$19333_compbranch6504388_result%next\ <= \$19333_compbranch6504388_result\;
      \$19441_arg%next\ <= \$19441_arg\;
      \$18920_binop_int6434362_arg%next\ <= \$18920_binop_int6434362_arg\;
      \$v5080%next\ <= \$v5080\;
      \$18790_loop666_id%next\ <= \$18790_loop666_id\;
      \$v5763%next\ <= \$v5763\;
      \$v5618%next\ <= \$v5618\;
      \$18613_copy_root_in_ram6634346_result%next\ <= \$18613_copy_root_in_ram6634346_result\;
      \$19498_loop665_arg%next\ <= \$19498_loop665_arg\;
      \$19467_sp%next\ <= \$19467_sp\;
      \$v4799%next\ <= \$v4799\;
      \$19187_compare6444358_arg%next\ <= \$19187_compare6444358_arg\;
      \$v4860%next\ <= \$v4860\;
      \$18849%next\ <= \$18849\;
      \$18749%next\ <= \$18749\;
      \$18907_modulo6684356_id%next\ <= \$18907_modulo6684356_id\;
      \$19794%next\ <= \$19794\;
      \$18863%next\ <= \$18863\;
      \$19910_hd%next\ <= \$19910_hd\;
      \$18958_binop_int6434364_id%next\ <= \$18958_binop_int6434364_id\;
      \$v5135%next\ <= \$v5135\;
      \$v4495%next\ <= \$v4495\;
      \$19320_forever6704386_id%next\ <= \$19320_forever6704386_id\;
      \$19300%next\ <= \$19300\;
      \$19116_binop_int6434373_arg%next\ <= \$19116_binop_int6434373_arg\;
      \$v5147%next\ <= \$v5147\;
      \$v4899%next\ <= \$v4899\;
      \$19333_compbranch6504388_id%next\ <= \$19333_compbranch6504388_id\;
      \$19880_w%next\ <= \$19880_w\;
      \$v5730%next\ <= \$v5730\;
      \$19366_compbranch6504391_arg%next\ <= \$19366_compbranch6504391_arg\;
      \$v5007%next\ <= \$v5007\;
      \$19377_compare6444359_result%next\ <= \$19377_compare6444359_result\;
      \$19203_compare6444358_result%next\ <= \$19203_compare6444358_result\;
      \$v5570%next\ <= \$v5570\;
      \$19664%next\ <= \$19664\;
      \$19637%next\ <= \$19637\;
      \$18926_modulo6684356_result%next\ <= \$18926_modulo6684356_result\;
      \$v4431%next\ <= \$v4431\;
      \$18854_sp%next\ <= \$18854_sp\;
      \$19710%next\ <= \$19710\;
      \$19771%next\ <= \$19771\;
      \$19057_res%next\ <= \$19057_res\;
      \$18907_modulo6684356_arg%next\ <= \$18907_modulo6684356_arg\;
      \$18537%next\ <= \$18537\;
      \$19785%next\ <= \$19785\;
      \$18792_wait662_result%next\ <= \$18792_wait662_result\;
      \$18826%next\ <= \$18826\;
      \$19307_v%next\ <= \$19307_v\;
      \$19354_v%next\ <= \$19354_v\;
      \$19463%next\ <= \$19463\;
      \$19734%next\ <= \$19734\;
      \rdy4929%next\ <= rdy4929;
      \$18799_w1656_id%next\ <= \$18799_w1656_id\;
      \$19589_copy_root_in_ram6634353_result%next\ <= \$19589_copy_root_in_ram6634353_result\;
      \$18472%next\ <= \$18472\;
      \$v4666%next\ <= \$v4666\;
      \$19129_modulo6684357_arg%next\ <= \$19129_modulo6684357_arg\;
      \$v4458%next\ <= \$v4458\;
      \$18873_v%next\ <= \$18873_v\;
      \$19038_res%next\ <= \$19038_res\;
      \$19595%next\ <= \$19595\;
      \$19883%next\ <= \$19883\;
      \$18677%next\ <= \$18677\;
      \$19249%next\ <= \$19249\;
      \$v5266%next\ <= \$v5266\;
      \$19546%next\ <= \$19546\;
      \$v4767%next\ <= \$v4767\;
      \$v5189%next\ <= \$v5189\;
      \$v4442%next\ <= \$v4442\;
      \$19891%next\ <= \$19891\;
      \$v5649%next\ <= \$v5649\;
      \$v5199%next\ <= \$v5199\;
      \$19559_w%next\ <= \$19559_w\;
      \$19920%next\ <= \$19920\;
      \$v4549%next\ <= \$v4549\;
      \$18990_modulo6684357_id%next\ <= \$18990_modulo6684357_id\;
      \$19107_modulo6684349_arg%next\ <= \$19107_modulo6684349_arg\;
      \$18520%next\ <= \$18520\;
      \$19420_w06554397_result%next\ <= \$19420_w06554397_result\;
      \$18884_v%next\ <= \$18884_v\;
      \$18925_r%next\ <= \$18925_r\;
      \$19179_compare6444358_result%next\ <= \$19179_compare6444358_result\;
      \$19078_modulo6684356_arg%next\ <= \$19078_modulo6684356_arg\;
      \$v5103%next\ <= \$v5103\;
      \$19522%next\ <= \$19522\;
      \$19544%next\ <= \$19544\;
      \$19243%next\ <= \$19243\;
      \$19718%next\ <= \$19718\;
      \$19148_modulo6684357_arg%next\ <= \$19148_modulo6684357_arg\;
      \$19538%next\ <= \$19538\;
      \$19255%next\ <= \$19255\;
      \$v4571%next\ <= \$v4571\;
      \$19275%next\ <= \$19275\;
      \$19281%next\ <= \$19281\;
      \$18599_hd%next\ <= \$18599_hd\;
      \$19836%next\ <= \$19836\;
      \$v4872%next\ <= \$v4872\;
      \$19043_modulo6684349_id%next\ <= \$19043_modulo6684349_id\;
      \$19884%next\ <= \$19884\;
      \$19871%next\ <= \$19871\;
      \$18851%next\ <= \$18851\;
      \$19557%next\ <= \$19557\;
      \$19517%next\ <= \$19517\;
      \$19532_forever6704350_id%next\ <= \$19532_forever6704350_id\;
      \$18782%next\ <= \$18782\;
      \$18526_aux664_id%next\ <= \$18526_aux664_id\;
      \$v4696%next\ <= \$v4696\;
      \$19238_w6514383_id%next\ <= \$19238_w6514383_id\;
      \$19582%next\ <= \$19582\;
      \$v5344%next\ <= \$v5344\;
      \$19570%next\ <= \$19570\;
      \$v4619%next\ <= \$v4619\;
      \$19888%next\ <= \$19888\;
      \$18794_apply638_id%next\ <= \$18794_apply638_id\;
      \$19497_loop666_id%next\ <= \$19497_loop666_id\;
      \$v4651%next\ <= \$v4651\;
      \$18521_loop666_result%next\ <= \$18521_loop666_result\;
      \$19901%next\ <= \$19901\;
      \$18442_cy%next\ <= \$18442_cy\;
      \$19444%next\ <= \$19444\;
      \$18549%next\ <= \$18549\;
      \$v5468%next\ <= \$v5468\;
      \$18604%next\ <= \$18604\;
      \$18540%next\ <= \$18540\;
      \$18575%next\ <= \$18575\;
      \$19330_compare6444359_id%next\ <= \$19330_compare6444359_id\;
      \$19085_modulo6684357_arg%next\ <= \$19085_modulo6684357_arg\;
      \$19040_modulo6684356_result%next\ <= \$19040_modulo6684356_result\;
      \$19324_f0%next\ <= \$19324_f0\;
      \$v5083%next\ <= \$v5083\;
      \$19540%next\ <= \$19540\;
      \$v5817%next\ <= \$v5817\;
      \$19554%next\ <= \$19554\;
      \$19295%next\ <= \$19295\;
      \$19120_res%next\ <= \$19120_res\;
      \$18475%next\ <= \$18475\;
      \$18580%next\ <= \$18580\;
      \$v4612%next\ <= \$v4612\;
      \$19005_modulo6684349_arg%next\ <= \$19005_modulo6684349_arg\;
      \$v4518%next\ <= \$v4518\;
      \$v5637%next\ <= \$v5637\;
      \$18848%next\ <= \$18848\;
      \$19801%next\ <= \$19801\;
      \$18893_v%next\ <= \$18893_v\;
      \$19913%next\ <= \$19913\;
      \$19262_forever6704385_id%next\ <= \$19262_forever6704385_id\;
      \$19210_res%next\ <= \$19210_res\;
      \$v5169%next\ <= \$v5169\;
      \$18514%next\ <= \$18514\;
      \$18747%next\ <= \$18747\;
      \$v5402%next\ <= \$v5402\;
      \$v5090%next\ <= \$v5090\;
      \$v4408%next\ <= \$v4408\;
      \$19304%next\ <= \$19304\;
      \$v5523%next\ <= \$v5523\;
      \$18505%next\ <= \$18505\;
      \$18888_next_acc%next\ <= \$18888_next_acc\;
      \$19376_b%next\ <= \$19376_b\;
      \$18688%next\ <= \$18688\;
      \$19100_modulo6684349_arg%next\ <= \$19100_modulo6684349_arg\;
      \$19412_sp%next\ <= \$19412_sp\;
      \$v4407%next\ <= \$v4407\;
      \$v5447%next\ <= \$v5447\;
      \$19798%next\ <= \$19798\;
      \$v5003%next\ <= \$v5003\;
      \$v5873%next\ <= \$v5873\;
      \$19097_modulo6684356_arg%next\ <= \$19097_modulo6684356_arg\;
      \$v5550%next\ <= \$v5550\;
      \$19626%next\ <= \$19626\;
      \$19471%next\ <= \$19471\;
      \$18721%next\ <= \$18721\;
      \$18971_modulo6684357_id%next\ <= \$18971_modulo6684357_id\;
      \$18797_branch_if648_id%next\ <= \$18797_branch_if648_id\;
      \$v4704%next\ <= \$v4704\;
      \$19288_v%next\ <= \$19288_v\;
      \$v5390%next\ <= \$v5390\;
      \$19366_compbranch6504391_result%next\ <= \$19366_compbranch6504391_result\;
      \$v5462%next\ <= \$v5462\;
      \$19914%next\ <= \$19914\;
      \$v5311%next\ <= \$v5311\;
      \$18608%next\ <= \$18608\;
      \$19317%next\ <= \$19317\;
      \$19141_modulo6684356_result%next\ <= \$19141_modulo6684356_result\;
      \$18511%next\ <= \$18511\;
      \$v4671%next\ <= \$v4671\;
      \$19487%next\ <= \$19487\;
      \$18522_loop665_arg%next\ <= \$18522_loop665_arg\;
      \$v4420%next\ <= \$v4420\;
      \$19625%next\ <= \$19625\;
      \$v5576%next\ <= \$v5576\;
      \$19886%next\ <= \$19886\;
      \$v5482%next\ <= \$v5482\;
      \result4928%next\ <= result4928;
      \$19773%next\ <= \$19773\;
      \$v4424%next\ <= \$v4424\;
      \$19787%next\ <= \$19787\;
      \$19104_modulo6684357_result%next\ <= \$19104_modulo6684357_result\;
      \$v5769%next\ <= \$v5769\;
      \$19496_aux664_result%next\ <= \$19496_aux664_result\;
      \$19717%next\ <= \$19717\;
      \$18647%next\ <= \$18647\;
      \$19155%next\ <= \$19155\;
      \$18661%next\ <= \$18661\;
      \$v4587%next\ <= \$v4587\;
      \$19939%next\ <= \$19939\;
      \$18832_v%next\ <= \$18832_v\;
      \$19227%next\ <= \$19227\;
      \$19650%next\ <= \$19650\;
      \$18495%next\ <= \$18495\;
      \$18551%next\ <= \$18551\;
      \$v5658%next\ <= \$v5658\;
      \$19276%next\ <= \$19276\;
      \$19859%next\ <= \$19859\;
      \$19325%next\ <= \$19325\;
      \$18977_binop_int6434365_result%next\ <= \$18977_binop_int6434365_result\;
      \$18944_r%next\ <= \$18944_r\;
      \$18527%next\ <= \$18527\;
      \$19119_v%next\ <= \$19119_v\;
      \$18648%next\ <= \$18648\;
      \$19793%next\ <= \$19793\;
      \$18877_v%next\ <= \$18877_v\;
      \$18939_binop_int6434363_id%next\ <= \$18939_binop_int6434363_id\;
      \$v5673%next\ <= \$v5673\;
      \$19190_binop_compare6454380_id%next\ <= \$19190_binop_compare6454380_id\;
      \$19842%next\ <= \$19842\;
      \$19144_modulo6684349_id%next\ <= \$19144_modulo6684349_id\;
      \$v5536%next\ <= \$v5536\;
      \$v5299%next\ <= \$v5299\;
      \$19601_copy_root_in_ram6634352_arg%next\ <= \$19601_copy_root_in_ram6634352_arg\;
      \$18539%next\ <= \$18539\;
      \$18936_modulo6684349_id%next\ <= \$18936_modulo6684349_id\;
      \$19015_binop_int6434367_result%next\ <= \$19015_binop_int6434367_result\;
      \$19171_compare6444358_id%next\ <= \$19171_compare6444358_id\;
      \$19597%next\ <= \$19597\;
      \$19581%next\ <= \$19581\;
      \$v4338%next\ <= \$v4338\;
      \$19384_compare6444359_result%next\ <= \$19384_compare6444359_result\;
      \$19748%next\ <= \$19748\;
      \$18522_loop665_id%next\ <= \$18522_loop665_id\;
      \$18461%next\ <= \$18461\;
      \$19256_v%next\ <= \$19256_v\;
      \$v5206%next\ <= \$v5206\;
      \$18824_v%next\ <= \$18824_v\;
      \$v5059%next\ <= \$v5059\;
      \$18657%next\ <= \$18657\;
      \$v5026%next\ <= \$v5026\;
      \$v4996%next\ <= \$v4996\;
      \$v5036%next\ <= \$v5036\;
      \$18825%next\ <= \$18825\;
      \$18806%next\ <= \$18806\;
      \$v4866%next\ <= \$v4866\;
      \$v4647%next\ <= \$v4647\;
      \$18891%next\ <= \$18891\;
      \$18843%next\ <= \$18843\;
      \$v4330%next\ <= \$v4330\;
      \$19370_compare6444359_id%next\ <= \$19370_compare6444359_id\;
      \$19601_copy_root_in_ram6634352_id%next\ <= \$19601_copy_root_in_ram6634352_id\;
      \$v5281%next\ <= \$v5281\;
      \$v4546%next\ <= \$v4546\;
      \$v4779%next\ <= \$v4779\;
      \$v4636%next\ <= \$v4636\;
      \$v4812%next\ <= \$v4812\;
      \$v5574%next\ <= \$v5574\;
      \$18526_aux664_arg%next\ <= \$18526_aux664_arg\;
      \$19308_v%next\ <= \$19308_v\;
      \$18793_make_block579_arg%next\ <= \$18793_make_block579_arg\;
      \$18437_loop666_arg%next\ <= \$18437_loop666_arg\;
      \$19206_binop_compare6454382_result%next\ <= \$19206_binop_compare6454382_result\;
      \$18444%next\ <= \$18444\;
      \$19066_modulo6684357_id%next\ <= \$19066_modulo6684357_id\;
      \$19046_r%next\ <= \$19046_r\;
      \$19837%next\ <= \$19837\;
      \$v5429%next\ <= \$v5429\;
      \$19571%next\ <= \$19571\;
      \$v4978%next\ <= \$v4978\;
      \$v4920%next\ <= \$v4920\;
      \$v5799%next\ <= \$v5799\;
      \$18524_loop666_arg%next\ <= \$18524_loop666_arg\;
      \$18810%next\ <= \$18810\;
      \$19944%next\ <= \$19944\;
      \$18880%next\ <= \$18880\;
      \$18869%next\ <= \$18869\;
      \$v5490%next\ <= \$v5490\;
      \$18659%next\ <= \$18659\;
      \$v5257%next\ <= \$v5257\;
      \$18945_modulo6684356_id%next\ <= \$18945_modulo6684356_id\;
      \$18683_hd%next\ <= \$18683_hd\;
      \$v4428%next\ <= \$v4428\;
      \$v5055%next\ <= \$v5055\;
      \$19774%next\ <= \$19774\;
      \$v5522%next\ <= \$v5522\;
      \$19783%next\ <= \$19783\;
      \$19125_modulo6684349_result%next\ <= \$19125_modulo6684349_result\;
      \$19097_modulo6684356_id%next\ <= \$19097_modulo6684356_id\;
      \$19507_next%next\ <= \$19507_next\;
      \rdy4400%next\ <= rdy4400;
      \$19542%next\ <= \$19542\;
      \$v5042%next\ <= \$v5042\;
      \$18813%next\ <= \$18813\;
      \$19220%next\ <= \$19220\;
      \$v4667%next\ <= \$v4667\;
      \$v4678%next\ <= \$v4678\;
      \$19211_compare6444358_result%next\ <= \$19211_compare6444358_result\;
      \$18790_loop666_result%next\ <= \$18790_loop666_result\;
      \$19804%next\ <= \$19804\;
      \$18622%next\ <= \$18622\;
      \$v4519%next\ <= \$v4519\;
      \$19667%next\ <= \$19667\;
      \$v4593%next\ <= \$v4593\;
      \$19811_copy_root_in_ram6634341_arg%next\ <= \$19811_copy_root_in_ram6634341_arg\;
      \$18695%next\ <= \$18695\;
      \$19789_next%next\ <= \$19789_next\;
      \$19259%next\ <= \$19259\;
      \$18437_loop666_id%next\ <= \$18437_loop666_id\;
      \$19203_compare6444358_id%next\ <= \$19203_compare6444358_id\;
      \$19788%next\ <= \$19788\;
      \$19141_modulo6684356_arg%next\ <= \$19141_modulo6684356_arg\;
      \$18473%next\ <= \$18473\;
      \$v5134%next\ <= \$v5134\;
      \$19144_modulo6684349_result%next\ <= \$19144_modulo6684349_result\;
      \$19932%next\ <= \$19932\;
      \$18603%next\ <= \$18603\;
      \$v5365%next\ <= \$v5365\;
      \$19701%next\ <= \$19701\;
      \$19543%next\ <= \$19543\;
      \$v5168%next\ <= \$v5168\;
      \$v4529%next\ <= \$v4529\;
      \$v4839%next\ <= \$v4839\;
      \$v4679%next\ <= \$v4679\;
      \$19796%next\ <= \$19796\;
      \$18845%next\ <= \$18845\;
      \$v5233%next\ <= \$v5233\;
      \$18438_loop665_arg%next\ <= \$18438_loop665_arg\;
      \$19337_compare6444359_arg%next\ <= \$19337_compare6444359_arg\;
      \$v4632%next\ <= \$v4632\;
      \$v4957%next\ <= \$v4957\;
      \$19336_b%next\ <= \$19336_b\;
      \$19709%next\ <= \$19709\;
      \$19031_modulo6684349_result%next\ <= \$19031_modulo6684349_result\;
      \$19824_hd%next\ <= \$19824_hd\;
      \$19619%next\ <= \$19619\;
      \$18546%next\ <= \$18546\;
      \$v5872%next\ <= \$v5872\;
      \$19818%next\ <= \$19818\;
      \$18971_modulo6684357_arg%next\ <= \$18971_modulo6684357_arg\;
      \$v4502%next\ <= \$v4502\;
      \$19326_compbranch6504387_id%next\ <= \$19326_compbranch6504387_id\;
      \$18531%next\ <= \$18531\;
      \$v4802%next\ <= \$v4802\;
      \$18841%next\ <= \$18841\;
      \$v4639%next\ <= \$v4639\;
      \$19466_sp%next\ <= \$19466_sp\;
      \$18567%next\ <= \$18567\;
      \$v4683%next\ <= \$v4683\;
      \$19643_w%next\ <= \$19643_w\;
      \$18649%next\ <= \$18649\;
      \$18929_modulo6684349_arg%next\ <= \$18929_modulo6684349_arg\;
      \$v5184%next\ <= \$v5184\;
      \$v4335%next\ <= \$v4335\;
      \$v5915%next\ <= \$v5915\;
      \$19169_v%next\ <= \$19169_v\;
      \$v5487%next\ <= \$v5487\;
      \$v5552%next\ <= \$v5552\;
      \$19361_fill6544390_id%next\ <= \$19361_fill6544390_id\;
      \$v5811%next\ <= \$v5811\;
      \$19512%next\ <= \$19512\;
      \$v4471%next\ <= \$v4471\;
      \$19725%next\ <= \$19725\;
      \$19844%next\ <= \$19844\;
      \$18732%next\ <= \$18732\;
      \$18618%next\ <= \$18618\;
      \$19387_compbranch6504394_arg%next\ <= \$19387_compbranch6504394_arg\;
      \$19027_r%next\ <= \$19027_r\;
      \$v5471%next\ <= \$v5471\;
      \$19659_hd%next\ <= \$19659_hd\;
      \$19875%next\ <= \$19875\;
      \$19639%next\ <= \$19639\;
      \$18470%next\ <= \$18470\;
      \$19310%next\ <= \$19310\;
      \$19815%next\ <= \$19815\;
      \$v5696%next\ <= \$v5696\;
      \$19350_v%next\ <= \$19350_v\;
      \$19503%next\ <= \$19503\;
      \$19182_binop_compare6454379_result%next\ <= \$19182_binop_compare6454379_result\;
      \$18955_modulo6684349_result%next\ <= \$18955_modulo6684349_result\;
      \$18476%next\ <= \$18476\;
      \$18443%next\ <= \$18443\;
      \$19230_v%next\ <= \$19230_v\;
      \$19018_v%next\ <= \$19018_v\;
      \$19713%next\ <= \$19713\;
      \$19218_v%next\ <= \$19218_v\;
      \$19009_modulo6684357_arg%next\ <= \$19009_modulo6684357_arg\;
      \$19498_loop665_result%next\ <= \$19498_loop665_result\;
      \$v5198%next\ <= \$v5198\;
      \$19741%next\ <= \$19741\;
      \$v4581%next\ <= \$v4581\;
      \$19161%next\ <= \$19161\;
      \$19156%next\ <= \$19156\;
      \$19104_modulo6684357_arg%next\ <= \$19104_modulo6684357_arg\;
      \$18492%next\ <= \$18492\;
      \$v5571%next\ <= \$v5571\;
      \$v4615%next\ <= \$v4615\;
      \$19937%next\ <= \$19937\;
      \$18917_modulo6684349_arg%next\ <= \$18917_modulo6684349_arg\;
      \$v5384%next\ <= \$v5384\;
      \$18939_binop_int6434363_arg%next\ <= \$18939_binop_int6434363_arg\;
      \$19572%next\ <= \$19572\;
      \$18898%next\ <= \$18898\;
      \$19391_compare6444359_result%next\ <= \$19391_compare6444359_result\;
      \$v5563%next\ <= \$v5563\;
      \$18948_modulo6684349_id%next\ <= \$18948_modulo6684349_id\;
      \$v5897%next\ <= \$v5897\;
      \$19100_modulo6684349_id%next\ <= \$19100_modulo6684349_id\;
      \$19409_sp%next\ <= \$19409_sp\;
      \$18478%next\ <= \$18478\;
      \$19047_modulo6684357_result%next\ <= \$19047_modulo6684357_result\;
      \$19009_modulo6684357_result%next\ <= \$19009_modulo6684357_result\;
      \$v5072%next\ <= \$v5072\;
      \$18895_v%next\ <= \$18895_v\;
      \$18559_copy_root_in_ram6634347_id%next\ <= \$18559_copy_root_in_ram6634347_id\;
      \$18559_copy_root_in_ram6634347_arg%next\ <= \$18559_copy_root_in_ram6634347_arg\;
      \$19922%next\ <= \$19922\;
      \$19125_modulo6684349_id%next\ <= \$19125_modulo6684349_id\;
      \$18629%next\ <= \$18629\;
      \$v4887%next\ <= \$v4887\;
      \$v4556%next\ <= \$v4556\;
      \$v5453%next\ <= \$v5453\;
      \$19731%next\ <= \$19731\;
      \$19449%next\ <= \$19449\;
      \$18669%next\ <= \$18669\;
      \$18660%next\ <= \$18660\;
      \rdy4573%next\ <= rdy4573;
      \$18795_offsetclosure_n639_id%next\ <= \$18795_offsetclosure_n639_id\;
      \$19401_compbranch6504396_arg%next\ <= \$19401_compbranch6504396_arg\;
      \$19878%next\ <= \$19878\;
      \$v5066%next\ <= \$v5066\;
      \$18631%next\ <= \$18631\;
      \$v4327%next\ <= \$v4327\;
      \$19234_sp%next\ <= \$19234_sp\;
      \$18687%next\ <= \$18687\;
      \$19811_copy_root_in_ram6634341_result%next\ <= \$19811_copy_root_in_ram6634341_result\;
      \rdy4608%next\ <= rdy4608;
      \$19728%next\ <= \$19728\;
      \$v5492%next\ <= \$v5492\;
      \$19843%next\ <= \$19843\;
      \$19532_forever6704350_arg%next\ <= \$19532_forever6704350_arg\;
      \$19028_modulo6684357_id%next\ <= \$19028_modulo6684357_id\;
      \$18958_binop_int6434364_arg%next\ <= \$18958_binop_int6434364_arg\;
      \$v4700%next\ <= \$v4700\;
      \$19301_v%next\ <= \$19301_v\;
      \$v4940%next\ <= \$v4940\;
      \$19012_modulo6684349_result%next\ <= \$19012_modulo6684349_result\;
      \$19268%next\ <= \$19268\;
      \$19772%next\ <= \$19772\;
      \$19226%next\ <= \$19226\;
      \$v5727%next\ <= \$v5727\;
      \$18889_v%next\ <= \$18889_v\;
      \$19882%next\ <= \$19882\;
      \$19877%next\ <= \$19877\;
      \$19091_binop_int6434371_id%next\ <= \$19091_binop_int6434371_id\;
      \$v4796%next\ <= \$v4796\;
      \$18907_modulo6684356_result%next\ <= \$18907_modulo6684356_result\;
      \$19561%next\ <= \$19561\;
      \$19282_v%next\ <= \$19282_v\;
      \$19806%next\ <= \$19806\;
      \$19257_v%next\ <= \$19257_v\;
      \$19660%next\ <= \$19660\;
      \$18583_w%next\ <= \$18583_w\;
      \$v4818%next\ <= \$v4818\;
      \$v4750%next\ <= \$v4750\;
      \$19492%next\ <= \$19492\;
      \$18525_loop665_id%next\ <= \$18525_loop665_id\;
      \$19311%next\ <= \$19311\;
      \$19743%next\ <= \$19743\;
      \$v4775%next\ <= \$v4775\;
      \$v4713%next\ <= \$v4713\;
      \$19519%next\ <= \$19519\;
      \$19870%next\ <= \$19870\;
      \$v4540%next\ <= \$v4540\;
      \$19638%next\ <= \$19638\;
      \$v4821%next\ <= \$v4821\;
      \$v5664%next\ <= \$v5664\;
      \$19211_compare6444358_arg%next\ <= \$19211_compare6444358_arg\;
      \$18500%next\ <= \$18500\;
      \$18545_next%next\ <= \$18545_next\;
      \$19078_modulo6684356_result%next\ <= \$19078_modulo6684356_result\;
      \$19868%next\ <= \$19868\;
      \$19047_modulo6684357_id%next\ <= \$19047_modulo6684357_id\;
      \$18663%next\ <= \$18663\;
      \$18679%next\ <= \$18679\;
      \$19053_binop_int6434369_result%next\ <= \$19053_binop_int6434369_result\;
      \$v4937%next\ <= \$v4937\;
      \$v5305%next\ <= \$v5305\;
      \$18986_modulo6684349_result%next\ <= \$18986_modulo6684349_result\;
      \$19266%next\ <= \$19266\;
      \$19447_sp%next\ <= \$19447_sp\;
      \$19084_r%next\ <= \$19084_r\;
      \$19779_loop666_result%next\ <= \$19779_loop666_result\;
      \$v5825%next\ <= \$v5825\;
      \$18464_rdy%next\ <= \$18464_rdy\;
      \$19636%next\ <= \$19636\;
      \$19329_b%next\ <= \$19329_b\;
      \$v5596%next\ <= \$v5596\;
      \$19031_modulo6684349_id%next\ <= \$19031_modulo6684349_id\;
      \$19526_forever6704355_id%next\ <= \$19526_forever6704355_id\;
      \$19926%next\ <= \$19926\;
      \$19614_hd%next\ <= \$19614_hd\;
      \$19594%next\ <= \$19594\;
      \$18542_next%next\ <= \$18542_next\;
      \$18553_forever6704348_id%next\ <= \$18553_forever6704348_id\;
      \$19521%next\ <= \$19521\;
      \$19832%next\ <= \$19832\;
      \$v4455%next\ <= \$v4455\;
      \$v4640%next\ <= \$v4640\;
      \$19053_binop_int6434369_arg%next\ <= \$19053_binop_int6434369_arg\;
      \$18508%next\ <= \$18508\;
      \$19684%next\ <= \$19684\;
      \$19315%next\ <= \$19315\;
      \$19166_binop_compare6454377_id%next\ <= \$19166_binop_compare6454377_id\;
      \$19110%next\ <= \$19110\;
      \$19678%next\ <= \$19678\;
      \$v5405%next\ <= \$v5405\;
      \$v5622%next\ <= \$v5622\;
      \$v5188%next\ <= \$v5188\;
      \$v5138%next\ <= \$v5138\;
      \$19198_binop_compare6454381_result%next\ <= \$19198_binop_compare6454381_result\;
      \$v4972%next\ <= \$v4972\;
      \$19872%next\ <= \$19872\;
      \$19031_modulo6684349_arg%next\ <= \$19031_modulo6684349_arg\;
      \$19405_compare6444359_arg%next\ <= \$19405_compare6444359_arg\;
      \$v4754%next\ <= \$v4754\;
      \$v5254%next\ <= \$v5254\;
      \$v5275%next\ <= \$v5275\;
      \$18642%next\ <= \$18642\;
      \$19892%next\ <= \$19892\;
      \$v4339%next\ <= \$v4339\;
      \$v4532%next\ <= \$v4532\;
      \$v5260%next\ <= \$v5260\;
      \$19021_modulo6684356_arg%next\ <= \$19021_modulo6684356_arg\;
      \$18996_binop_int6434366_result%next\ <= \$18996_binop_int6434366_result\;
      \$19005_modulo6684349_id%next\ <= \$19005_modulo6684349_id\;
      \$18522_loop665_result%next\ <= \$18522_loop665_result\;
      \$18682_w%next\ <= \$18682_w\;
      \$18914_modulo6684357_id%next\ <= \$18914_modulo6684357_id\;
      \$18673%next\ <= \$18673\;
      \$19766%next\ <= \$19766\;
      \$v4558%next\ <= \$v4558\;
      \$19214%next\ <= \$19214\;
      \$19566%next\ <= \$19566\;
      \$v4337%next\ <= \$v4337\;
      \$v5096%next\ <= \$v5096\;
      \$v5359%next\ <= \$v5359\;
      \$19174_binop_compare6454378_result%next\ <= \$19174_binop_compare6454378_result\;
      \$19563%next\ <= \$19563\;
      \$v4606%next\ <= \$v4606\;
      \$v5141%next\ <= \$v5141\;
      \$18639%next\ <= \$18639\;
      \$19154%next\ <= \$19154\;
      \$18562%next\ <= \$18562\;
      \$v4449%next\ <= \$v4449\;
      \$v4605%next\ <= \$v4605\;
      \$v4539%next\ <= \$v4539\;
      \$18666%next\ <= \$18666\;
      \$19781_aux664_id%next\ <= \$19781_aux664_id\;
      \$18904_v%next\ <= \$18904_v\;
      \$18498%next\ <= \$18498\;
      \$v4562%next\ <= \$v4562\;
      \$19497_loop666_arg%next\ <= \$19497_loop666_arg\;
      \$18564%next\ <= \$18564\;
      \$v5335%next\ <= \$v5335\;
      \$19834%next\ <= \$19834\;
      \$19700%next\ <= \$19700\;
      \$19769%next\ <= \$19769\;
      \$19907%next\ <= \$19907\;
      \$18724%next\ <= \$18724\;
      \$19425%next\ <= \$19425\;
      \$19293%next\ <= \$19293\;
      \$19147_r%next\ <= \$19147_r\;
      \$19950%next\ <= \$19950\;
      \$19355%next\ <= \$19355\;
      \$19024_modulo6684349_id%next\ <= \$19024_modulo6684349_id\;
      \$19665%next\ <= \$19665\;
      \$19351%next\ <= \$19351\;
      \$19500%next\ <= \$19500\;
      \$v4833%next\ <= \$v4833\;
      \$v4791%next\ <= \$v4791\;
      \$v4746%next\ <= \$v4746\;
      \$v5524%next\ <= \$v5524\;
      \$19856%next\ <= \$19856\;
      \$18456%next\ <= \$18456\;
      \$19021_modulo6684356_result%next\ <= \$19021_modulo6684356_result\;
      \$v5560%next\ <= \$v5560\;
      \$v4751%next\ <= \$v4751\;
      \$18487%next\ <= \$18487\;
      \$19755%next\ <= \$19755\;
      \$19233%next\ <= \$19233\;
      \$18654%next\ <= \$18654\;
      \$v4911%next\ <= \$v4911\;
      \$v5743%next\ <= \$v5743\;
      \$19414%next\ <= \$19414\;
      \$19649%next\ <= \$19649\;
      \$18702%next\ <= \$18702\;
      \$18897%next\ <= \$18897\;
      \$v4496%next\ <= \$v4496\;
      \$18967_modulo6684349_result%next\ <= \$18967_modulo6684349_result\;
      \$v5477%next\ <= \$v5477\;
      \$v4675%next\ <= \$v4675\;
      \$v5107%next\ <= \$v5107\;
      \$19485%next\ <= \$19485\;
      \$v5597%next\ <= \$v5597\;
      \$19132_modulo6684349_arg%next\ <= \$19132_modulo6684349_arg\;
      \$18781%next\ <= \$18781\;
      \$19252_forever6704384_id%next\ <= \$19252_forever6704384_id\;
      \$v4984%next\ <= \$v4984\;
      \$v5753%next\ <= \$v5753\;
      \$18896_v%next\ <= \$18896_v\;
      \$18737%next\ <= \$18737\;
      \$18439_wait662_result%next\ <= \$18439_wait662_result\;
      \$v5102%next\ <= \$v5102\;
      \$v4813%next\ <= \$v4813\;
      \$v5432%next\ <= \$v5432\;
      \$19642%next\ <= \$19642\;
      \$18446_dur%next\ <= \$18446_dur\;
      \$18625_copy_root_in_ram6634345_id%next\ <= \$18625_copy_root_in_ram6634345_id\;
      \$v5314%next\ <= \$v5314\;
      \$v5540%next\ <= \$v5540\;
      \$19617%next\ <= \$19617\;
      \$19451%next\ <= \$19451\;
      \$18556_forever6704344_id%next\ <= \$18556_forever6704344_id\;
      \$19585%next\ <= \$19585\;
      \$18886%next\ <= \$18886\;
      \$18439_wait662_id%next\ <= \$18439_wait662_id\;
      \$v5441%next\ <= \$v5441\;
      \$19737%next\ <= \$19737\;
      \$19879%next\ <= \$19879\;
      \$19072_binop_int6434370_id%next\ <= \$19072_binop_int6434370_id\;
      \$19462%next\ <= \$19462\;
      \$18516%next\ <= \$18516\;
      \$18838_v%next\ <= \$18838_v\;
      \$v5502%next\ <= \$v5502\;
      \$v5814%next\ <= \$v5814\;
      \$v5845%next\ <= \$v5845\;
      \$18438_loop665_result%next\ <= \$18438_loop665_result\;
      \$19658_w%next\ <= \$19658_w\;
      \$19182_binop_compare6454379_arg%next\ <= \$19182_binop_compare6454379_arg\;
      \$18901_binop_int6434361_result%next\ <= \$18901_binop_int6434361_result\;
      \$18453%next\ <= \$18453\;
      \$19260%next\ <= \$19260\;
      \$v5605%next\ <= \$v5605\;
      \$18971_modulo6684357_result%next\ <= \$18971_modulo6684357_result\;
      \$19853%next\ <= \$19853\;
      \$v5131%next\ <= \$v5131\;
      \$18820_v%next\ <= \$18820_v\;
      \$18571_copy_root_in_ram6634345_result%next\ <= \$18571_copy_root_in_ram6634345_result\;
      \$18515%next\ <= \$18515\;
      \$v4689%next\ <= \$v4689\;
      \$18914_modulo6684357_result%next\ <= \$18914_modulo6684357_result\;
      \$v5497%next\ <= \$v5497\;
      \$19951%next\ <= \$19951\;
      \$19807%next\ <= \$19807\;
      \$19241_v%next\ <= \$19241_v\;
      \$19242%next\ <= \$19242\;
      \$19539%next\ <= \$19539\;
      \$18752%next\ <= \$18752\;
      \$v5544%next\ <= \$v5544\;
      \result4607%next\ <= result4607;
      \$19091_binop_int6434371_arg%next\ <= \$19091_binop_int6434371_arg\;
      \$19345%next\ <= \$19345\;
      \$v5491%next\ <= \$v5491\;
      \$18844%next\ <= \$18844\;
      \$18963_r%next\ <= \$18963_r\;
      \$v5652%next\ <= \$v5652\;
      \$v5876%next\ <= \$v5876\;
      \$19113_forever6704372_id%next\ <= \$19113_forever6704372_id\;
      \$19383_b%next\ <= \$19383_b\;
      \$19584%next\ <= \$19584\;
      \$19942%next\ <= \$19942\;
      \$19615%next\ <= \$19615\;
      \$18676%next\ <= \$18676\;
      \$v4514%next\ <= \$v4514\;
      \$19316%next\ <= \$19316\;
      \$19148_modulo6684357_id%next\ <= \$19148_modulo6684357_id\;
      \$v4492%next\ <= \$v4492\;
      \$v5347%next\ <= \$v5347\;
      \$v5411%next\ <= \$v5411\;
      \$18756%next\ <= \$18756\;
      \$19865_w%next\ <= \$19865_w\;
      \$18533%next\ <= \$18533\;
      \$19297_v%next\ <= \$19297_v\;
      \$18497%next\ <= \$18497\;
      \$19062_modulo6684349_arg%next\ <= \$19062_modulo6684349_arg\;
      \$19456%next\ <= \$19456\;
      \$v5909%next\ <= \$v5909\;
      \$v5356%next\ <= \$v5356\;
      \$v5584%next\ <= \$v5584\;
      \$v5023%next\ <= \$v5023\;
      \$18766%next\ <= \$18766\;
      \$19770%next\ <= \$19770\;
      \$v4960%next\ <= \$v4960\;
      \$18674%next\ <= \$18674\;
      \$18595%next\ <= \$18595\;
      \$19927%next\ <= \$19927\;
      \$v5293%next\ <= \$v5293\;
      \$v5525%next\ <= \$v5525\;
      \$18786%next\ <= \$18786\;
      \$19592%next\ <= \$19592\;
      \$18748%next\ <= \$18748\;
      \$18448_dis%next\ <= \$18448_dis\;
      \$19398_compare6444359_result%next\ <= \$19398_compare6444359_result\;
      \$19202_res%next\ <= \$19202_res\;
      \$18951_r%next\ <= \$18951_r\;
      \$19040_modulo6684356_arg%next\ <= \$19040_modulo6684356_arg\;
      \$v5724%next\ <= \$v5724\;
      \$18780%next\ <= \$18780\;
      \$18651%next\ <= \$18651\;
      \$19518_next%next\ <= \$19518_next\;
      \$19005_modulo6684349_result%next\ <= \$19005_modulo6684349_result\;
      \$18808%next\ <= \$18808\;
      \$18715%next\ <= \$18715\;
      \$19799%next\ <= \$19799\;
      \$v5505%next\ <= \$v5505\;
      \$v5867%next\ <= \$v5867\;
      \$19646%next\ <= \$19646\;
      \$19833%next\ <= \$19833\;
      \$19182_binop_compare6454379_id%next\ <= \$19182_binop_compare6454379_id\;
      \$v5000%next\ <= \$v5000\;
      \$v5185%next\ <= \$v5185\;
      \$v5034%next\ <= \$v5034\;
      \$18467_loop665_result%next\ <= \$18467_loop665_result\;
      \$v5222%next\ <= \$v5222\;
      \$v4782%next\ <= \$v4782\;
      \$19547_copy_root_in_ram6634352_id%next\ <= \$19547_copy_root_in_ram6634352_id\;
      \$19915%next\ <= \$19915\;
      \$19719%next\ <= \$19719\;
      \$18777%next\ <= \$18777\;
      \$18550%next\ <= \$18550\;
      \$18842%next\ <= \$18842\;
      \$18489%next\ <= \$18489\;
      \$18439_wait662_arg%next\ <= \$18439_wait662_arg\;
      \$19100_modulo6684349_result%next\ <= \$19100_modulo6684349_result\;
      \$19135_binop_int6434374_id%next\ <= \$19135_binop_int6434374_id\;
      \$18796_make_block_n646_arg%next\ <= \$18796_make_block_n646_arg\;
      \$v5084%next\ <= \$v5084\;
      \$v4654%next\ <= \$v4654\;
      \$19820%next\ <= \$19820\;
      \$18901_binop_int6434361_arg%next\ <= \$18901_binop_int6434361_arg\;
      \$18701%next\ <= \$18701\;
      \$18768_w%next\ <= \$18768_w\;
      \$19586%next\ <= \$19586\;
      \$v5709%next\ <= \$v5709\;
      \$18613_copy_root_in_ram6634346_arg%next\ <= \$18613_copy_root_in_ram6634346_arg\;
      \$19917%next\ <= \$19917\;
      \$19138_v%next\ <= \$19138_v\;
      \$19697%next\ <= \$19697\;
      \$v4423%next\ <= \$v4423\;
      \result4963%next\ <= result4963;
      \$18794_apply638_arg%next\ <= \$18794_apply638_arg\;
      \$18792_wait662_arg%next\ <= \$18792_wait662_arg\;
      \$18741%next\ <= \$18741\;
      \$18735%next\ <= \$18735\;
      \$v5039%next\ <= \$v5039\;
      \$19677%next\ <= \$19677\;
      \$v5296%next\ <= \$v5296\;
      \$18714%next\ <= \$18714\;
      \$19231%next\ <= \$19231\;
      \$v5689%next\ <= \$v5689\;
      \$v5251%next\ <= \$v5251\;
      \$19876%next\ <= \$19876\;
      \$v5606%next\ <= \$v5606\;
      \$v5670%next\ <= \$v5670\;
      \$18794_apply638_result%next\ <= \$18794_apply638_result\;
      \$19921%next\ <= \$19921\;
      \$19420_w06554397_id%next\ <= \$19420_w06554397_id\;
      \$v4719%next\ <= \$v4719\;
      \$19059_modulo6684356_id%next\ <= \$19059_modulo6684356_id\;
      \$19864%next\ <= \$19864\;
      \$19347_fill6534389_result%next\ <= \$19347_fill6534389_result\;
      \$v5099%next\ <= \$v5099\;
      \$19860%next\ <= \$19860\;
      \$19781_aux664_arg%next\ <= \$19781_aux664_arg\;
      \$v4827%next\ <= \$v4827\;
      \$18964_modulo6684356_arg%next\ <= \$18964_modulo6684356_arg\;
      \$v5802%next\ <= \$v5802\;
      \$v4917%next\ <= \$v4917\;
      \$19302%next\ <= \$19302\;
      \$v5368%next\ <= \$v5368\;
      \$19823_w%next\ <= \$19823_w\;
      \$v5494%next\ <= \$v5494\;
      \$19668%next\ <= \$19668\;
      \$19398_compare6444359_id%next\ <= \$19398_compare6444359_id\;
      \$18574%next\ <= \$18574\;
      \$19228_v%next\ <= \$19228_v\;
      \$v5079%next\ <= \$v5079\;
      \$19749%next\ <= \$19749\;
      \$19795%next\ <= \$19795\;
      \$19203_compare6444358_arg%next\ <= \$19203_compare6444358_arg\;
      \$19768%next\ <= \$19768\;
      \$v4809%next\ <= \$v4809\;
      \$19941%next\ <= \$19941\;
      \$v4902%next\ <= \$v4902\;
      \$18899%next\ <= \$18899\;
      \$19605%next\ <= \$19605\;
      \$19514%next\ <= \$19514\;
      \$v4836%next\ <= \$v4836\;
      \$18640%next\ <= \$18640\;
      \$v4716%next\ <= \$v4716\;
      \$v5396%next\ <= \$v5396\;
      \$19341%next\ <= \$19341\;
      \$18870_v%next\ <= \$18870_v\;
      \$19722%next\ <= \$19722\;
      \$19475%next\ <= \$19475\;
      \$v5353%next\ <= \$v5353\;
      \$v4953%next\ <= \$v4953\;
      \$19460%next\ <= \$19460\;
      \$19470%next\ <= \$19470\;
      \$19580%next\ <= \$19580\;
      \$19893%next\ <= \$19893\;
      \$v4597%next\ <= \$v4597\;
      \$v5051%next\ <= \$v5051\;
      \$v5679%next\ <= \$v5679\;
      \$v5630%next\ <= \$v5630\;
      \$19889%next\ <= \$19889\;
      \$18812%next\ <= \$18812\;
      \$v5543%next\ <= \$v5543\;
      \$18955_modulo6684349_id%next\ <= \$18955_modulo6684349_id\;
      \$19529_forever6704351_arg%next\ <= \$19529_forever6704351_arg\;
      \$v5556%next\ <= \$v5556\;
      \$19497_loop666_result%next\ <= \$19497_loop666_result\;
      \$18536%next\ <= \$18536\;
      \$19433%next\ <= \$19433\;
      \$v4857%next\ <= \$v4857\;
      \$19286%next\ <= \$19286\;
      \$19621%next\ <= \$19621\;
      \$18758%next\ <= \$18758\;
      \$19261%next\ <= \$19261\;
      \$v5566%next\ <= \$v5566\;
      \$v4881%next\ <= \$v4881\;
      \$19148_modulo6684357_result%next\ <= \$19148_modulo6684357_result\;
      \$v4795%next\ <= \$v4795\;
      \$19945%next\ <= \$19945\;
      \$v4466%next\ <= \$v4466\;
      \$v4824%next\ <= \$v4824\;
      \$19747%next\ <= \$19747\;
      \$19081_modulo6684349_id%next\ <= \$19081_modulo6684349_id\;
      \$19285%next\ <= \$19285\;
      \$v4884%next\ <= \$v4884\;
      \$v5863%next\ <= \$v5863\;
      \$19394_compbranch6504395_result%next\ <= \$19394_compbranch6504395_result\;
      \$19535_copy_root_in_ram6634354_result%next\ <= \$19535_copy_root_in_ram6634354_result\;
      \$v4758%next\ <= \$v4758\;
      \$v4488%next\ <= \$v4488\;
      \$19012_modulo6684349_arg%next\ <= \$19012_modulo6684349_arg\;
      \$18607%next\ <= \$18607\;
      \$19753%next\ <= \$19753\;
      \$18785%next\ <= \$18785\;
      \$19394_compbranch6504395_id%next\ <= \$19394_compbranch6504395_id\;
      \$v5894%next\ <= \$v5894\;
      \$18799_w1656_arg%next\ <= \$18799_w1656_arg\;
      \$18856_loop_push6494360_id%next\ <= \$18856_loop_push6494360_id\;
      \$v4981%next\ <= \$v4981\;
      \$19391_compare6444359_arg%next\ <= \$19391_compare6444359_arg\;
      \$19366_compbranch6504391_id%next\ <= \$19366_compbranch6504391_id\;
      \$v4771%next\ <= \$v4771\;
      \$19781_aux664_result%next\ <= \$19781_aux664_result\;
      \$19174_binop_compare6454378_id%next\ <= \$19174_binop_compare6454378_id\;
      \$19416_w36574398_arg%next\ <= \$19416_w36574398_arg\;
      \$v5627%next\ <= \$v5627\;
      \$19271%next\ <= \$19271\;
      \$v5126%next\ <= \$v5126\;
      \$18708%next\ <= \$18708\;
      \$19780_loop665_id%next\ <= \$19780_loop665_id\;
      \$18827%next\ <= \$18827\;
      \$v5890%next\ <= \$v5890\;
      \$18882_v%next\ <= \$18882_v\;
      \$18525_loop665_arg%next\ <= \$18525_loop665_arg\;
      \$v5623%next\ <= \$v5623\;
      \$19344%next\ <= \$19344\;
      \$19576%next\ <= \$19576\;
      \$19171_compare6444358_arg%next\ <= \$19171_compare6444358_arg\;
      \$19838_copy_root_in_ram6634340_id%next\ <= \$19838_copy_root_in_ram6634340_id\;
      \$v5387%next\ <= \$v5387\;
      \$19373_compbranch6504392_arg%next\ <= \$19373_compbranch6504392_arg\;
      \$v5602%next\ <= \$v5602\;
      \$18544%next\ <= \$18544\;
      \$v5773%next\ <= \$v5773\;
      \$18493%next\ <= \$18493\;
      \$18579%next\ <= \$18579\;
      \$v5444%next\ <= \$v5444\;
      \$19524%next\ <= \$19524\;
      \$19247%next\ <= \$19247\;
      \$19122_modulo6684356_id%next\ <= \$19122_modulo6684356_id\;
      \$v5585%next\ <= \$v5585\;
      \$19494_loop666_result%next\ <= \$19494_loop666_result\;
      \$19284%next\ <= \$19284\;
      \$19373_compbranch6504392_id%next\ <= \$19373_compbranch6504392_id\;
      \$19287_v%next\ <= \$19287_v\;
      \$19808_forever6704342_id%next\ <= \$19808_forever6704342_id\;
      \$v5459%next\ <= \$v5459\;
      \$19767%next\ <= \$19767\;
      \$v5181%next\ <= \$v5181\;
      \$19494_loop666_id%next\ <= \$19494_loop666_id\;
      \$19529_forever6704351_id%next\ <= \$19529_forever6704351_id\;
      \$v5782%next\ <= \$v5782\;
      \$19053_binop_int6434369_id%next\ <= \$19053_binop_int6434369_id\;
      \$v4478%next\ <= \$v4478\;
      \$v5495%next\ <= \$v5495\;
      \$v4505%next\ <= \$v4505\;
      \$18621%next\ <= \$18621\;
      \$19598%next\ <= \$19598\;
      \$v4774%next\ <= \$v4774\;
      \$18523_aux664_result%next\ <= \$18523_aux664_result\;
      \$v5919%next\ <= \$v5919\;
      \$19298_v%next\ <= \$19298_v\;
      \$18872_v%next\ <= \$18872_v\;
      \$18817_v%next\ <= \$18817_v\;
      \$19762%next\ <= \$19762\;
      \$19002_modulo6684356_id%next\ <= \$19002_modulo6684356_id\;
      \$v5695%next\ <= \$v5695\;
      \$v5770%next\ <= \$v5770\;
      \$19024_modulo6684349_arg%next\ <= \$19024_modulo6684349_arg\;
      \$18936_modulo6684349_result%next\ <= \$18936_modulo6684349_result\;
      \$19428%next\ <= \$19428\;
      \$18890_v%next\ <= \$18890_v\;
      \$v5561%next\ <= \$v5561\;
      \$18535%next\ <= \$18535\;
      \$19151_modulo6684349_arg%next\ <= \$19151_modulo6684349_arg\;
      \result4399%next\ <= result4399;
      \$19278%next\ <= \$19278\;
      \rdy4435%next\ <= rdy4435;
      \$19000_res%next\ <= \$19000_res\;
      \$18609%next\ <= \$18609\;
      \$18720%next\ <= \$18720\;
      \$19552%next\ <= \$19552\;
      \$18757%next\ <= \$18757\;
      \$v4459%next\ <= \$v4459\;
      \$19305%next\ <= \$19305\;
      \$18874%next\ <= \$18874\;
      \$18800%next\ <= \$18800\;
      \$19607%next\ <= \$19607\;
      \$v4557%next\ <= \$v4557\;
      \$19757%next\ <= \$19757\;
      \$v4536%next\ <= \$v4536\;
      \$19933_w%next\ <= \$19933_w\;
      \$v4487%next\ <= \$v4487\;
      \$19258%next\ <= \$19258\;
      \$v4720%next\ <= \$v4720\;
      \$19151_modulo6684349_id%next\ <= \$19151_modulo6684349_id\;
      \$19744_w%next\ <= \$19744_w\;
      \result4572%next\ <= result4572;
      \$19103_r%next\ <= \$19103_r\;
      \$v5562%next\ <= \$v5562\;
      \$19178_res%next\ <= \$19178_res\;
      \$19160%next\ <= \$19160\;
      \$19663%next\ <= \$19663\;
      \$18871%next\ <= \$18871\;
      \$v5332%next\ <= \$v5332\;
      \$v5045%next\ <= \$v5045\;
      \$19193_v%next\ <= \$19193_v\;
      \$v4670%next\ <= \$v4670\;
      \$v5880%next\ <= \$v5880\;
      \$v5030%next\ <= \$v5030\;
      \$18883_v%next\ <= \$18883_v\;
      \$v4333%next\ <= \$v4333\;
      \$v5572%next\ <= \$v5572\;
      \$18983_modulo6684356_result%next\ <= \$18983_modulo6684356_result\;
      \$19493%next\ <= \$19493\;
      \$19095_res%next\ <= \$19095_res\;
      \$v5756%next\ <= \$v5756\;
      \$18983_modulo6684356_arg%next\ <= \$18983_modulo6684356_arg\;
      \$v5114%next\ <= \$v5114\;
      \$v5192%next\ <= \$v5192\;
      \$19461%next\ <= \$19461\;
      \$19107_modulo6684349_result%next\ <= \$19107_modulo6684349_result\;
      \$18839%next\ <= \$18839\;
      \$v5341%next\ <= \$v5341\;
      \$v5626%next\ <= \$v5626\;
      \$19050_modulo6684349_id%next\ <= \$19050_modulo6684349_id\;
      \$18787%next\ <= \$18787\;
      \$18716%next\ <= \$18716\;
      \$19121_r%next\ <= \$19121_r\;
      \$19206_binop_compare6454382_id%next\ <= \$19206_binop_compare6454382_id\;
      \$18885_v%next\ <= \$18885_v\;
      \$18658%next\ <= \$18658\;
      \$v5851%next\ <= \$v5851\;
      \$19069_modulo6684349_result%next\ <= \$19069_modulo6684349_result\;
      \$v5111%next\ <= \$v5111\;
      \$18678%next\ <= \$18678\;
      \$19822%next\ <= \$19822\;
      \$v5510%next\ <= \$v5510\;
      \$18753%next\ <= \$18753\;
      \$v5848%next\ <= \$v5848\;
      \$19113_forever6704372_arg%next\ <= \$19113_forever6704372_arg\;
      \$18840_v%next\ <= \$18840_v\;
      \$v5362%next\ <= \$v5362\;
      \$v4905%next\ <= \$v4905\;
      \$18596%next\ <= \$18596\;
      \$v4553%next\ <= \$v4553\;
      \$v5218%next\ <= \$v5218\;
      \$18440_make_block579_result%next\ <= \$18440_make_block579_result\;
      \$19401_compbranch6504396_id%next\ <= \$19401_compbranch6504396_id\;
      \$19380_compbranch6504393_result%next\ <= \$19380_compbranch6504393_result\;
      \$19047_modulo6684357_arg%next\ <= \$19047_modulo6684357_arg\;
      \$18861%next\ <= \$18861\;
      \$19931%next\ <= \$19931\;
      \$19340_argument2%next\ <= \$19340_argument2\;
      \$v4991%next\ <= \$v4991\;
      \$18983_modulo6684356_id%next\ <= \$18983_modulo6684356_id\;
      \$v5591%next\ <= \$v5591\;
      \$v5211%next\ <= \$v5211\;
      \$18920_binop_int6434362_id%next\ <= \$18920_binop_int6434362_id\;
      \$v5531%next\ <= \$v5531\;
      \$19002_modulo6684356_result%next\ <= \$19002_modulo6684356_result\;
      \$v4890%next\ <= \$v4890\;
      \$18589%next\ <= \$18589\;
      \$19144_modulo6684349_arg%next\ <= \$19144_modulo6684349_arg\;
      \$v4600%next\ <= \$v4600\;
      \$19476_v%next\ <= \$19476_v\;
      \$19587%next\ <= \$19587\;
      \$19919%next\ <= \$19919\;
      \$19574_w%next\ <= \$19574_w\;
      \$19237_v%next\ <= \$19237_v\;
      \$19037_v%next\ <= \$19037_v\;
      \$v5483%next\ <= \$v5483\;
      \$19634%next\ <= \$19634\;
      \$18585%next\ <= \$18585\;
      \$v4432%next\ <= \$v4432\;
      \$19365%next\ <= \$19365\;
      \$v5736%next\ <= \$v5736\;
      \$v4332%next\ <= \$v4332\;
      \$19857%next\ <= \$19857\;
      \$v5868%next\ <= \$v5868\;
      \$18803%next\ <= \$18803\;
      \$19346_sp%next\ <= \$19346_sp\;
      \$18691%next\ <= \$18691\;
      \$19846%next\ <= \$19846\;
      \$v5841%next\ <= \$v5841\;
      \$19695%next\ <= \$19695\;
      \$19494_loop666_arg%next\ <= \$19494_loop666_arg\;
      \$v5177%next\ <= \$v5177\;
      \$v4707%next\ <= \$v4707\;
      \$19122_modulo6684356_arg%next\ <= \$19122_modulo6684356_arg\;
      \$v4737%next\ <= \$v4737\;
      \$v5712%next\ <= \$v5712\;
      \$19370_compare6444359_arg%next\ <= \$19370_compare6444359_arg\;
      \$19622%next\ <= \$19622\;
      \$v4567%next\ <= \$v4567\;
      \$v5500%next\ <= \$v5500\;
      \$19899%next\ <= \$19899\;
      \$v5918%next\ <= \$v5918\;
      \$v5408%next\ <= \$v5408\;
      \$19039_r%next\ <= \$19039_r\;
      \$18814%next\ <= \$18814\;
      \$19738%next\ <= \$19738\;
      \$19670%next\ <= \$19670\;
      \$19457%next\ <= \$19457\;
      \$19377_compare6444359_id%next\ <= \$19377_compare6444359_id\;
      \$19556%next\ <= \$19556\;
      \$19711%next\ <= \$19711\;
      \$v5808%next\ <= \$v5808\;
      \$19377_compare6444359_arg%next\ <= \$19377_compare6444359_arg\;
      \$19405_compare6444359_result%next\ <= \$19405_compare6444359_result\;
      \$v5593%next\ <= \$v5593\;
      \$19903_next%next\ <= \$19903_next\;
      \$18818_v%next\ <= \$18818_v\;
      \$18633%next\ <= \$18633\;
      \$18466_loop666_arg%next\ <= \$18466_loop666_arg\;
      \$19459%next\ <= \$19459\;
      \$19705%next\ <= \$19705\;
      \$19629_hd%next\ <= \$19629_hd\;
      \$18836_v%next\ <= \$18836_v\;
      \$19384_compare6444359_arg%next\ <= \$19384_compare6444359_arg\;
      \$18736%next\ <= \$18736\;
      \$v5110%next\ <= \$v5110\;
      \$18671%next\ <= \$18671\;
      \$18686%next\ <= \$18686\;
      \$v4526%next\ <= \$v4526\;
      \$18990_modulo6684357_arg%next\ <= \$18990_modulo6684357_arg\;
      \$v5493%next\ <= \$v5493\;
      \$19632%next\ <= \$19632\;
      \$v5871%next\ <= \$v5871\;
      \$18823_v%next\ <= \$18823_v\;
      \$18593%next\ <= \$18593\;
      \$v5229%next\ <= \$v5229\;
      \$v5302%next\ <= \$v5302\;
      \$18652_w%next\ <= \$18652_w\;
      \$19506%next\ <= \$19506\;
      \$19337_compare6444359_result%next\ <= \$19337_compare6444359_result\;
      \$v4411%next\ <= \$v4411\;
      \$19680%next\ <= \$19680\;
      \rdy4964%next\ <= rdy4964;
      \$18690%next\ <= \$18690\;
      \$v4755%next\ <= \$v4755\;
      \$v5615%next\ <= \$v5615\;
      \$19195_compare6444358_id%next\ <= \$19195_compare6444358_id\;
      \$19912%next\ <= \$19912\;
      \$18469_make_block579_arg%next\ <= \$18469_make_block579_arg\;
      \$18743%next\ <= \$18743\;
      \$19791%next\ <= \$19791\;
      \$19604%next\ <= \$19604\;
      \$v5805%next\ <= \$v5805\;
      \$19510%next\ <= \$19510\;
      \$18728%next\ <= \$18728\;
      \$19869%next\ <= \$19869\;
      \$19900%next\ <= \$19900\;
      \$19898%next\ <= \$19898\;
      \$19111%next\ <= \$19111\;
      \$18586%next\ <= \$18586\;
      \$18986_modulo6684349_id%next\ <= \$18986_modulo6684349_id\;
      \$18468_wait662_id%next\ <= \$18468_wait662_id\;
      \$19244_v%next\ <= \$19244_v\;
      \$19612%next\ <= \$19612\;
      \$v4785%next\ <= \$v4785\;
      \$19847%next\ <= \$19847\;
      \$19398_compare6444359_arg%next\ <= \$19398_compare6444359_arg\;
      \$v4987%next\ <= \$v4987\;
      \$19830%next\ <= \$19830\;
      \$19034_binop_int6434368_id%next\ <= \$19034_binop_int6434368_id\;
      \$18856_loop_push6494360_result%next\ <= \$18856_loop_push6494360_result\;
      \$19687_w%next\ <= \$19687_w\;
      \$19745_hd%next\ <= \$19745_hd\;
      \$18894_v%next\ <= \$18894_v\;
      \$v5887%next\ <= \$v5887\;
      \$18672%next\ <= \$18672\;
      \$18617%next\ <= \$18617\;
      \$19938%next\ <= \$19938\;
      \$18892_v%next\ <= \$18892_v\;
      \$19437%next\ <= \$19437\;
      \$18636%next\ <= \$18636\;
      \$18611%next\ <= \$18611\;
      \$19225%next\ <= \$19225\;
      \$19420_w06554397_arg%next\ <= \$19420_w06554397_arg\;
      \$18713%next\ <= \$18713\;
      \$18616%next\ <= \$18616\;
      \$18771%next\ <= \$18771\;
      \$v4635%next\ <= \$v4635\;
      \$v5792%next\ <= \$v5792\;
      \$18868_v%next\ <= \$18868_v\;
      \$v5106%next\ <= \$v5106\;
      \$18693%next\ <= \$18693\;
      \$18597%next\ <= \$18597\;
      \$18437_loop666_result%next\ <= \$18437_loop666_result\;
      \$19426%next\ <= \$19426\;
      \$19763%next\ <= \$19763\;
      \$v5575%next\ <= \$v5575\;
      \$v4747%next\ <= \$v4747\;
      \$v5381%next\ <= \$v5381\;
      \$19151_modulo6684349_result%next\ <= \$19151_modulo6684349_result\;
      \$v5474%next\ <= \$v5474\;
      \$18850%next\ <= \$18850\;
      \$18445_x%next\ <= \$18445_x\;
      \$18798_w652_arg%next\ <= \$18798_w652_arg\;
      \$18878%next\ <= \$18878\;
      \$v5820%next\ <= \$v5820\;
      \$v5022%next\ <= \$v5022\;
      \$v4968%next\ <= \$v4968\;
      \$v4686%next\ <= \$v4686\;
      \$19472%next\ <= \$19472\;
      \$v5718%next\ <= \$v5718\;
      \$19404_b%next\ <= \$19404_b\;
      \$v4446%next\ <= \$v4446\;
      \$19624%next\ <= \$19624\;
      \$18587%next\ <= \$18587\;
      \$v5906%next\ <= \$v5906\;
      \$18970_r%next\ <= \$18970_r\;
      \$19545%next\ <= \$19545\;
      \$18534_next%next\ <= \$18534_next\;
      \$19219%next\ <= \$19219\;
      \$18792_wait662_id%next\ <= \$18792_wait662_id\;
      \$19265_ofs%next\ <= \$19265_ofs\;
      \$19618%next\ <= \$19618\;
      \$19411%next\ <= \$19411\;
      \$19468_sp%next\ <= \$19468_sp\;
      \$18547%next\ <= \$18547\;
      \$19116_binop_int6434373_id%next\ <= \$19116_binop_int6434373_id\;
      \$19065_r%next\ <= \$19065_r\;
      \$19645%next\ <= \$19645\;
      \$19129_modulo6684357_result%next\ <= \$19129_modulo6684357_result\;
      \$v5155%next\ <= \$v5155\;
      \$v5219%next\ <= \$v5219\;
      \$19756%next\ <= \$19756\;
      \$18490%next\ <= \$18490\;
      \$18523_aux664_arg%next\ <= \$18523_aux664_arg\;
      \$v5375%next\ <= \$v5375\;
      \$19215_argument1%next\ <= \$19215_argument1\;
      \$18860%next\ <= \$18860\;
      \$v5898%next\ <= \$v5898\;
      \$v4643%next\ <= \$v4643\;
      \$19174_binop_compare6454378_arg%next\ <= \$19174_binop_compare6454378_arg\;
      \$v5581%next\ <= \$v5581\;
      \$v4999%next\ <= \$v4999\;
      \$18466_loop666_result%next\ <= \$18466_loop666_result\;
      \$18469_make_block579_result%next\ <= \$18469_make_block579_result\;
      \$18625_copy_root_in_ram6634345_result%next\ <= \$18625_copy_root_in_ram6634345_result\;
      \$19640%next\ <= \$19640\;
      \$v4657%next\ <= \$v4657\;
      \$v5501%next\ <= \$v5501\;
      \$19323%next\ <= \$19323\;
      \$v5631%next\ <= \$v5631\;
      \$19270%next\ <= \$19270\;
      \$19473%next\ <= \$19473\;
      \$19318%next\ <= \$19318\;
      \$19132_modulo6684349_result%next\ <= \$19132_modulo6684349_result\;
      \$18548%next\ <= \$18548\;
      \$18967_modulo6684349_id%next\ <= \$18967_modulo6684349_id\;
      \$18772%next\ <= \$18772\;
      \$18628%next\ <= \$18628\;
      \$19562%next\ <= \$19562\;
      \$18538%next\ <= \$18538\;
      \$18819_v%next\ <= \$18819_v\;
      \$19198_binop_compare6454381_arg%next\ <= \$19198_binop_compare6454381_arg\;
      \$19465_sp%next\ <= \$19465_sp\;
      \$18526_aux664_result%next\ <= \$18526_aux664_result\;
      \$19911%next\ <= \$19911\;
      \$v4914%next\ <= \$v4914\;
      \$19446_sp%next\ <= \$19446_sp\;
      \$18932_r%next\ <= \$18932_r\;
      \$v4463%next\ <= \$v4463\;
      \$19946%next\ <= \$19946\;
      \$19943%next\ <= \$19943\;
      \$v5372%next\ <= \$v5372\;
      \$19577%next\ <= \$19577\;
      \$18641%next\ <= \$18641\;
      \$18773%next\ <= \$18773\;
      \$v5740%next\ <= \$v5740\;
      \$18524_loop666_id%next\ <= \$18524_loop666_id\;
      \$18964_modulo6684356_result%next\ <= \$18964_modulo6684356_result\;
      \$v4427%next\ <= \$v4427\;
      \$19655%next\ <= \$19655\;
      \$19028_modulo6684357_arg%next\ <= \$19028_modulo6684357_arg\;
      \$v4788%next\ <= \$v4788\;
      \$19520%next\ <= \$19520\;
      \$v4875%next\ <= \$v4875\;
      \$19306_v%next\ <= \$19306_v\;
      \$v5567%next\ <= \$v5567\;
      \$v5521%next\ <= \$v5521\;
      \$v4644%next\ <= \$v4644\;
      \$19343_sp%next\ <= \$19343_sp\;
      \$18722%next\ <= \$18722\;
      \$19935%next\ <= \$19935\;
      \$19056_v%next\ <= \$19056_v\;
      \$18513%next\ <= \$18513\;
      \$18989_r%next\ <= \$18989_r\;
      \$18879_v%next\ <= \$18879_v\;
      \$v4956%next\ <= \$v4956\;
      \$19730%next\ <= \$19730\;
      \$18665%next\ <= \$18665\;
      \$v4452%next\ <= \$v4452\;
      \$v5783%next\ <= \$v5783\;
      \$18710%next\ <= \$18710\;
      \$v5676%next\ <= \$v5676\;
      \$19009_modulo6684357_id%next\ <= \$19009_modulo6684357_id\;
      \$19712%next\ <= \$19712\;
      \$19841%next\ <= \$19841\;
      \$18556_forever6704344_arg%next\ <= \$18556_forever6704344_arg\;
      \$19780_loop665_result%next\ <= \$19780_loop665_result\;
      \$19236_v%next\ <= \$19236_v\;
      \$19330_compare6444359_result%next\ <= \$19330_compare6444359_result\;
      \$v5600%next\ <= \$v5600\;
      \$19330_compare6444359_arg%next\ <= \$19330_compare6444359_arg\;
      \$18592%next\ <= \$18592\;
      \$19289%next\ <= \$19289\;
      \$19589_copy_root_in_ram6634353_arg%next\ <= \$19589_copy_root_in_ram6634353_arg\;
      \$v4778%next\ <= \$v4778\;
      \$19356%next\ <= \$19356\;
      \$19050_modulo6684349_arg%next\ <= \$19050_modulo6684349_arg\;
      \$v5241%next\ <= \$v5241\;
      \$18594%next\ <= \$18594\;
      \$v5680%next\ <= \$v5680\;
      \$18866_v%next\ <= \$18866_v\;
      \$v5877%next\ <= \$v5877\;
      \$19424%next\ <= \$19424\;
      \$v5587%next\ <= \$v5587\;
      \$19369_b%next\ <= \$19369_b\;
      \$18481%next\ <= \$18481\;
      \$19050_modulo6684349_result%next\ <= \$19050_modulo6684349_result\;
      \$19691%next\ <= \$19691\;
      \$18471%next\ <= \$18471\;
      \$19058_r%next\ <= \$19058_r\;
      \$19560_hd%next\ <= \$19560_hd\;
      \$19405_compare6444359_id%next\ <= \$19405_compare6444359_id\;
      \$v5901%next\ <= \$v5901\;
      \$v5435%next\ <= \$v5435\;
      \$19353%next\ <= \$19353\;
      \$19059_modulo6684356_result%next\ <= \$19059_modulo6684356_result\;
      \$18910_modulo6684349_arg%next\ <= \$18910_modulo6684349_arg\;
      \$v5706%next\ <= \$v5706\;
      \$18486%next\ <= \$18486\;
      \$18501%next\ <= \$18501\;
      \$18532%next\ <= \$18532\;
      \$v4764%next\ <= \$v4764\;
      \$19216_v%next\ <= \$19216_v\;
      \$19613_w%next\ <= \$19613_w\;
      \$18528%next\ <= \$18528\;
      \$19283%next\ <= \$19283\;
      \$v5338%next\ <= \$v5338\;
      \$19091_binop_int6434371_result%next\ <= \$19091_binop_int6434371_result\;
      \$v4962%next\ <= \$v4962\;
      \$19654%next\ <= \$19654\;
      \$v5842%next\ <= \$v5842\;
      \$v5527%next\ <= \$v5527\;
      \$18920_binop_int6434362_result%next\ <= \$18920_binop_int6434362_result\;
      \$19195_compare6444358_arg%next\ <= \$19195_compare6444358_arg\;
      \$v5910%next\ <= \$v5910\;
      \$18705_next%next\ <= \$18705_next\;
      \$19511%next\ <= \$19511\;
      \$v5902%next\ <= \$v5902\;
      \$19410%next\ <= \$19410\;
      \$18468_wait662_arg%next\ <= \$18468_wait662_arg\;
      \$v5504%next\ <= \$v5504\;
      \$v4522%next\ <= \$v4522\;
      \$18797_branch_if648_arg%next\ <= \$18797_branch_if648_arg\;
      \$19696%next\ <= \$19696\;
      \$18955_modulo6684349_arg%next\ <= \$18955_modulo6684349_arg\;
      \$19652%next\ <= \$19652\;
      \$19606%next\ <= \$19606\;
      \$19195_compare6444358_result%next\ <= \$19195_compare6444358_result\;
      \$v5006%next\ <= \$v5006\;
      \$18804%next\ <= \$18804\;
      \$18910_modulo6684349_result%next\ <= \$18910_modulo6684349_result\;
      \$19502%next\ <= \$19502\;
      \$v5583%next\ <= \$v5583\;
      \$18853_hd%next\ <= \$18853_hd\;
      \$v5746%next\ <= \$v5746\;
      \$v5048%next\ <= \$v5048\;
      \$19831%next\ <= \$19831\;
      \$19481%next\ <= \$19481\;
      \$18774%next\ <= \$18774\;
      \$19708%next\ <= \$19708\;
      \$18632%next\ <= \$18632\;
      \$18625_copy_root_in_ram6634345_arg%next\ <= \$18625_copy_root_in_ram6634345_arg\;
      \$v5834%next\ <= \$v5834\;
      \$19568%next\ <= \$19568\;
      \$v4723%next\ <= \$v4723\;
      \$18519%next\ <= \$18519\;
      \$v4580%next\ <= \$v4580\;
      \$19547_copy_root_in_ram6634352_arg%next\ <= \$19547_copy_root_in_ram6634352_arg\;
      \$19477_v%next\ <= \$19477_v\;
      \$18704%next\ <= \$18704\;
      \$18503%next\ <= \$18503\;
      \$18790_loop666_arg%next\ <= \$18790_loop666_arg\;
      \$v5854%next\ <= \$v5854\;
      \$19690%next\ <= \$19690\;
      \$v5786%next\ <= \$v5786\;
      \$19498_loop665_id%next\ <= \$19498_loop665_id\;
      \$v5864%next\ <= \$v5864\;
      \$v5886%next\ <= \$v5886\;
      \$18923_v%next\ <= \$18923_v\;
      \$v5914%next\ <= \$v5914\;
      \$v5798%next\ <= \$v5798\;
      \$v5016%next\ <= \$v5016\;
      \$19499_aux664_result%next\ <= \$19499_aux664_result\;
      \$v5554%next\ <= \$v5554\;
      \$18675%next\ <= \$18675\;
      \$18463%next\ <= \$18463\;
      \$19469%next\ <= \$19469\;
      \$18700%next\ <= \$18700\;
      \$18744_w%next\ <= \$18744_w\;
      \$v5087%next\ <= \$v5087\;
      \$18530%next\ <= \$18530\;
      \$v5423%next\ <= \$v5423\;
      \$v5215%next\ <= \$v5215\;
      \$18929_modulo6684349_result%next\ <= \$18929_modulo6684349_result\;
      \$19733%next\ <= \$19733\;
      \$18653_hd%next\ <= \$18653_hd\;
      \$19429%next\ <= \$19429\;
      \$18833%next\ <= \$18833\;
      \$v5165%next\ <= \$v5165\;
      \$18454%next\ <= \$18454\;
      \$18847%next\ <= \$18847\;
      \$v5553%next\ <= \$v5553\;
      \$v5075%next\ <= \$v5075\;
      \$18692%next\ <= \$18692\;
      \$18719%next\ <= \$18719\;
      \$19940%next\ <= \$19940\;
      \$18712_hd%next\ <= \$18712_hd\;
      \$v5417%next\ <= \$v5417\;
      \$19125_modulo6684349_arg%next\ <= \$19125_modulo6684349_arg\;
      \$18634%next\ <= \$18634\;
      \$19484%next\ <= \$19484\;
      \$18929_modulo6684349_id%next\ <= \$18929_modulo6684349_id\;
      \$19198_binop_compare6454381_id%next\ <= \$19198_binop_compare6454381_id\;
      \$19416_w36574398_id%next\ <= \$19416_w36574398_id\;
      \$18798_w652_id%next\ <= \$18798_w652_id\;
      \$v5056%next\ <= \$v5056\;
      \$v4439%next\ <= \$v4439\;
      \$v5503%next\ <= \$v5503\;
      \$19608%next\ <= \$19608\;
      \$v5779%next\ <= \$v5779\;
      \$19277%next\ <= \$19277\;
      \$19223%next\ <= \$19223\;
      \$18499%next\ <= \$18499\;
      \$18796_make_block_n646_result%next\ <= \$18796_make_block_n646_result\;
      \$19085_modulo6684357_id%next\ <= \$19085_modulo6684357_id\;
      \$v5399%next\ <= \$v5399\;
      \$v4808%next\ <= \$v4808\;
      \$18811%next\ <= \$18811\;
      \$19808_forever6704342_arg%next\ <= \$19808_forever6704342_arg\;
      \$v4508%next\ <= \$v4508\;
      \$v5207%next\ <= \$v5207\;
      \$v5093%next\ <= \$v5093\;
      \$19034_binop_int6434368_result%next\ <= \$19034_binop_int6434368_result\;
      \$19627%next\ <= \$19627\;
      \$19881_hd%next\ <= \$19881_hd\;
      \$19291_v%next\ <= \$19291_v\;
      \$18901_binop_int6434361_id%next\ <= \$18901_binop_int6434361_id\;
      \$19387_compbranch6504394_result%next\ <= \$19387_compbranch6504394_result\;
      \$19644_hd%next\ <= \$19644_hd\;
      \$19347_fill6534389_id%next\ <= \$19347_fill6534389_id\;
      \$v5917%next\ <= \$v5917\;
      \$19792%next\ <= \$19792\;
      \$19541%next\ <= \$19541\;
      \$v5480%next\ <= \$v5480\;
      \$19415_sp%next\ <= \$19415_sp\;
      \$19262_forever6704385_arg%next\ <= \$19262_forever6704385_arg\;
      \$18477%next\ <= \$18477\;
      \$19635%next\ <= \$19635\;
      \$v4933%next\ <= \$v4933\;
      \$19633%next\ <= \$19633\;
      \$v4566%next\ <= \$v4566\;
      \$18917_modulo6684349_id%next\ <= \$18917_modulo6684349_id\;
      \$18451%next\ <= \$18451\;
      \$19802%next\ <= \$19802\;
      \$19221%next\ <= \$19221\;
      \$19224%next\ <= \$19224\;
      \$v5240%next\ <= \$v5240\;
      \$19516%next\ <= \$19516\;
      \$18656%next\ <= \$18656\;
      \$19693%next\ <= \$19693\;
      \$18496%next\ <= \$18496\;
      \$18588%next\ <= \$18588\;
      \$18887_v%next\ <= \$18887_v\;
      \$19360_sp%next\ <= \$19360_sp\;
      \$19171_compare6444358_result%next\ <= \$19171_compare6444358_result\;
      \$19688_hd%next\ <= \$19688_hd\;
      \$18491%next\ <= \$18491\;
      \$18541%next\ <= \$18541\;
      \$19380_compbranch6504393_arg%next\ <= \$19380_compbranch6504393_arg\;
      \$19782%next\ <= \$19782\;
      \$v5517%next\ <= \$v5517\;
      \$19141_modulo6684356_id%next\ <= \$19141_modulo6684356_id\;
      \$19107_modulo6684349_id%next\ <= \$19107_modulo6684349_id\;
      \$v4971%next\ <= \$v4971\;
      \$v4848%next\ <= \$v4848\;
      \$19166_binop_compare6454377_result%next\ <= \$19166_binop_compare6454377_result\;
      \$19593%next\ <= \$19593\;
      \$18568%next\ <= \$18568\;
      \$v4625%next\ <= \$v4625\;
      \$18452%next\ <= \$18452\;
      \$19742%next\ <= \$19742\;
      \$v4869%next\ <= \$v4869\;
      \$v5590%next\ <= \$v5590\;
      \$18468_wait662_result%next\ <= \$18468_wait662_result\;
      \$19575_hd%next\ <= \$19575_hd\;
      \$19229_v%next\ <= \$19229_v\;
      \$18981_res%next\ <= \$18981_res\;
      \$v4622%next\ <= \$v4622\;
      \$18942_v%next\ <= \$18942_v\;
      \$18543%next\ <= \$18543\;
      \$19513%next\ <= \$19513\;
      \$19555%next\ <= \$19555\;
      \$19692%next\ <= \$19692\;
      \$19370_compare6444359_result%next\ <= \$19370_compare6444359_result\;
      \$v4896%next\ <= \$v4896\;
      \$v5661%next\ <= \$v5661\;
      \$v5520%next\ <= \$v5520\;
      \$18917_modulo6684349_result%next\ <= \$18917_modulo6684349_result\;
      \$19116_binop_int6434373_result%next\ <= \$19116_binop_int6434373_result\;
      \$v4404%next\ <= \$v4404\;
      \$19862%next\ <= \$19862\;
      \$18449%next\ <= \$18449\;
      \$19573%next\ <= \$19573\;
      \$19729%next\ <= \$19729\;
      \$18952_modulo6684357_id%next\ <= \$18952_modulo6684357_id\;
      \$19252_forever6704384_arg%next\ <= \$19252_forever6704384_arg\;
      \$19805%next\ <= \$19805\;
      \$18943_res%next\ <= \$18943_res\;
      \$v4564%next\ <= \$v4564\;
      \$18926_modulo6684356_arg%next\ <= \$18926_modulo6684356_arg\;
      \$v5438%next\ <= \$v5438\;
      \$19567%next\ <= \$19567\;
      \$18761%next\ <= \$18761\;
      \$v5350%next\ <= \$v5350\;
      \$v5230%next\ <= \$v5230\;
      \$v4731%next\ <= \$v4731\;
      \$19838_copy_root_in_ram6634340_arg%next\ <= \$19838_copy_root_in_ram6634340_arg\;
      \$v5667%next\ <= \$v5667\;
      \$v5535%next\ <= \$v5535\;
      \$19008_r%next\ <= \$19008_r\;
      \$v5547%next\ <= \$v5547\;
      \$19669%next\ <= \$19669\;
      \$18862%next\ <= \$18862\;
      \$19699%next\ <= \$19699\;
      \$19630%next\ <= \$19630\;
      \$ram_lock%next\ <= \$ram_lock\;
      \$global_end_lock%next\ <= \$global_end_lock\;
      \$code_lock%next\ <= \$code_lock\;
      
      
      result <= result4399;
      end process;
  end architecture;
