-- code generated from the following source code:
--   stdlib.ecl
--   ../ocaml-vm/vm/mlvalue.ecl
--   ../ocaml-vm/vm/fail.ecl
--   ../ocaml-vm/vm/ram.ecl
--   ../ocaml-vm/vm/runtime.ecl
--   ../ocaml-vm/vm/debug.ecl
--   ../ocaml-vm/vm/alloc.ecl
--   ../ocaml-vm/vm/prims.ecl
--   ../ocaml-vm/bytecode.ecl
--   ../ocaml-vm/vm/vm.ecl
--   ../ocaml-vm/vm/target-specific/intel-max10/IOs.ecl
--   ../ocaml-vm/vm/target-specific/intel-max10/main.ecl
--
-- with the following command:
--
--    ./eclat -arg ((true,true,true,true,true,true,true,true,true,true),(true,false)) ../ocaml-vm/vm/mlvalue.ecl ../ocaml-vm/vm/fail.ecl ../ocaml-vm/vm/ram.ecl ../ocaml-vm/vm/runtime.ecl ../ocaml-vm/vm/debug.ecl ../ocaml-vm/vm/alloc.ecl ../ocaml-vm/vm/prims.ecl ../ocaml-vm/bytecode.ecl ../ocaml-vm/vm/vm.ecl ../ocaml-vm/vm/target-specific/intel-max10/IOs.ecl ../ocaml-vm/vm/target-specific/intel-max10/main.ecl

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.runtime.all;


entity main is
  
  port(signal clk    : in std_logic;
       signal reset  : in std_logic;
       signal argument : in value(0 to 11);
       signal result : out value(0 to 57));
       
end entity;
architecture rtl of main is

  type t_state is (IDLE5941, \$12520_LOOP666\, \$12521_LOOP665\, \$12522_WAIT662\, \$12523_MAKE_BLOCK579\, PAUSE_GET5945, PAUSE_GET5961, PAUSE_GET5965, PAUSE_GET5969, PAUSE_SET5942, PAUSE_SET5949, PAUSE_SET5952, PAUSE_SET5955, PAUSE_SET5958, PAUSE_SET6100, Q_WAIT5943, Q_WAIT5946, Q_WAIT5950, Q_WAIT5953, Q_WAIT5956, Q_WAIT5959, Q_WAIT5962, Q_WAIT5966, Q_WAIT5970, Q_WAIT6101);
  signal \state%now\, \state%next\: t_state;
  type t_state_var7464 is (IDLE5976, \$18632_LOOP666\, \$18633_LOOP665\, \$18634_AUX664\, \$18679_FOREVER6705881\, \$18686_COPY_ROOT_IN_RAM6635880\, \$18793_COPY_ROOT_IN_RAM6635879\, PAUSE_GET5980, PAUSE_GET5996, PAUSE_GET6000, PAUSE_GET6004, PAUSE_GET6008, PAUSE_GET6025, PAUSE_GET6029, PAUSE_GET6033, PAUSE_GET6037, PAUSE_GET6052, PAUSE_GET6056, PAUSE_GET6060, PAUSE_GET6073, PAUSE_GET6077, PAUSE_GET6090, PAUSE_GET6094, PAUSE_SET5977, PAUSE_SET5984, PAUSE_SET5987, PAUSE_SET5990, PAUSE_SET5993, PAUSE_SET6013, PAUSE_SET6016, PAUSE_SET6019, PAUSE_SET6022, PAUSE_SET6040, PAUSE_SET6043, PAUSE_SET6046, PAUSE_SET6049, PAUSE_SET6064, PAUSE_SET6067, PAUSE_SET6070, PAUSE_SET6081, PAUSE_SET6084, PAUSE_SET6087, Q_WAIT5978, Q_WAIT5981, Q_WAIT5985, Q_WAIT5988, Q_WAIT5991, Q_WAIT5994, Q_WAIT5997, Q_WAIT6001, Q_WAIT6005, Q_WAIT6009, Q_WAIT6014, Q_WAIT6017, Q_WAIT6020, Q_WAIT6023, Q_WAIT6026, Q_WAIT6030, Q_WAIT6034, Q_WAIT6038, Q_WAIT6041, Q_WAIT6044, Q_WAIT6047, Q_WAIT6050, Q_WAIT6053, Q_WAIT6057, Q_WAIT6061, Q_WAIT6065, Q_WAIT6068, Q_WAIT6071, Q_WAIT6074, Q_WAIT6078, Q_WAIT6082, Q_WAIT6085, Q_WAIT6088, Q_WAIT6091, Q_WAIT6095);
  signal \state_var7464%now\, \state_var7464%next\: t_state_var7464;
  type t_state_var7463 is (IDLE6149, \$12803_LOOP666\, \$12804_LOOP665\, \$12805_AUX664\, \$12806_LOOP666\, \$12807_LOOP665\, \$12808_AUX664\, \$12853_FOREVER6705887\, \$12857_FOREVER6705883\, \$12864_COPY_ROOT_IN_RAM6635886\, \$12891_COPY_ROOT_IN_RAM6635884\, \$13078_COPY_ROOT_IN_RAM6635885\, \$13105_COPY_ROOT_IN_RAM6635884\, PAUSE_GET6153, PAUSE_GET6169, PAUSE_GET6173, PAUSE_GET6177, PAUSE_GET6181, PAUSE_GET6188, PAUSE_GET6204, PAUSE_GET6208, PAUSE_GET6212, PAUSE_GET6216, PAUSE_GET6233, PAUSE_GET6237, PAUSE_GET6241, PAUSE_GET6257, PAUSE_GET6261, PAUSE_GET6265, PAUSE_GET6269, PAUSE_GET6284, PAUSE_GET6288, PAUSE_GET6292, PAUSE_GET6308, PAUSE_GET6312, PAUSE_GET6316, PAUSE_GET6329, PAUSE_GET6333, PAUSE_GET6346, PAUSE_GET6350, PAUSE_SET6150, PAUSE_SET6157, PAUSE_SET6160, PAUSE_SET6163, PAUSE_SET6166, PAUSE_SET6185, PAUSE_SET6192, PAUSE_SET6195, PAUSE_SET6198, PAUSE_SET6201, PAUSE_SET6221, PAUSE_SET6224, PAUSE_SET6227, PAUSE_SET6230, PAUSE_SET6245, PAUSE_SET6248, PAUSE_SET6251, PAUSE_SET6254, PAUSE_SET6272, PAUSE_SET6275, PAUSE_SET6278, PAUSE_SET6281, PAUSE_SET6296, PAUSE_SET6299, PAUSE_SET6302, PAUSE_SET6305, PAUSE_SET6320, PAUSE_SET6323, PAUSE_SET6326, PAUSE_SET6337, PAUSE_SET6340, PAUSE_SET6343, Q_WAIT6151, Q_WAIT6154, Q_WAIT6158, Q_WAIT6161, Q_WAIT6164, Q_WAIT6167, Q_WAIT6170, Q_WAIT6174, Q_WAIT6178, Q_WAIT6182, Q_WAIT6186, Q_WAIT6189, Q_WAIT6193, Q_WAIT6196, Q_WAIT6199, Q_WAIT6202, Q_WAIT6205, Q_WAIT6209, Q_WAIT6213, Q_WAIT6217, Q_WAIT6222, Q_WAIT6225, Q_WAIT6228, Q_WAIT6231, Q_WAIT6234, Q_WAIT6238, Q_WAIT6242, Q_WAIT6246, Q_WAIT6249, Q_WAIT6252, Q_WAIT6255, Q_WAIT6258, Q_WAIT6262, Q_WAIT6266, Q_WAIT6270, Q_WAIT6273, Q_WAIT6276, Q_WAIT6279, Q_WAIT6282, Q_WAIT6285, Q_WAIT6289, Q_WAIT6293, Q_WAIT6297, Q_WAIT6300, Q_WAIT6303, Q_WAIT6306, Q_WAIT6309, Q_WAIT6313, Q_WAIT6317, Q_WAIT6321, Q_WAIT6324, Q_WAIT6327, Q_WAIT6330, Q_WAIT6334, Q_WAIT6338, Q_WAIT6341, Q_WAIT6344, Q_WAIT6347, Q_WAIT6351);
  signal \state_var7463%now\, \state_var7463%next\: t_state_var7463;
  type t_state_var7462 is (IDLE6114, \$12679_LOOP666\, \$12680_LOOP665\, \$12681_WAIT662\, \$12682_MAKE_BLOCK579\, PAUSE_GET6118, PAUSE_GET6134, PAUSE_GET6138, PAUSE_GET6142, PAUSE_SET6115, PAUSE_SET6122, PAUSE_SET6125, PAUSE_SET6128, PAUSE_SET6131, PAUSE_SET6356, PAUSE_SET6359, PAUSE_SET6362, PAUSE_SET6365, PAUSE_SET6368, PAUSE_SET6371, PAUSE_SET6374, PAUSE_SET6377, PAUSE_SET6380, PAUSE_SET6383, PAUSE_SET6386, PAUSE_SET6389, PAUSE_SET6392, PAUSE_SET6395, PAUSE_SET6398, PAUSE_SET6401, PAUSE_SET6404, PAUSE_SET6407, PAUSE_SET6410, PAUSE_SET6413, PAUSE_SET6416, PAUSE_SET6419, PAUSE_SET6422, PAUSE_SET6425, PAUSE_SET6428, PAUSE_SET6431, PAUSE_SET6434, PAUSE_SET6437, PAUSE_SET6440, PAUSE_SET6443, PAUSE_SET6446, PAUSE_SET6449, PAUSE_SET6452, PAUSE_SET6455, PAUSE_SET6458, PAUSE_SET6461, PAUSE_SET6464, Q_WAIT6116, Q_WAIT6119, Q_WAIT6123, Q_WAIT6126, Q_WAIT6129, Q_WAIT6132, Q_WAIT6135, Q_WAIT6139, Q_WAIT6143, Q_WAIT6357, Q_WAIT6360, Q_WAIT6363, Q_WAIT6366, Q_WAIT6369, Q_WAIT6372, Q_WAIT6375, Q_WAIT6378, Q_WAIT6381, Q_WAIT6384, Q_WAIT6387, Q_WAIT6390, Q_WAIT6393, Q_WAIT6396, Q_WAIT6399, Q_WAIT6402, Q_WAIT6405, Q_WAIT6408, Q_WAIT6411, Q_WAIT6414, Q_WAIT6417, Q_WAIT6420, Q_WAIT6423, Q_WAIT6426, Q_WAIT6429, Q_WAIT6432, Q_WAIT6435, Q_WAIT6438, Q_WAIT6441, Q_WAIT6444, Q_WAIT6447, Q_WAIT6450, Q_WAIT6453, Q_WAIT6456, Q_WAIT6459, Q_WAIT6462, Q_WAIT6465);
  signal \state_var7462%now\, \state_var7462%next\: t_state_var7462;
  type t_state_var7461 is (IDLE6505, \$17455_LOOP666\, \$17456_LOOP665\, \$17457_AUX664\, \$17458_LOOP666\, \$17459_LOOP665\, \$17460_AUX664\, \$17505_FOREVER6705894\, \$17509_FOREVER6705890\, \$17513_FOREVER6705889\, \$17520_COPY_ROOT_IN_RAM6635893\, \$17547_COPY_ROOT_IN_RAM6635891\, \$17734_COPY_ROOT_IN_RAM6635892\, \$17761_COPY_ROOT_IN_RAM6635891\, PAUSE_GET6509, PAUSE_GET6525, PAUSE_GET6529, PAUSE_GET6533, PAUSE_GET6537, PAUSE_GET6544, PAUSE_GET6560, PAUSE_GET6564, PAUSE_GET6568, PAUSE_GET6572, PAUSE_GET6589, PAUSE_GET6593, PAUSE_GET6597, PAUSE_GET6613, PAUSE_GET6617, PAUSE_GET6621, PAUSE_GET6625, PAUSE_GET6640, PAUSE_GET6644, PAUSE_GET6648, PAUSE_GET6664, PAUSE_GET6668, PAUSE_GET6672, PAUSE_GET6685, PAUSE_GET6689, PAUSE_GET6702, PAUSE_GET6706, PAUSE_SET6506, PAUSE_SET6513, PAUSE_SET6516, PAUSE_SET6519, PAUSE_SET6522, PAUSE_SET6541, PAUSE_SET6548, PAUSE_SET6551, PAUSE_SET6554, PAUSE_SET6557, PAUSE_SET6577, PAUSE_SET6580, PAUSE_SET6583, PAUSE_SET6586, PAUSE_SET6601, PAUSE_SET6604, PAUSE_SET6607, PAUSE_SET6610, PAUSE_SET6628, PAUSE_SET6631, PAUSE_SET6634, PAUSE_SET6637, PAUSE_SET6652, PAUSE_SET6655, PAUSE_SET6658, PAUSE_SET6661, PAUSE_SET6676, PAUSE_SET6679, PAUSE_SET6682, PAUSE_SET6693, PAUSE_SET6696, PAUSE_SET6699, Q_WAIT6507, Q_WAIT6510, Q_WAIT6514, Q_WAIT6517, Q_WAIT6520, Q_WAIT6523, Q_WAIT6526, Q_WAIT6530, Q_WAIT6534, Q_WAIT6538, Q_WAIT6542, Q_WAIT6545, Q_WAIT6549, Q_WAIT6552, Q_WAIT6555, Q_WAIT6558, Q_WAIT6561, Q_WAIT6565, Q_WAIT6569, Q_WAIT6573, Q_WAIT6578, Q_WAIT6581, Q_WAIT6584, Q_WAIT6587, Q_WAIT6590, Q_WAIT6594, Q_WAIT6598, Q_WAIT6602, Q_WAIT6605, Q_WAIT6608, Q_WAIT6611, Q_WAIT6614, Q_WAIT6618, Q_WAIT6622, Q_WAIT6626, Q_WAIT6629, Q_WAIT6632, Q_WAIT6635, Q_WAIT6638, Q_WAIT6641, Q_WAIT6645, Q_WAIT6649, Q_WAIT6653, Q_WAIT6656, Q_WAIT6659, Q_WAIT6662, Q_WAIT6665, Q_WAIT6669, Q_WAIT6673, Q_WAIT6677, Q_WAIT6680, Q_WAIT6683, Q_WAIT6686, Q_WAIT6690, Q_WAIT6694, Q_WAIT6697, Q_WAIT6700, Q_WAIT6703, Q_WAIT6707);
  signal \state_var7461%now\, \state_var7461%next\: t_state_var7461;
  type t_state_var7460 is (IDLE6470, \$13920_LOOP666\, \$13921_LOOP665\, \$13922_WAIT662\, \$13923_MAKE_BLOCK579\, \$13924_APPLY638\, \$13925_OFFSETCLOSURE_N639\, \$13926_MAKE_BLOCK_N646\, \$13927_BRANCH_IF648\, \$13928_W652\, \$14207_LOOP_PUSH6495899\, \$14564_BINOP_INT6435900\, \$14589_MODULO6685895\, \$14597_MODULO6685888\, \$14613_MODULO6685896\, \$14621_MODULO6685888\, \$14644_BINOP_INT6435901\, \$14669_MODULO6685895\, \$14677_MODULO6685888\, \$14693_MODULO6685896\, \$14701_MODULO6685888\, \$14724_BINOP_INT6435902\, \$14749_MODULO6685895\, \$14757_MODULO6685888\, \$14773_MODULO6685896\, \$14781_MODULO6685888\, \$14804_BINOP_INT6435903\, \$14829_MODULO6685895\, \$14837_MODULO6685888\, \$14853_MODULO6685896\, \$14861_MODULO6685888\, \$14884_BINOP_INT6435904\, \$14909_MODULO6685895\, \$14917_MODULO6685888\, \$14933_MODULO6685896\, \$14941_MODULO6685888\, \$14964_BINOP_INT6435905\, \$14989_MODULO6685895\, \$14997_MODULO6685888\, \$15013_MODULO6685896\, \$15021_MODULO6685888\, \$15044_BINOP_INT6435906\, \$15069_MODULO6685895\, \$15077_MODULO6685888\, \$15093_MODULO6685896\, \$15101_MODULO6685888\, \$15124_BINOP_INT6435907\, \$15149_MODULO6685895\, \$15157_MODULO6685888\, \$15173_MODULO6685896\, \$15181_MODULO6685888\, \$15204_BINOP_INT6435908\, \$15229_MODULO6685895\, \$15237_MODULO6685888\, \$15253_MODULO6685896\, \$15261_MODULO6685888\, \$15284_BINOP_INT6435909\, \$15309_MODULO6685895\, \$15317_MODULO6685888\, \$15333_MODULO6685896\, \$15341_MODULO6685888\, \$15364_BINOP_INT6435910\, \$15389_MODULO6685895\, \$15397_MODULO6685888\, \$15413_MODULO6685896\, \$15421_MODULO6685888\, \$15447_FOREVER6705911\, \$15451_BINOP_INT6435912\, \$15476_MODULO6685895\, \$15484_MODULO6685888\, \$15500_MODULO6685896\, \$15508_MODULO6685888\, \$15531_BINOP_INT6435913\, \$15556_MODULO6685895\, \$15564_MODULO6685888\, \$15580_MODULO6685896\, \$15588_MODULO6685888\, \$15614_FOREVER6705914\, \$15621_FOREVER6705915\, \$15625_BINOP_COMPARE6455916\, \$15648_COMPARE6445897\, \$15661_BINOP_COMPARE6455917\, \$15684_COMPARE6445897\, \$15697_BINOP_COMPARE6455918\, \$15720_COMPARE6445897\, \$15733_BINOP_COMPARE6455919\, \$15756_COMPARE6445897\, \$15769_BINOP_COMPARE6455920\, \$15792_COMPARE6445897\, \$15805_BINOP_COMPARE6455921\, \$15828_COMPARE6445897\, \$16063_W6515922\, \$16158_FOREVER6705923\, \$16195_FOREVER6705924\, \$16510_FOREVER6705925\, \$16551_COMPBRANCH6505926\, \$16574_COMPARE6445898\, \$16589_COMPBRANCH6505927\, \$16612_COMPARE6445898\, \$16662_FILL6535928\, \$16752_FILL6545929\, \$16788_COMPBRANCH6505930\, \$16811_COMPARE6445898\, \$16823_COMPBRANCH6505931\, \$16846_COMPARE6445898\, \$16858_COMPBRANCH6505932\, \$16881_COMPARE6445898\, \$16893_COMPBRANCH6505933\, \$16916_COMPARE6445898\, \$16928_COMPBRANCH6505934\, \$16951_COMPARE6445898\, \$16963_COMPBRANCH6505935\, \$16986_COMPARE6445898\, \$17018_W36575938\, \$17048_W16565937\, \$17105_W06555936\, PAUSE_GET6474, PAUSE_GET6490, PAUSE_GET6494, PAUSE_GET6498, PAUSE_GET6715, PAUSE_GET6740, PAUSE_GET6744, PAUSE_GET6748, PAUSE_GET6756, PAUSE_GET6763, PAUSE_GET6771, PAUSE_GET6778, PAUSE_GET6782, PAUSE_GET6785, PAUSE_GET6788, PAUSE_GET6791, PAUSE_GET6794, PAUSE_GET6797, PAUSE_GET6800, PAUSE_GET6803, PAUSE_GET6812, PAUSE_GET6818, PAUSE_GET6824, PAUSE_GET6830, PAUSE_GET6836, PAUSE_GET6842, PAUSE_GET6848, PAUSE_GET6854, PAUSE_GET6857, PAUSE_GET6860, PAUSE_GET6863, PAUSE_GET6866, PAUSE_GET6872, PAUSE_GET6878, PAUSE_GET6884, PAUSE_GET6890, PAUSE_GET6896, PAUSE_GET6900, PAUSE_GET6915, PAUSE_GET6918, PAUSE_GET6921, PAUSE_GET6924, PAUSE_GET6930, PAUSE_GET6936, PAUSE_GET6942, PAUSE_GET6948, PAUSE_GET6951, PAUSE_GET6954, PAUSE_GET6957, PAUSE_GET6963, PAUSE_GET6966, PAUSE_GET6969, PAUSE_GET6972, PAUSE_GET6978, PAUSE_GET6981, PAUSE_GET6984, PAUSE_GET6987, PAUSE_GET6990, PAUSE_GET6993, PAUSE_GET6996, PAUSE_GET7018, PAUSE_GET7028, PAUSE_GET7038, PAUSE_GET7048, PAUSE_GET7058, PAUSE_GET7068, PAUSE_GET7078, PAUSE_GET7088, PAUSE_GET7098, PAUSE_GET7108, PAUSE_GET7118, PAUSE_GET7128, PAUSE_GET7138, PAUSE_GET7142, PAUSE_GET7146, PAUSE_GET7150, PAUSE_GET7154, PAUSE_GET7158, PAUSE_GET7162, PAUSE_GET7165, PAUSE_GET7168, PAUSE_GET7177, PAUSE_GET7180, PAUSE_GET7195, PAUSE_GET7198, PAUSE_GET7201, PAUSE_GET7204, PAUSE_GET7207, PAUSE_GET7211, PAUSE_GET7214, PAUSE_GET7217, PAUSE_GET7223, PAUSE_GET7237, PAUSE_GET7240, PAUSE_GET7252, PAUSE_GET7258, PAUSE_GET7261, PAUSE_GET7264, PAUSE_GET7280, PAUSE_GET7287, PAUSE_GET7294, PAUSE_GET7297, PAUSE_GET7304, PAUSE_GET7307, PAUSE_GET7310, PAUSE_GET7317, PAUSE_GET7320, PAUSE_GET7323, PAUSE_GET7326, PAUSE_GET7333, PAUSE_GET7336, PAUSE_GET7339, PAUSE_GET7342, PAUSE_GET7351, PAUSE_GET7356, PAUSE_GET7362, PAUSE_GET7373, PAUSE_GET7376, PAUSE_GET7379, PAUSE_GET7382, PAUSE_GET7391, PAUSE_GET7414, PAUSE_GET7424, PAUSE_GET7435, PAUSE_GET7439, PAUSE_GET7443, PAUSE_GET7447, PAUSE_GET7451, PAUSE_SET6471, PAUSE_SET6478, PAUSE_SET6481, PAUSE_SET6484, PAUSE_SET6487, PAUSE_SET6712, PAUSE_SET6718, PAUSE_SET6722, PAUSE_SET6726, PAUSE_SET6730, PAUSE_SET6733, PAUSE_SET6736, PAUSE_SET6753, PAUSE_SET6760, PAUSE_SET6767, PAUSE_SET6775, PAUSE_SET6806, PAUSE_SET6809, PAUSE_SET6815, PAUSE_SET6821, PAUSE_SET6827, PAUSE_SET6833, PAUSE_SET6839, PAUSE_SET6845, PAUSE_SET6851, PAUSE_SET6869, PAUSE_SET6875, PAUSE_SET6881, PAUSE_SET6887, PAUSE_SET6893, PAUSE_SET6903, PAUSE_SET6906, PAUSE_SET6909, PAUSE_SET6912, PAUSE_SET6927, PAUSE_SET6933, PAUSE_SET6939, PAUSE_SET6945, PAUSE_SET6960, PAUSE_SET6975, PAUSE_SET6999, PAUSE_SET7002, PAUSE_SET7005, PAUSE_SET7008, PAUSE_SET7171, PAUSE_SET7174, PAUSE_SET7183, PAUSE_SET7186, PAUSE_SET7189, PAUSE_SET7192, PAUSE_SET7220, PAUSE_SET7227, PAUSE_SET7230, PAUSE_SET7234, PAUSE_SET7243, PAUSE_SET7246, PAUSE_SET7249, PAUSE_SET7255, PAUSE_SET7268, PAUSE_SET7271, PAUSE_SET7274, PAUSE_SET7277, PAUSE_SET7284, PAUSE_SET7291, PAUSE_SET7301, PAUSE_SET7314, PAUSE_SET7330, PAUSE_SET7345, PAUSE_SET7348, PAUSE_SET7359, PAUSE_SET7366, PAUSE_SET7369, PAUSE_SET7385, PAUSE_SET7388, PAUSE_SET7395, PAUSE_SET7404, PAUSE_SET7408, PAUSE_SET7411, PAUSE_SET7417, PAUSE_SET7421, PAUSE_SET7428, PAUSE_SET7431, Q_WAIT6472, Q_WAIT6475, Q_WAIT6479, Q_WAIT6482, Q_WAIT6485, Q_WAIT6488, Q_WAIT6491, Q_WAIT6495, Q_WAIT6499, Q_WAIT6713, Q_WAIT6716, Q_WAIT6719, Q_WAIT6723, Q_WAIT6727, Q_WAIT6731, Q_WAIT6734, Q_WAIT6737, Q_WAIT6741, Q_WAIT6745, Q_WAIT6749, Q_WAIT6754, Q_WAIT6757, Q_WAIT6761, Q_WAIT6764, Q_WAIT6768, Q_WAIT6772, Q_WAIT6776, Q_WAIT6779, Q_WAIT6783, Q_WAIT6786, Q_WAIT6789, Q_WAIT6792, Q_WAIT6795, Q_WAIT6798, Q_WAIT6801, Q_WAIT6804, Q_WAIT6807, Q_WAIT6810, Q_WAIT6813, Q_WAIT6816, Q_WAIT6819, Q_WAIT6822, Q_WAIT6825, Q_WAIT6828, Q_WAIT6831, Q_WAIT6834, Q_WAIT6837, Q_WAIT6840, Q_WAIT6843, Q_WAIT6846, Q_WAIT6849, Q_WAIT6852, Q_WAIT6855, Q_WAIT6858, Q_WAIT6861, Q_WAIT6864, Q_WAIT6867, Q_WAIT6870, Q_WAIT6873, Q_WAIT6876, Q_WAIT6879, Q_WAIT6882, Q_WAIT6885, Q_WAIT6888, Q_WAIT6891, Q_WAIT6894, Q_WAIT6897, Q_WAIT6901, Q_WAIT6904, Q_WAIT6907, Q_WAIT6910, Q_WAIT6913, Q_WAIT6916, Q_WAIT6919, Q_WAIT6922, Q_WAIT6925, Q_WAIT6928, Q_WAIT6931, Q_WAIT6934, Q_WAIT6937, Q_WAIT6940, Q_WAIT6943, Q_WAIT6946, Q_WAIT6949, Q_WAIT6952, Q_WAIT6955, Q_WAIT6958, Q_WAIT6961, Q_WAIT6964, Q_WAIT6967, Q_WAIT6970, Q_WAIT6973, Q_WAIT6976, Q_WAIT6979, Q_WAIT6982, Q_WAIT6985, Q_WAIT6988, Q_WAIT6991, Q_WAIT6994, Q_WAIT6997, Q_WAIT7000, Q_WAIT7003, Q_WAIT7006, Q_WAIT7009, Q_WAIT7019, Q_WAIT7029, Q_WAIT7039, Q_WAIT7049, Q_WAIT7059, Q_WAIT7069, Q_WAIT7079, Q_WAIT7089, Q_WAIT7099, Q_WAIT7109, Q_WAIT7119, Q_WAIT7129, Q_WAIT7139, Q_WAIT7143, Q_WAIT7147, Q_WAIT7151, Q_WAIT7155, Q_WAIT7159, Q_WAIT7163, Q_WAIT7166, Q_WAIT7169, Q_WAIT7172, Q_WAIT7175, Q_WAIT7178, Q_WAIT7181, Q_WAIT7184, Q_WAIT7187, Q_WAIT7190, Q_WAIT7193, Q_WAIT7196, Q_WAIT7199, Q_WAIT7202, Q_WAIT7205, Q_WAIT7208, Q_WAIT7212, Q_WAIT7215, Q_WAIT7218, Q_WAIT7221, Q_WAIT7224, Q_WAIT7228, Q_WAIT7231, Q_WAIT7235, Q_WAIT7238, Q_WAIT7241, Q_WAIT7244, Q_WAIT7247, Q_WAIT7250, Q_WAIT7253, Q_WAIT7256, Q_WAIT7259, Q_WAIT7262, Q_WAIT7265, Q_WAIT7269, Q_WAIT7272, Q_WAIT7275, Q_WAIT7278, Q_WAIT7281, Q_WAIT7285, Q_WAIT7288, Q_WAIT7292, Q_WAIT7295, Q_WAIT7298, Q_WAIT7302, Q_WAIT7305, Q_WAIT7308, Q_WAIT7311, Q_WAIT7315, Q_WAIT7318, Q_WAIT7321, Q_WAIT7324, Q_WAIT7327, Q_WAIT7331, Q_WAIT7334, Q_WAIT7337, Q_WAIT7340, Q_WAIT7343, Q_WAIT7346, Q_WAIT7349, Q_WAIT7352, Q_WAIT7357, Q_WAIT7360, Q_WAIT7363, Q_WAIT7367, Q_WAIT7370, Q_WAIT7374, Q_WAIT7377, Q_WAIT7380, Q_WAIT7383, Q_WAIT7386, Q_WAIT7389, Q_WAIT7392, Q_WAIT7396, Q_WAIT7405, Q_WAIT7409, Q_WAIT7412, Q_WAIT7415, Q_WAIT7418, Q_WAIT7422, Q_WAIT7425, Q_WAIT7429, Q_WAIT7432, Q_WAIT7436, Q_WAIT7440, Q_WAIT7444, Q_WAIT7448, Q_WAIT7452);
  signal \state_var7460%now\, \state_var7460%next\: t_state_var7460;
  type array_value_16 is array (natural range <>) of value(0 to 15);
  type array_value_31 is array (natural range <>) of value(0 to 30);
  type array_value_32 is array (natural range <>) of value(0 to 31);
  signal ram : array_value_32(0 to 16383);
  signal \$ram_value\ : value(0 to 31) := (others => '0');
  signal \$ram_ptr\ : natural range 0 to 16383 := 0;
  signal \$ram_ptr_write\ : natural range 0 to 16383 := 0;
  signal \$ram_write\ : value(0 to 31) := (others => '0');
  signal \$ram_write_request\ : std_logic := '0';
  signal global_end : array_value_16(0 to 0);
  signal \$global_end_value\ : value(0 to 15) := (others => '0');
  signal \$global_end_ptr\ : natural range 0 to 0 := 0;
  signal \$global_end_ptr_write\ : natural range 0 to 0 := 0;
  signal \$global_end_write\ : value(0 to 15) := (others => '0');
  signal \$global_end_write_request\ : std_logic := '0';
  signal code : array_value_31(0 to 34);
  signal \$code_value\ : value(0 to 30) := (others => '0');
  signal \$code_ptr\ : natural range 0 to 34 := 0;
  signal \$code_ptr_write\ : natural range 0 to 34 := 0;
  signal \$code_write\ : value(0 to 30) := (others => '0');
  signal \$code_write_request\ : std_logic := '0';
  signal \$12670%next\, \$12670%now\ : value(0 to 1) := (others => '0');
  signal \$12807_loop665_arg%next\, \$12807_loop665_arg%now\, \$16651%next\, 
         \$16651%now\, \$17456_loop665_arg%next\, \$17456_loop665_arg%now\, 
         \$13921_loop665_arg%next\, \$13921_loop665_arg%now\, 
         \$12523_make_block579_result%next\, 
         \$12523_make_block579_result%now\, \$17105_w06555936_arg%next\, 
         \$17105_w06555936_arg%now\, \$16741%next\, \$16741%now\, 
         \$12680_loop665_arg%next\, \$12680_loop665_arg%now\, 
         \$12804_loop665_arg%next\, \$12804_loop665_arg%now\, \$17232%next\, 
         \$17232%now\, \$13923_make_block579_result%next\, 
         \$13923_make_block579_result%now\, 
         \$12682_make_block579_result%next\, 
         \$12682_make_block579_result%now\, \$18633_loop665_arg%next\, 
         \$18633_loop665_arg%now\, \$16024%next\, \$16024%now\, 
         \$12521_loop665_arg%next\, \$12521_loop665_arg%now\, \$17001%next\, 
         \$17001%now\, \$17459_loop665_arg%next\, \$17459_loop665_arg%now\ : value(0 to 95) := (others => '0');
  signal \$13928_w652_arg%next\, \$13928_w652_arg%now\, 
         \$16063_w6515922_arg%next\, \$16063_w6515922_arg%now\, 
         \$12805_aux664_arg%next\, \$12805_aux664_arg%now\, 
         \$12806_loop666_arg%next\, \$12806_loop666_arg%now\, 
         \$12808_aux664_arg%next\, \$12808_aux664_arg%now\, 
         \$14207_loop_push6495899_arg%next\, 
         \$14207_loop_push6495899_arg%now\, \$17460_aux664_arg%next\, 
         \$17460_aux664_arg%now\, \$18634_aux664_arg%next\, 
         \$18634_aux664_arg%now\, \$12803_loop666_arg%next\, 
         \$12803_loop666_arg%now\, \$12679_loop666_arg%next\, 
         \$12679_loop666_arg%now\, \$18632_loop666_arg%next\, 
         \$18632_loop666_arg%now\, \$17458_loop666_arg%next\, 
         \$17458_loop666_arg%now\, \$17457_aux664_arg%next\, 
         \$17457_aux664_arg%now\, \$12520_loop666_arg%next\, 
         \$12520_loop666_arg%now\, \$17455_loop666_arg%next\, 
         \$17455_loop666_arg%now\, \$13920_loop666_arg%next\, 
         \$13920_loop666_arg%now\ : value(0 to 63) := (others => '0');
  signal \$18323%next\, \$18323%now\, \$17780%next\, \$17780%now\, 
         \$17753%next\, \$17753%now\, \$13097%next\, \$13097%now\, 
         \$13124%next\, \$13124%now\, \$13791%next\, \$13791%now\, 
         \$18812%next\, \$18812%now\, \$18705%next\, \$18705%now\, 
         \$17539%next\, \$17539%now\, \$17566%next\, \$17566%now\, 
         \$19239%next\, \$19239%now\, \$12548_dis%next\, \$12548_dis%now\, 
         \$17324%next\, \$17324%now\, \$12835%next\, \$12835%now\, 
         \$18661%next\, \$18661%now\, \$13507%next\, \$13507%now\, 
         \$12818%next\, \$12818%now\, \$19115%next\, \$19115%now\, 
         \$17327%next\, \$17327%now\, \$12910%next\, \$12910%now\, 
         \$18163%next\, \$18163%now\, \$17321%next\, \$17321%now\, 
         \$17487%next\, \$17487%now\, \$13667%next\, \$13667%now\, 
         \$18644%next\, \$18644%now\, \$18447%next\, \$18447%now\, 
         \$17470%next\, \$17470%now\, \$12883%next\, \$12883%now\ : value(0 to 47) := (others => '0');
  signal \$15648_compare6445897_arg%next\, \$15648_compare6445897_arg%now\, 
         \$16846_compare6445898_arg%next\, \$16846_compare6445898_arg%now\, 
         \$15684_compare6445897_arg%next\, \$15684_compare6445897_arg%now\, 
         \$16986_compare6445898_arg%next\, \$16986_compare6445898_arg%now\, 
         \$15792_compare6445897_arg%next\, \$15792_compare6445897_arg%now\, 
         \$16612_compare6445898_arg%next\, \$16612_compare6445898_arg%now\, 
         \$16574_compare6445898_arg%next\, \$16574_compare6445898_arg%now\, 
         \$16916_compare6445898_arg%next\, \$16916_compare6445898_arg%now\, 
         \$15828_compare6445897_arg%next\, \$15828_compare6445897_arg%now\, 
         \$16881_compare6445898_arg%next\, \$16881_compare6445898_arg%now\, 
         \$15720_compare6445897_arg%next\, \$15720_compare6445897_arg%now\, 
         \$16951_compare6445898_arg%next\, \$16951_compare6445898_arg%now\, 
         \$15756_compare6445897_arg%next\, \$15756_compare6445897_arg%now\, 
         \$16811_compare6445898_arg%next\, \$16811_compare6445898_arg%now\ : value(0 to 93) := (others => '0');
  signal \$13911%next\, \$13911%now\, \$13897%next\, \$13897%now\, 
         \$13917%next\, \$13917%now\, \$13927_branch_if648_arg%next\, 
         \$13927_branch_if648_arg%now\ : value(0 to 122) := (others => '0');
  signal \$17547_copy_root_in_ram6635891_result%next\, 
         \$17547_copy_root_in_ram6635891_result%now\, \$16659_sp%next\, 
         \$16659_sp%now\, \$12840_next%next\, \$12840_next%now\, 
         \$18665%next\, \$18665%now\, \$17330_sp%next\, \$17330_sp%now\, 
         \$18793_copy_root_in_ram6635879_result%next\, 
         \$18793_copy_root_in_ram6635879_result%now\, 
         \$13105_copy_root_in_ram6635884_result%next\, 
         \$13105_copy_root_in_ram6635884_result%now\, 
         \$18686_copy_root_in_ram6635880_result%next\, 
         \$18686_copy_root_in_ram6635880_result%now\, 
         \$16662_fill6535928_result%next\, \$16662_fill6535928_result%now\, 
         \$13921_loop665_result%next\, \$13921_loop665_result%now\, 
         \$17105_w06555936_result%next\, \$17105_w06555936_result%now\, 
         \$12891_copy_root_in_ram6635884_result%next\, 
         \$12891_copy_root_in_ram6635884_result%now\, 
         \$17520_copy_root_in_ram6635893_result%next\, 
         \$17520_copy_root_in_ram6635893_result%now\, \$17331_sp%next\, 
         \$17331_sp%now\, \$17492_next%next\, \$17492_next%now\, 
         \$17459_loop665_result%next\, \$17459_loop665_result%now\, 
         \$13472_next%next\, \$13472_next%now\, \$18664_next%next\, 
         \$18664_next%now\, \$13078_copy_root_in_ram6635885_result%next\, 
         \$13078_copy_root_in_ram6635885_result%now\, \$18670_next%next\, 
         \$18670_next%now\, \$17490_next%next\, \$17490_next%now\, 
         \$18666_next%next\, \$18666_next%now\, \$17237_sp%next\, 
         \$17237_sp%now\, \$17734_copy_root_in_ram6635892_result%next\, 
         \$17734_copy_root_in_ram6635892_result%now\, 
         \$17018_w36575938_result%next\, \$17018_w36575938_result%now\, 
         \$18633_loop665_result%next\, \$18633_loop665_result%now\, 
         \$16650_sp%next\, \$16650_sp%now\, \$17332_sp%next\, 
         \$17332_sp%now\, \$12864_copy_root_in_ram6635886_result%next\, 
         \$12864_copy_root_in_ram6635886_result%now\, \$16749_sp%next\, 
         \$16749_sp%now\, \$17009_sp%next\, \$17009_sp%now\, 
         \$12804_loop665_result%next\, \$12804_loop665_result%now\, 
         \$12807_loop665_result%next\, \$12807_loop665_result%now\, 
         \$17456_loop665_result%next\, \$17456_loop665_result%now\, 
         \$16063_w6515922_result%next\, \$16063_w6515922_result%now\, 
         \$17000_sp%next\, \$17000_sp%now\, \$17460_aux664_result%next\, 
         \$17460_aux664_result%now\, \$16202_ofs%next\, \$16202_ofs%now\, 
         \$12521_loop665_result%next\, \$12521_loop665_result%now\, 
         \$18288_next%next\, \$18288_next%now\, \$16036_sp%next\, 
         \$16036_sp%now\, \$12838_next%next\, \$12838_next%now\, 
         \$17491%next\, \$17491%now\, \$12844_next%next\, \$12844_next%now\, 
         \$12680_loop665_result%next\, \$12680_loop665_result%now\, 
         \$18634_aux664_result%next\, \$18634_aux664_result%now\, 
         \$17012_sp%next\, \$17012_sp%now\, \$17333_sp%next\, 
         \$17333_sp%now\, \$17761_copy_root_in_ram6635891_result%next\, 
         \$17761_copy_root_in_ram6635891_result%now\, \$18128_next%next\, 
         \$18128_next%now\, \$14207_loop_push6495899_result%next\, 
         \$14207_loop_push6495899_result%now\, \$17238_sp%next\, 
         \$17238_sp%now\, \$14181_sp%next\, \$14181_sp%now\, 
         \$17457_aux664_result%next\, \$17457_aux664_result%now\, 
         \$12808_aux664_result%next\, \$12808_aux664_result%now\, 
         \$12805_aux664_result%next\, \$12805_aux664_result%now\, 
         \$12839%next\, \$12839%now\, \$13632_next%next\, \$13632_next%now\, 
         \$16752_fill6545929_result%next\, \$16752_fill6545929_result%now\, 
         \$19080_next%next\, \$19080_next%now\, \$17496_next%next\, 
         \$17496_next%now\ : value(0 to 15) := (others => '0');
  signal \$12563%next\, \$12563%now\, \$12558%next\, \$12558%now\, 
         \$12562%next\, \$12562%now\, \$12561%next\, \$12561%now\, 
         \$v7438%next\, \$v7438%now\, \$v7442%next\, \$v7442%now\, 
         \$v7450%next\, \$v7450%now\, \$12560%next\, \$12560%now\, 
         \$v7446%next\, \$v7446%now\, \$12559%next\, \$12559%now\ : value(0 to 7) := (others => '0');
  signal \$14613_modulo6685896_arg%next\, \$14613_modulo6685896_arg%now\, 
         \$15013_modulo6685896_arg%next\, \$15013_modulo6685896_arg%now\, 
         \$15253_modulo6685896_arg%next\, \$15253_modulo6685896_arg%now\, 
         \$14997_modulo6685888_arg%next\, \$14997_modulo6685888_arg%now\, 
         \$15149_modulo6685895_arg%next\, \$15149_modulo6685895_arg%now\, 
         \$14757_modulo6685888_arg%next\, \$14757_modulo6685888_arg%now\, 
         \$14933_modulo6685896_arg%next\, \$14933_modulo6685896_arg%now\, 
         \$15333_modulo6685896_arg%next\, \$15333_modulo6685896_arg%now\, 
         \$15556_modulo6685895_arg%next\, \$15556_modulo6685895_arg%now\, 
         \$15101_modulo6685888_arg%next\, \$15101_modulo6685888_arg%now\, 
         \$14829_modulo6685895_arg%next\, \$14829_modulo6685895_arg%now\, 
         \$15508_modulo6685888_arg%next\, \$15508_modulo6685888_arg%now\, 
         \$15588_modulo6685888_arg%next\, \$15588_modulo6685888_arg%now\, 
         \$15181_modulo6685888_arg%next\, \$15181_modulo6685888_arg%now\, 
         \$14781_modulo6685888_arg%next\, \$14781_modulo6685888_arg%now\, 
         \$15173_modulo6685896_arg%next\, \$15173_modulo6685896_arg%now\, 
         \$15077_modulo6685888_arg%next\, \$15077_modulo6685888_arg%now\, 
         \$15413_modulo6685896_arg%next\, \$15413_modulo6685896_arg%now\, 
         \$14589_modulo6685895_arg%next\, \$14589_modulo6685895_arg%now\, 
         \$14621_modulo6685888_arg%next\, \$14621_modulo6685888_arg%now\, 
         \$14861_modulo6685888_arg%next\, \$14861_modulo6685888_arg%now\, 
         \$15157_modulo6685888_arg%next\, \$15157_modulo6685888_arg%now\, 
         \$15564_modulo6685888_arg%next\, \$15564_modulo6685888_arg%now\, 
         \$14909_modulo6685895_arg%next\, \$14909_modulo6685895_arg%now\, 
         \$15421_modulo6685888_arg%next\, \$15421_modulo6685888_arg%now\, 
         \$15580_modulo6685896_arg%next\, \$15580_modulo6685896_arg%now\, 
         \$14669_modulo6685895_arg%next\, \$14669_modulo6685895_arg%now\, 
         \$15309_modulo6685895_arg%next\, \$15309_modulo6685895_arg%now\, 
         \$14941_modulo6685888_arg%next\, \$14941_modulo6685888_arg%now\, 
         \$14693_modulo6685896_arg%next\, \$14693_modulo6685896_arg%now\, 
         \$15237_modulo6685888_arg%next\, \$15237_modulo6685888_arg%now\, 
         \$15093_modulo6685896_arg%next\, \$15093_modulo6685896_arg%now\, 
         \$15341_modulo6685888_arg%next\, \$15341_modulo6685888_arg%now\, 
         \$15317_modulo6685888_arg%next\, \$15317_modulo6685888_arg%now\, 
         \$14853_modulo6685896_arg%next\, \$14853_modulo6685896_arg%now\, 
         \$14837_modulo6685888_arg%next\, \$14837_modulo6685888_arg%now\, 
         \$15484_modulo6685888_arg%next\, \$15484_modulo6685888_arg%now\, 
         \$15021_modulo6685888_arg%next\, \$15021_modulo6685888_arg%now\, 
         \$15261_modulo6685888_arg%next\, \$15261_modulo6685888_arg%now\, 
         \$15500_modulo6685896_arg%next\, \$15500_modulo6685896_arg%now\, 
         \$14773_modulo6685896_arg%next\, \$14773_modulo6685896_arg%now\, 
         \$15229_modulo6685895_arg%next\, \$15229_modulo6685895_arg%now\, 
         \$15397_modulo6685888_arg%next\, \$15397_modulo6685888_arg%now\, 
         \$14677_modulo6685888_arg%next\, \$14677_modulo6685888_arg%now\, 
         \$15476_modulo6685895_arg%next\, \$15476_modulo6685895_arg%now\, 
         \$14701_modulo6685888_arg%next\, \$14701_modulo6685888_arg%now\, 
         \$14749_modulo6685895_arg%next\, \$14749_modulo6685895_arg%now\, 
         \$15389_modulo6685895_arg%next\, \$15389_modulo6685895_arg%now\, 
         \$14597_modulo6685888_arg%next\, \$14597_modulo6685888_arg%now\, 
         \$14989_modulo6685895_arg%next\, \$14989_modulo6685895_arg%now\, 
         \$14917_modulo6685888_arg%next\, \$14917_modulo6685888_arg%now\, 
         \$15069_modulo6685895_arg%next\, \$15069_modulo6685895_arg%now\ : value(0 to 61) := (others => '0');
  signal \$13922_wait662_arg%next\, \$13922_wait662_arg%now\, 
         \$12681_wait662_arg%next\, \$12681_wait662_arg%now\, 
         \$12522_wait662_arg%next\, \$12522_wait662_arg%now\ : value(0 to 96) := (others => '0');
  signal \result5939%next\, \result5939%now\ : value(0 to 57) := (others => '0');
  signal \$12539%next\, \$12539%now\, \$v6107%next\, \$v6107%now\, 
         \$12662%next\, \$12662%now\, \$v6106%next\, \$v6106%now\, 
         \$v6104%next\, \$v6104%now\, \$v6103%next\, \$v6103%now\, 
         \$v6108%next\, \$v6108%now\, \$v6105%next\, \$v6105%now\ : value(0 to 3) := (others => '0');
  signal \$15508_modulo6685888_id%next\, \$15508_modulo6685888_id%now\, 
         \$13925_offsetclosure_n639_id%next\, 
         \$13925_offsetclosure_n639_id%now\, \$15229_modulo6685895_id%next\, 
         \$15229_modulo6685895_id%now\, \$15013_modulo6685896_id%next\, 
         \$15013_modulo6685896_id%now\, 
         \$15697_binop_compare6455918_id%next\, 
         \$15697_binop_compare6455918_id%now\, 
         \$14207_loop_push6495899_id%next\, \$14207_loop_push6495899_id%now\, 
         \$13923_make_block579_id%next\, \$13923_make_block579_id%now\, 
         \$17456_loop665_id%next\, \$17456_loop665_id%now\, 
         \$15805_binop_compare6455921_id%next\, 
         \$15805_binop_compare6455921_id%now\, 
         \$14884_binop_int6435904_id%next\, \$14884_binop_int6435904_id%now\, 
         \$15564_modulo6685888_id%next\, \$15564_modulo6685888_id%now\, 
         \$15451_binop_int6435912_id%next\, \$15451_binop_int6435912_id%now\, 
         \$15317_modulo6685888_id%next\, \$15317_modulo6685888_id%now\, 
         \$15588_modulo6685888_id%next\, \$15588_modulo6685888_id%now\, 
         \$16951_compare6445898_id%next\, \$16951_compare6445898_id%now\, 
         \$15733_binop_compare6455919_id%next\, 
         \$15733_binop_compare6455919_id%now\, 
         \$14941_modulo6685888_id%next\, \$14941_modulo6685888_id%now\, 
         \$14621_modulo6685888_id%next\, \$14621_modulo6685888_id%now\, 
         \$14853_modulo6685896_id%next\, \$14853_modulo6685896_id%now\, 
         \$15621_forever6705915_id%next\, \$15621_forever6705915_id%now\, 
         \$15756_compare6445897_id%next\, \$15756_compare6445897_id%now\, 
         \$16788_compbranch6505930_id%next\, 
         \$16788_compbranch6505930_id%now\, \$14589_modulo6685895_id%next\, 
         \$14589_modulo6685895_id%now\, \$14781_modulo6685888_id%next\, 
         \$14781_modulo6685888_id%now\, \$14701_modulo6685888_id%next\, 
         \$14701_modulo6685888_id%now\, \$13924_apply638_id%next\, 
         \$13924_apply638_id%now\, \$15309_modulo6685895_id%next\, 
         \$15309_modulo6685895_id%now\, \$15181_modulo6685888_id%next\, 
         \$15181_modulo6685888_id%now\, 
         \$12891_copy_root_in_ram6635884_id%next\, 
         \$12891_copy_root_in_ram6635884_id%now\, 
         \$15556_modulo6685895_id%next\, \$15556_modulo6685895_id%now\, 
         \$17459_loop665_id%next\, \$17459_loop665_id%now\, 
         \$15500_modulo6685896_id%next\, \$15500_modulo6685896_id%now\, 
         \$15093_modulo6685896_id%next\, \$15093_modulo6685896_id%now\, 
         \$17048_w16565937_id%next\, \$17048_w16565937_id%now\, 
         \$13927_branch_if648_id%next\, \$13927_branch_if648_id%now\, 
         \$16662_fill6535928_id%next\, \$16662_fill6535928_id%now\, 
         \$16811_compare6445898_id%next\, \$16811_compare6445898_id%now\, 
         \$18634_aux664_id%next\, \$18634_aux664_id%now\, 
         \$17505_forever6705894_id%next\, \$17505_forever6705894_id%now\, 
         \$12857_forever6705883_id%next\, \$12857_forever6705883_id%now\, 
         \$15413_modulo6685896_id%next\, \$15413_modulo6685896_id%now\, 
         \$18632_loop666_id%next\, \$18632_loop666_id%now\, 
         \$13105_copy_root_in_ram6635884_id%next\, 
         \$13105_copy_root_in_ram6635884_id%now\, 
         \$15021_modulo6685888_id%next\, \$15021_modulo6685888_id%now\, 
         \$16752_fill6545929_id%next\, \$16752_fill6545929_id%now\, 
         \$15684_compare6445897_id%next\, \$15684_compare6445897_id%now\, 
         \$14597_modulo6685888_id%next\, \$14597_modulo6685888_id%now\, 
         \$14644_binop_int6435901_id%next\, \$14644_binop_int6435901_id%now\, 
         \$16881_compare6445898_id%next\, \$16881_compare6445898_id%now\, 
         \$15792_compare6445897_id%next\, \$15792_compare6445897_id%now\, 
         \$16858_compbranch6505932_id%next\, 
         \$16858_compbranch6505932_id%now\, \$12803_loop666_id%next\, 
         \$12803_loop666_id%now\, \$15614_forever6705914_id%next\, 
         \$15614_forever6705914_id%now\, \$14693_modulo6685896_id%next\, 
         \$14693_modulo6685896_id%now\, \$15397_modulo6685888_id%next\, 
         \$15397_modulo6685888_id%now\, \$12804_loop665_id%next\, 
         \$12804_loop665_id%now\, \$15661_binop_compare6455917_id%next\, 
         \$15661_binop_compare6455917_id%now\, 
         \$16612_compare6445898_id%next\, \$16612_compare6445898_id%now\, 
         \$15149_modulo6685895_id%next\, \$15149_modulo6685895_id%now\, 
         \$18793_copy_root_in_ram6635879_id%next\, 
         \$18793_copy_root_in_ram6635879_id%now\, \$12522_wait662_id%next\, 
         \$12522_wait662_id%now\, \$14989_modulo6685895_id%next\, 
         \$14989_modulo6685895_id%now\, \$15173_modulo6685896_id%next\, 
         \$15173_modulo6685896_id%now\, \$14804_binop_int6435903_id%next\, 
         \$14804_binop_int6435903_id%now\, \$12681_wait662_id%next\, 
         \$12681_wait662_id%now\, \$13928_w652_id%next\, 
         \$13928_w652_id%now\, \$17509_forever6705890_id%next\, 
         \$17509_forever6705890_id%now\, \$15333_modulo6685896_id%next\, 
         \$15333_modulo6685896_id%now\, \$16986_compare6445898_id%next\, 
         \$16986_compare6445898_id%now\, \$12853_forever6705887_id%next\, 
         \$12853_forever6705887_id%now\, \$14861_modulo6685888_id%next\, 
         \$14861_modulo6685888_id%now\, \$13920_loop666_id%next\, 
         \$13920_loop666_id%now\, \$14564_binop_int6435900_id%next\, 
         \$14564_binop_int6435900_id%now\, \$17458_loop666_id%next\, 
         \$17458_loop666_id%now\, \$15077_modulo6685888_id%next\, 
         \$15077_modulo6685888_id%now\, \$15447_forever6705911_id%next\, 
         \$15447_forever6705911_id%now\, \$15157_modulo6685888_id%next\, 
         \$15157_modulo6685888_id%now\, 
         \$17547_copy_root_in_ram6635891_id%next\, 
         \$17547_copy_root_in_ram6635891_id%now\, 
         \$14909_modulo6685895_id%next\, \$14909_modulo6685895_id%now\, 
         \$13926_make_block_n646_id%next\, \$13926_make_block_n646_id%now\, 
         \$16846_compare6445898_id%next\, \$16846_compare6445898_id%now\, 
         \$12864_copy_root_in_ram6635886_id%next\, 
         \$12864_copy_root_in_ram6635886_id%now\, 
         \$14757_modulo6685888_id%next\, \$14757_modulo6685888_id%now\, 
         \$14773_modulo6685896_id%next\, \$14773_modulo6685896_id%now\, 
         \$15389_modulo6685895_id%next\, \$15389_modulo6685895_id%now\, 
         \$16928_compbranch6505934_id%next\, 
         \$16928_compbranch6505934_id%now\, 
         \$18686_copy_root_in_ram6635880_id%next\, 
         \$18686_copy_root_in_ram6635880_id%now\, \$16063_w6515922_id%next\, 
         \$16063_w6515922_id%now\, \$13922_wait662_id%next\, 
         \$13922_wait662_id%now\, \$15101_modulo6685888_id%next\, 
         \$15101_modulo6685888_id%now\, \$16158_forever6705923_id%next\, 
         \$16158_forever6705923_id%now\, \$14837_modulo6685888_id%next\, 
         \$14837_modulo6685888_id%now\, \$15364_binop_int6435910_id%next\, 
         \$15364_binop_int6435910_id%now\, \$15284_binop_int6435909_id%next\, 
         \$15284_binop_int6435909_id%now\, \$15531_binop_int6435913_id%next\, 
         \$15531_binop_int6435913_id%now\, \$16195_forever6705924_id%next\, 
         \$16195_forever6705924_id%now\, \$16916_compare6445898_id%next\, 
         \$16916_compare6445898_id%now\, \$15421_modulo6685888_id%next\, 
         \$15421_modulo6685888_id%now\, \$14917_modulo6685888_id%next\, 
         \$14917_modulo6685888_id%now\, \$12806_loop666_id%next\, 
         \$12806_loop666_id%now\, \$15253_modulo6685896_id%next\, 
         \$15253_modulo6685896_id%now\, \$15341_modulo6685888_id%next\, 
         \$15341_modulo6685888_id%now\, \$15580_modulo6685896_id%next\, 
         \$15580_modulo6685896_id%now\, \$15476_modulo6685895_id%next\, 
         \$15476_modulo6685895_id%now\, 
         \$17761_copy_root_in_ram6635891_id%next\, 
         \$17761_copy_root_in_ram6635891_id%now\, 
         \$16823_compbranch6505931_id%next\, 
         \$16823_compbranch6505931_id%now\, 
         \$15769_binop_compare6455920_id%next\, 
         \$15769_binop_compare6455920_id%now\, 
         \$15828_compare6445897_id%next\, \$15828_compare6445897_id%now\, 
         \$14669_modulo6685895_id%next\, \$14669_modulo6685895_id%now\, 
         \$13078_copy_root_in_ram6635885_id%next\, 
         \$13078_copy_root_in_ram6635885_id%now\, 
         \$14613_modulo6685896_id%next\, \$14613_modulo6685896_id%now\, 
         \$15648_compare6445897_id%next\, \$15648_compare6445897_id%now\, 
         \$14964_binop_int6435905_id%next\, \$14964_binop_int6435905_id%now\, 
         \$17513_forever6705889_id%next\, \$17513_forever6705889_id%now\, 
         \$15204_binop_int6435908_id%next\, \$15204_binop_int6435908_id%now\, 
         \$17018_w36575938_id%next\, \$17018_w36575938_id%now\, 
         \$17520_copy_root_in_ram6635893_id%next\, 
         \$17520_copy_root_in_ram6635893_id%now\, 
         \$15484_modulo6685888_id%next\, \$15484_modulo6685888_id%now\, 
         \$14933_modulo6685896_id%next\, \$14933_modulo6685896_id%now\, 
         \$14724_binop_int6435902_id%next\, \$14724_binop_int6435902_id%now\, 
         \$14749_modulo6685895_id%next\, \$14749_modulo6685895_id%now\, 
         \$12679_loop666_id%next\, \$12679_loop666_id%now\, 
         \$17105_w06555936_id%next\, \$17105_w06555936_id%now\, 
         \$15069_modulo6685895_id%next\, \$15069_modulo6685895_id%now\, 
         \$12807_loop665_id%next\, \$12807_loop665_id%now\, 
         \$17460_aux664_id%next\, \$17460_aux664_id%now\, 
         \$16510_forever6705925_id%next\, \$16510_forever6705925_id%now\, 
         \$16589_compbranch6505927_id%next\, 
         \$16589_compbranch6505927_id%now\, \$12808_aux664_id%next\, 
         \$12808_aux664_id%now\, \$15720_compare6445897_id%next\, 
         \$15720_compare6445897_id%now\, \$18679_forever6705881_id%next\, 
         \$18679_forever6705881_id%now\, \$15237_modulo6685888_id%next\, 
         \$15237_modulo6685888_id%now\, \$14677_modulo6685888_id%next\, 
         \$14677_modulo6685888_id%now\, \$14829_modulo6685895_id%next\, 
         \$14829_modulo6685895_id%now\, 
         \$15625_binop_compare6455916_id%next\, 
         \$15625_binop_compare6455916_id%now\, \$18633_loop665_id%next\, 
         \$18633_loop665_id%now\, \$15124_binop_int6435907_id%next\, 
         \$15124_binop_int6435907_id%now\, 
         \$16551_compbranch6505926_id%next\, 
         \$16551_compbranch6505926_id%now\, \$12520_loop666_id%next\, 
         \$12520_loop666_id%now\, \$16963_compbranch6505935_id%next\, 
         \$16963_compbranch6505935_id%now\, 
         \$15044_binop_int6435906_id%next\, \$15044_binop_int6435906_id%now\, 
         \$16574_compare6445898_id%next\, \$16574_compare6445898_id%now\, 
         \$17455_loop666_id%next\, \$17455_loop666_id%now\, 
         \$17734_copy_root_in_ram6635892_id%next\, 
         \$17734_copy_root_in_ram6635892_id%now\, 
         \$15261_modulo6685888_id%next\, \$15261_modulo6685888_id%now\, 
         \$14997_modulo6685888_id%next\, \$14997_modulo6685888_id%now\, 
         \$16893_compbranch6505933_id%next\, 
         \$16893_compbranch6505933_id%now\ : value(0 to 11) := (others => '0');
  signal \$16893_compbranch6505933_arg%next\, 
         \$16893_compbranch6505933_arg%now\, 
         \$16928_compbranch6505934_arg%next\, 
         \$16928_compbranch6505934_arg%now\, 
         \$16589_compbranch6505927_arg%next\, 
         \$16589_compbranch6505927_arg%now\, 
         \$16551_compbranch6505926_arg%next\, 
         \$16551_compbranch6505926_arg%now\, 
         \$16963_compbranch6505935_arg%next\, 
         \$16963_compbranch6505935_arg%now\, 
         \$16823_compbranch6505931_arg%next\, 
         \$16823_compbranch6505931_arg%now\, 
         \$16788_compbranch6505930_arg%next\, 
         \$16788_compbranch6505930_arg%now\, 
         \$16858_compbranch6505932_arg%next\, 
         \$16858_compbranch6505932_arg%now\ : value(0 to 215) := (others => '0');
  signal \$14690_r%next\, \$14690_r%now\, \$14770_r%next\, \$14770_r%now\, 
         \$14662_res%next\, \$14662_res%now\, \$15226_r%next\, 
         \$15226_r%now\, \$14822_res%next\, \$14822_res%now\, 
         \$15549_res%next\, \$15549_res%now\, \$17062%next\, \$17062%now\, 
         \$15146_r%next\, \$15146_r%now\, \$14850_r%next\, \$14850_r%now\, 
         \$15157_modulo6685888_result%next\, 
         \$15157_modulo6685888_result%now\, \$15066_r%next\, \$15066_r%now\, 
         \$14586_r%next\, \$14586_r%now\, \$14742_res%next\, 
         \$14742_res%now\, \$v7329%next\, \$v7329%now\, \$15469_res%next\, 
         \$15469_res%now\, \$15222_res%next\, \$15222_res%now\, 
         \$15149_modulo6685895_result%next\, 
         \$15149_modulo6685895_result%now\, \$14906_r%next\, \$14906_r%now\, 
         \$15090_r%next\, \$15090_r%now\, \$15473_r%next\, \$15473_r%now\, 
         \$15093_modulo6685896_result%next\, 
         \$15093_modulo6685896_result%now\, \$13965%next\, \$13965%now\, 
         \$15013_modulo6685896_result%next\, 
         \$15013_modulo6685896_result%now\, \$16998_argument3%next\, 
         \$16998_argument3%now\, \$14982_res%next\, \$14982_res%now\, 
         \$15069_modulo6685895_result%next\, 
         \$15069_modulo6685895_result%now\, \$16624_argument2%next\, 
         \$16624_argument2%now\, \$14669_modulo6685895_result%next\, 
         \$14669_modulo6685895_result%now\, \$15851_argument1%next\, 
         \$15851_argument1%now\, \$15142_res%next\, \$15142_res%now\, 
         \$15062_res%next\, \$15062_res%now\, \$15410_r%next\, 
         \$15410_r%now\, \$17207_arg%next\, \$17207_arg%now\, 
         \$15497_r%next\, \$15497_r%now\, \$14693_modulo6685896_result%next\, 
         \$14693_modulo6685896_result%now\, 
         \$14917_modulo6685888_result%next\, 
         \$14917_modulo6685888_result%now\, \$15306_r%next\, \$15306_r%now\, 
         \$15173_modulo6685896_result%next\, 
         \$15173_modulo6685896_result%now\, \$14826_r%next\, \$14826_r%now\, 
         \$14853_modulo6685896_result%next\, 
         \$14853_modulo6685896_result%now\, 
         \$15421_modulo6685888_result%next\, 
         \$15421_modulo6685888_result%now\, 
         \$14997_modulo6685888_result%next\, 
         \$14997_modulo6685888_result%now\, \$15250_r%next\, \$15250_r%now\, 
         \$15588_modulo6685888_result%next\, 
         \$15588_modulo6685888_result%now\, 
         \$14773_modulo6685896_result%next\, 
         \$14773_modulo6685896_result%now\, \$15302_res%next\, 
         \$15302_res%now\, \$15170_r%next\, \$15170_r%now\, 
         \$14902_res%next\, \$14902_res%now\, 
         \$14701_modulo6685888_result%next\, 
         \$14701_modulo6685888_result%now\, \$15577_r%next\, \$15577_r%now\, 
         \$15564_modulo6685888_result%next\, 
         \$15564_modulo6685888_result%now\, 
         \$14989_modulo6685895_result%next\, 
         \$14989_modulo6685895_result%now\, 
         \$15229_modulo6685895_result%next\, 
         \$15229_modulo6685895_result%now\, \$16203%next\, \$16203%now\, 
         \$15508_modulo6685888_result%next\, 
         \$15508_modulo6685888_result%now\, 
         \$15500_modulo6685896_result%next\, 
         \$15500_modulo6685896_result%now\, 
         \$14909_modulo6685895_result%next\, 
         \$14909_modulo6685895_result%now\, 
         \$14941_modulo6685888_result%next\, 
         \$14941_modulo6685888_result%now\, 
         \$15261_modulo6685888_result%next\, 
         \$15261_modulo6685888_result%now\, \$14610_r%next\, \$14610_r%now\, 
         \$15580_modulo6685896_result%next\, 
         \$15580_modulo6685896_result%now\, 
         \$14757_modulo6685888_result%next\, 
         \$14757_modulo6685888_result%now\, 
         \$15253_modulo6685896_result%next\, 
         \$15253_modulo6685896_result%now\, 
         \$14621_modulo6685888_result%next\, 
         \$14621_modulo6685888_result%now\, \$14930_r%next\, \$14930_r%now\, 
         \$v7283%next\, \$v7283%now\, \$15309_modulo6685895_result%next\, 
         \$15309_modulo6685895_result%now\, \$17165%next\, \$17165%now\, 
         \$15382_res%next\, \$15382_res%now\, 
         \$14677_modulo6685888_result%next\, 
         \$14677_modulo6685888_result%now\, 
         \$15341_modulo6685888_result%next\, 
         \$15341_modulo6685888_result%now\, 
         \$15556_modulo6685895_result%next\, 
         \$15556_modulo6685895_result%now\, \$14746_r%next\, \$14746_r%now\, 
         \$15413_modulo6685896_result%next\, 
         \$15413_modulo6685896_result%now\, 
         \$14829_modulo6685895_result%next\, 
         \$14829_modulo6685895_result%now\, \$15010_r%next\, \$15010_r%now\, 
         \$14933_modulo6685896_result%next\, 
         \$14933_modulo6685896_result%now\, \$14986_r%next\, \$14986_r%now\, 
         \$15181_modulo6685888_result%next\, 
         \$15181_modulo6685888_result%now\, 
         \$15333_modulo6685896_result%next\, 
         \$15333_modulo6685896_result%now\, 
         \$15101_modulo6685888_result%next\, 
         \$15101_modulo6685888_result%now\, 
         \$15317_modulo6685888_result%next\, 
         \$15317_modulo6685888_result%now\, \$15386_r%next\, \$15386_r%now\, 
         \$v7290%next\, \$v7290%now\, \$15476_modulo6685895_result%next\, 
         \$15476_modulo6685895_result%now\, 
         \$15021_modulo6685888_result%next\, 
         \$15021_modulo6685888_result%now\, \$14582_res%next\, 
         \$14582_res%now\, \$14597_modulo6685888_result%next\, 
         \$14597_modulo6685888_result%now\, 
         \$14837_modulo6685888_result%next\, 
         \$14837_modulo6685888_result%now\, 
         \$15389_modulo6685895_result%next\, 
         \$15389_modulo6685895_result%now\, \$v7300%next\, \$v7300%now\, 
         \$15397_modulo6685888_result%next\, 
         \$15397_modulo6685888_result%now\, \$15330_r%next\, \$15330_r%now\, 
         \$14861_modulo6685888_result%next\, 
         \$14861_modulo6685888_result%now\, 
         \$14781_modulo6685888_result%next\, 
         \$14781_modulo6685888_result%now\, 
         \$14613_modulo6685896_result%next\, 
         \$14613_modulo6685896_result%now\, 
         \$15237_modulo6685888_result%next\, 
         \$15237_modulo6685888_result%now\, \$15553_r%next\, \$15553_r%now\, 
         \$15484_modulo6685888_result%next\, 
         \$15484_modulo6685888_result%now\, \$v7313%next\, \$v7313%now\, 
         \$14749_modulo6685895_result%next\, 
         \$14749_modulo6685895_result%now\, 
         \$15077_modulo6685888_result%next\, 
         \$15077_modulo6685888_result%now\, 
         \$14589_modulo6685895_result%next\, 
         \$14589_modulo6685895_result%now\, \$14666_r%next\, \$14666_r%now\ : value(0 to 30) := (others => '0');
  signal \$13925_offsetclosure_n639_arg%next\, 
         \$13925_offsetclosure_n639_arg%now\ : value(0 to 137) := (others => '0');
  signal \$13923_make_block579_arg%next\, \$13923_make_block579_arg%now\ : value(0 to 103) := (others => '0');
  signal \result6147%next\, \result6147%now\, \result5974%next\, 
         \result5974%now\, \$12523_make_block579_arg%next\, 
         \$12523_make_block579_arg%now\, \result6503%next\, \result6503%now\, 
         \$12682_make_block579_arg%next\, \$12682_make_block579_arg%now\ : value(0 to 127) := (others => '0');
  signal \$code_lock%next\, \$code_lock%now\, \$global_end_lock%next\, 
         \$global_end_lock%now\, \$ram_lock%next\, \$ram_lock%now\, 
         \$v6311%next\, \$v6311%now\, \$v7071%next\, \$v7071%now\, 
         \$13537%next\, \$13537%now\, \$15751_res%next\, \$15751_res%now\, 
         \$17784%next\, \$17784%now\, \$12718%next\, \$12718%now\, 
         \$14368%next\, \$14368%now\, \$v6028%next\, \$v6028%now\, 
         \$12812%next\, \$12812%now\, \$13465%next\, \$13465%now\, 
         \$v6349%next\, \$v6349%now\, \$13690%next\, \$13690%now\, 
         \$v5971%next\, \$v5971%now\, \$17965%next\, \$17965%now\, 
         \$v6010%next\, \$v6010%now\, \$v6592%next\, \$v6592%now\, 
         \$v6932%next\, \$v6932%now\, \$13020%next\, \$13020%now\, 
         \$12690%next\, \$12690%now\, \$v7316%next\, \$v7316%now\, 
         \$13128%next\, \$13128%now\, \$v7209%next\, \$v7209%now\, 
         \$17236%next\, \$17236%now\, \$v7239%next\, \$v7239%now\, 
         \$v7053%next\, \$v7053%now\, \$v6168%next\, \$v6168%now\, 
         \$17810%next\, \$17810%now\, \$v6120%next\, \$v6120%now\, 
         \$v6063%next\, \$v6063%now\, \$v6636%next\, \$v6636%now\, 
         \$v7312%next\, \$v7312%now\, \$14355%next\, \$14355%now\, 
         \$13622%next\, \$13622%now\, \$v7063%next\, \$v7063%now\, 
         \$v7384%next\, \$v7384%now\, \$v7124%next\, \$v7124%now\, 
         \$v6630%next\, \$v6630%now\, \$12661%next\, \$12661%now\, 
         \$v6687%next\, \$v6687%now\, \$18656%next\, \$18656%now\, 
         \$12876%next\, \$12876%now\, \$v6944%next\, \$v6944%now\, 
         \$13699%next\, \$13699%now\, \$v6674%next\, \$v6674%now\, 
         \$v6923%next\, \$v6923%now\, \$v7225%next\, \$v7225%now\, 
         \$18477%next\, \$18477%now\, \$12850%next\, \$12850%now\, 
         \$v7043%next\, \$v7043%now\, \$16910_b%next\, \$16910_b%now\, 
         \$v6929%next\, \$v6929%now\, \$v7152%next\, \$v7152%now\, 
         \$13534%next\, \$13534%now\, \$v7286%next\, \$v7286%now\, 
         \$18469%next\, \$18469%now\, \$19056%next\, \$19056%now\, 
         \$13230%next\, \$13230%now\, \$13305%next\, \$13305%now\, 
         \$v6612%next\, \$v6612%now\, \$17806%next\, \$17806%now\, 
         \$17396%next\, \$17396%now\, \$v7319%next\, \$v7319%now\, 
         \$v6226%next\, \$v6226%now\, \$v7065%next\, \$v7065%now\, 
         \$17161%next\, \$17161%now\, \$18923%next\, \$18923%now\, 
         \$19137%next\, \$19137%now\, \$15444%next\, \$15444%now\, 
         \$18422%next\, \$18422%now\, \$18632_loop666_result%next\, 
         \$18632_loop666_result%now\, \$v7148%next\, \$v7148%now\, 
         \$18840%next\, \$18840%now\, \$18847%next\, \$18847%now\, 
         \$14561%next\, \$14561%now\, \$v7073%next\, \$v7073%now\, 
         \$v7173%next\, \$v7173%now\, \$12940%next\, \$12940%now\, 
         \$v6777%next\, \$v6777%now\, \$18700%next\, \$18700%now\, 
         \$18347%next\, \$18347%now\, \$v7394%next\, \$v7394%now\, 
         \$v6615%next\, \$v6615%now\, \$v7325%next\, \$v7325%now\, 
         \$13819%next\, \$13819%now\, \$v6483%next\, \$v6483%now\, 
         \$v5864%next\, \$v5864%now\, \$12711%next\, \$12711%now\, 
         \$v6310%next\, \$v6310%now\, \$17601%next\, \$17601%now\, 
         \$18282%next\, \$18282%now\, \$18920%next\, \$18920%now\, 
         \$12721%next\, \$12721%now\, \$v6210%next\, \$v6210%now\, 
         \$16951_compare6445898_result%next\, 
         \$16951_compare6445898_result%now\, \$12700%next\, \$12700%now\, 
         \$v6877%next\, \$v6877%now\, \$15446%next\, \$15446%now\, 
         \$v6145%next\, \$v6145%now\, \$v6086%next\, \$v6086%now\, 
         \$13391%next\, \$13391%now\, \$v6141%next\, \$v6141%now\, 
         \$17756%next\, \$17756%now\, \$17352%next\, \$17352%now\, 
         \$v7052%next\, \$v7052%now\, \$16358%next\, \$16358%now\, 
         \$v6018%next\, \$v6018%now\, \$17757%next\, \$17757%now\, 
         \$17571%next\, \$17571%now\, \$13448%next\, \$13448%now\, 
         \$18039%next\, \$18039%now\, \$v6977%next\, \$v6977%now\, 
         \$13014%next\, \$13014%now\, \$18349%next\, \$18349%now\, 
         \$16980_b%next\, \$16980_b%now\, \$17811%next\, \$17811%now\, 
         \$v6540%next\, \$v6540%now\, \$18195%next\, \$18195%now\, 
         \$14015%next\, \$14015%now\, \$19072%next\, \$19072%now\, 
         \$19148%next\, \$19148%now\, \$17672%next\, \$17672%now\, 
         \$v6871%next\, \$v6871%now\, \$18817%next\, \$18817%now\, 
         \$16846_compare6445898_result%next\, 
         \$16846_compare6445898_result%now\, \$18914%next\, \$18914%now\, 
         \$15643_res%next\, \$15643_res%now\, \$v7309%next\, \$v7309%now\, 
         \$14260%next\, \$14260%now\, \$17483%next\, \$17483%now\, 
         \$v7055%next\, \$v7055%now\, \$16357%next\, \$16357%now\, 
         \$18350%next\, \$18350%now\, \$v7266%next\, \$v7266%now\, 
         \$v6793%next\, \$v6793%now\, \$18471%next\, \$18471%now\, 
         \$13130%next\, \$13130%now\, \$v6024%next\, \$v6024%now\, 
         \$13231%next\, \$13231%now\, \$v5877%next\, \$v5877%now\, 
         \$19000%next\, \$19000%now\, \$18468%next\, \$18468%now\, 
         \$v7001%next\, \$v7001%now\, \$16296%next\, \$16296%now\, 
         \$16706%next\, \$16706%now\, \$19141%next\, \$19141%now\, 
         \$16413%next\, \$16413%now\, \$17596%next\, \$17596%now\, 
         \$15620%next\, \$15620%now\, \$19073%next\, \$19073%now\, 
         \$v6006%next\, \$v6006%now\, \$v5979%next\, \$v5979%now\, 
         \$18710%next\, \$18710%now\, \$v6808%next\, \$v6808%now\, 
         \$15611%next\, \$15611%now\, \$v6039%next\, \$v6039%now\, 
         \$13015%next\, \$13015%now\, \$13953%next\, \$13953%now\, 
         \$13159%next\, \$13159%now\, \$16293%next\, \$16293%now\, 
         \$13920_loop666_result%next\, \$13920_loop666_result%now\, 
         \$v7106%next\, \$v7106%now\, \$12693%next\, \$12693%now\, 
         \$16155%next\, \$16155%now\, \$13152%next\, \$13152%now\, 
         \$v6486%next\, \$v6486%now\, \$v6191%next\, \$v6191%now\, 
         \$17680%next\, \$17680%now\, \$v7040%next\, \$v7040%now\, 
         \$v6770%next\, \$v6770%now\, \$v6886%next\, \$v6886%now\, 
         \$v6051%next\, \$v6051%now\, \$v6250%next\, \$v6250%now\, 
         \$v6418%next\, \$v6418%now\, \$v6671%next\, \$v6671%now\, 
         \$v7430%next\, \$v7430%now\, \$v6850%next\, \$v6850%now\, 
         \$19270%next\, \$19270%now\, \$13462%next\, \$13462%now\, 
         \$v7341%next\, \$v7341%now\, \$v6539%next\, \$v6539%now\, 
         \$13306%next\, \$13306%now\, \$v7390%next\, \$v7390%now\, 
         \$v7131%next\, \$v7131%now\, \$v7410%next\, \$v7410%now\, 
         \$v6331%next\, \$v6331%now\, \$17486%next\, \$17486%now\, 
         \$v6339%next\, \$v6339%now\, \$v5968%next\, \$v5968%now\, 
         \$v7136%next\, \$v7136%now\, \$16658%next\, \$16658%now\, 
         \$12831%next\, \$12831%now\, \$v6747%next\, \$v6747%now\, 
         \$v7407%next\, \$v7407%now\, \$v6412%next\, \$v6412%now\, 
         \$17061%next\, \$17061%now\, \$12687%next\, \$12687%now\, 
         \$v6556%next\, \$v6556%now\, \$13952%next\, \$13952%now\, 
         \$v6497%next\, \$v6497%now\, \$v7160%next\, \$v7160%now\, 
         \$15720_compare6445897_result%next\, 
         \$15720_compare6445897_result%now\, \$v6215%next\, \$v6215%now\, 
         \$17481%next\, \$17481%now\, \$v6124%next\, \$v6124%now\, 
         \$18573%next\, \$18573%now\, \$13024%next\, \$13024%now\, 
         \$v7075%next\, \$v7075%now\, \$v6698%next\, \$v6698%now\, 
         \$v7026%next\, \$v7026%now\, \$15908%next\, \$15908%now\, 
         \$v6076%next\, \$v6076%now\, \$18042%next\, \$18042%now\, 
         \$v7270%next\, \$v7270%now\, \rdy5975%next\, \rdy5975%now\, 
         \$v6260%next\, \$v6260%now\, \$19074%next\, \$19074%now\, 
         \$18672%next\, \$18672%now\, \$v6032%next\, \$v6032%now\, 
         \$13118%next\, \$13118%now\, \$v6663%next\, \$v6663%now\, 
         \$v7257%next\, \$v7257%now\, \$v6983%next\, \$v6983%now\, 
         \$17353%next\, \$17353%now\, \$v6620%next\, \$v6620%now\, 
         \$15648_compare6445897_result%next\, 
         \$15648_compare6445897_result%now\, \$v7024%next\, \$v7024%now\, 
         \$13951%next\, \$13951%now\, \$13119%next\, \$13119%now\, 
         \$12742%next\, \$12742%now\, \$v6244%next\, \$v6244%now\, 
         \$12916%next\, \$12916%now\, \$14265%next\, \$14265%now\, 
         \$16462%next\, \$16462%now\, \$13091%next\, \$13091%now\, 
         \$v6647%next\, \$v6647%now\, \$16157%next\, \$16157%now\, 
         \$18728%next\, \$18728%now\, \$v7423%next\, \$v7423%now\, 
         \$v6576%next\, \$v6576%now\, \$v6675%next\, \$v6675%now\, 
         \$v7080%next\, \$v7080%now\, \$v6566%next\, \$v6566%now\, 
         \$13698%next\, \$13698%now\, \$v7105%next\, \$v7105%now\, 
         \$16322%next\, \$16322%now\, \$13958%next\, \$13958%now\, 
         \$v5871%next\, \$v5871%now\, \$19338%next\, \$19338%now\, 
         \$13394%next\, \$13394%now\, \$17172%next\, \$17172%now\, 
         \$v6290%next\, \$v6290%now\, \$13821%next\, \$13821%now\, 
         \$v6220%next\, \$v6220%now\, \$17807%next\, \$17807%now\, 
         \$v7226%next\, \$v7226%now\, \$18671%next\, \$18671%now\, 
         \$18736%next\, \$18736%now\, \$v7122%next\, \$v7122%now\, 
         \$18345%next\, \$18345%now\, \$13017%next\, \$13017%now\, 
         \$17589%next\, \$17589%now\, \$16195_forever6705924_arg%next\, 
         \$16195_forever6705924_arg%now\, \$v6895%next\, \$v6895%now\, 
         \$v7347%next\, \$v7347%now\, \$18353%next\, \$18353%now\, 
         \$17884%next\, \$17884%now\, \$15621_forever6705915_arg%next\, 
         \$15621_forever6705915_arg%now\, \$v6079%next\, \$v6079%now\, 
         \$v6439%next\, \$v6439%now\, \$v6571%next\, \$v6571%now\, 
         \$v6194%next\, \$v6194%now\, \$v6345%next\, \$v6345%now\, 
         \$17542%next\, \$17542%now\, \rdy6113%next\, \rdy6113%now\, 
         \$13314%next\, \$13314%now\, \$19147%next\, \$19147%now\, 
         \$v5989%next\, \$v5989%now\, \$v6926%next\, \$v6926%now\, 
         \$17534%next\, \$17534%now\, \$v6980%next\, \$v6980%now\, 
         \$17599%next\, \$17599%now\, \$13813%next\, \$13813%now\, 
         \$18589%next\, \$18589%now\, \$17533%next\, \$17533%now\, 
         \$v6755%next\, \$v6755%now\, \$v7036%next\, \$v7036%now\, 
         \$19139%next\, \$19139%now\, \$13228%next\, \$13228%now\, 
         \$17184%next\, \$17184%now\, \$v6448%next\, \$v6448%now\, 
         \$v6524%next\, \$v6524%now\, \$16724%next\, \$16724%now\, 
         \$v6083%next\, \$v6083%now\, \$v6528%next\, \$v6528%now\, 
         \$v6720%next\, \$v6720%now\, \$v6762%next\, \$v6762%now\, 
         \$13022%next\, \$13022%now\, \$v6811%next\, \$v6811%now\, 
         \$v6774%next\, \$v6774%now\, \$16461%next\, \$16461%now\, 
         \$18678%next\, \$18678%now\, \$13025%next\, \$13025%now\, 
         \$v6477%next\, \$v6477%now\, \$17465%next\, \$17465%now\, 
         \$13386%next\, \$13386%now\, \$18658%next\, \$18658%now\, 
         \$v6267%next\, \$v6267%now\, \$12905%next\, \$12905%now\, 
         \$19146%next\, \$19146%now\, \$v7303%next\, \$v7303%now\, 
         \$18839%next\, \$18839%now\, \$16916_compare6445898_result%next\, 
         \$16916_compare6445898_result%now\, \$16193%next\, \$16193%now\, 
         \$v7130%next\, \$v7130%now\, \$12657%next\, \$12657%now\, 
         \$v6691%next\, \$v6691%now\, \$14342%next\, \$14342%now\, 
         \$v6264%next\, \$v6264%now\, \$v6600%next\, \$v6600%now\, 
         \$v6582%next\, \$v6582%now\, \$17545%next\, \$17545%now\, 
         \$v6361%next\, \$v6361%now\, \$12845%next\, \$12845%now\, 
         \$v6280%next\, \$v6280%now\, \$17969%next\, \$17969%now\, 
         \$16404%next\, \$16404%now\, \$17809%next\, \$17809%now\, 
         \$v7134%next\, \$v7134%now\, \$v7276%next\, \$v7276%now\, 
         \$12803_loop666_result%next\, \$12803_loop666_result%now\, 
         \$17970%next\, \$17970%now\, \$v6820%next\, \$v6820%now\, 
         \$17808%next\, \$17808%now\, \$13150%next\, \$13150%now\, 
         \$v6457%next\, \$v6457%now\, \$17499%next\, \$17499%now\, 
         \$12813%next\, \$12813%now\, \$v7282%next\, \$v7282%now\, 
         \$v7012%next\, \$v7012%now\, \$17011%next\, \$17011%now\, 
         \$19265%next\, \$19265%now\, \$v5982%next\, \$v5982%now\, 
         \$v6415%next\, \$v6415%now\, \$v7082%next\, \$v7082%now\, 
         \$v6294%next\, \$v6294%now\, \$13533%next\, \$13533%now\, 
         \$13820%next\, \$13820%now\, \$13812%next\, \$13812%now\, 
         \$17895%next\, \$17895%now\, \$v7111%next\, \$v7111%now\, 
         \$15684_compare6445897_result%next\, 
         \$15684_compare6445897_result%now\, \$12832%next\, \$12832%now\, 
         \$v6358%next\, \$v6358%now\, \$12703%next\, \$12703%now\, 
         \$v6059%next\, \$v6059%now\, \$17166%next\, \$17166%now\, 
         \$v6011%next\, \$v6011%now\, \$v6111%next\, \$v6111%now\, 
         \$12659%next\, \$12659%now\, \$18924%next\, \$18924%now\, 
         \$v6295%next\, \$v6295%now\, \$18190%next\, \$18190%now\, 
         \$v7060%next\, \$v7060%now\, \$v6639%next\, \$v6639%now\, 
         \$v7084%next\, \$v7084%now\, \$v5960%next\, \$v5960%now\, 
         \result6112%next\, \result6112%now\, \$v7032%next\, \$v7032%now\, 
         \$18344%next\, \$18344%now\, \$18992%next\, \$18992%now\, 
         \$13315%next\, \$13315%now\, \$16515%next\, \$16515%now\, 
         \$16156%next\, \$16156%now\, \$17560%next\, \$17560%now\, 
         \$17010%next\, \$17010%now\, \$12846%next\, \$12846%now\, 
         \$12674%next\, \$12674%now\, \$v6315%next\, \$v6315%now\, 
         \$v7031%next\, \$v7031%now\, \$12547%next\, \$12547%now\, 
         \$v7070%next\, \$v7070%now\, \$14471%next\, \$14471%now\, 
         \$18991%next\, \$18991%now\, \$18708%next\, \$18708%now\, 
         \$16508%next\, \$16508%now\, \$v7242%next\, \$v7242%now\, 
         \$v6769%next\, \$v6769%now\, \$v6735%next\, \$v6735%now\, 
         \$19271%next\, \$19271%now\, \$v5983%next\, \$v5983%now\, 
         \$v7033%next\, \$v7033%now\, \$13815%next\, \$13815%now\, 
         \$v5973%next\, \$v5973%now\, \$v6603%next\, \$v6603%now\, 
         \$13018%next\, \$13018%now\, \$v6144%next\, \$v6144%now\, 
         \$v6259%next\, \$v6259%now\, \$13147%next\, \$13147%now\, 
         \$17503%next\, \$17503%now\, \$v6781%next\, \$v6781%now\, 
         \$v6054%next\, \$v6054%now\, \$13232%next\, \$13232%now\, 
         \$v7113%next\, \$v7113%now\, \$v7233%next\, \$v7233%now\, 
         \$17786%next\, \$17786%now\, \$18040%next\, \$18040%now\, 
         \$v6704%next\, \$v6704%now\, \$17544%next\, \$17544%now\, 
         \$v7114%next\, \$v7114%now\, \$v6159%next\, \$v6159%now\, 
         \$13229%next\, \$13229%now\, \$v6332%next\, \$v6332%now\, 
         \$v6968%next\, \$v6968%now\, \$v7041%next\, \$v7041%now\, 
         \$19002%next\, \$19002%now\, \$v7191%next\, \$v7191%now\, 
         \$16534%next\, \$16534%now\, \$13390%next\, \$13390%now\, 
         \$19261%next\, \$19261%now\, \$v7103%next\, \$v7103%now\, 
         \$18047%next\, \$18047%now\, \rdy6148%next\, \rdy6148%now\, 
         \$v7072%next\, \$v7072%now\, \$v6187%next\, \$v6187%now\, 
         \$12708%next\, \$12708%now\, \$13239%next\, \$13239%now\, 
         \$v6476%next\, \$v6476%now\, \$v6002%next\, \$v6002%now\, 
         \$17894%next\, \$17894%now\, \$v6322%next\, \$v6322%now\, 
         \$v7419%next\, \$v7419%now\, \$v6814%next\, \$v6814%now\, 
         \$v6156%next\, \$v6156%now\, \$v7254%next\, \$v7254%now\, 
         \$13528%next\, \$13528%now\, \$18640%next\, \$18640%now\, 
         \$12933%next\, \$12933%now\, \$v6140%next\, \$v6140%now\, 
         \$13963%next\, \$13963%now\, \$18638%next\, \$18638%now\, 
         \$17748%next\, \$17748%now\, \$v6045%next\, \$v6045%now\, 
         \$17310%next\, \$17310%now\, \$v7120%next\, \$v7120%now\, 
         \$v6787%next\, \$v6787%now\, \$17966%next\, \$17966%now\, 
         \$v7096%next\, \$v7096%now\, \$19264%next\, \$19264%now\, 
         \$13311%next\, \$13311%now\, \$12744%next\, \$12744%now\, 
         \$16133%next\, \$16133%now\, \$16232%next\, \$16232%now\, 
         \$18351%next\, \$18351%now\, \$18262%next\, \$18262%now\, 
         \$v6527%next\, \$v6527%now\, \$16568_b%next\, \$16568_b%now\, 
         \$16840_b%next\, \$16840_b%now\, \$14552%next\, \$14552%now\, 
         \$13313%next\, \$13313%now\, \$v6905%next\, \$v6905%now\, 
         \$v6098%next\, \$v6098%now\, \$13023%next\, \$13023%now\, 
         \$v6511%next\, \$v6511%now\, \$v7182%next\, \$v7182%now\, 
         \$12842%next\, \$12842%now\, \$13536%next\, \$13536%now\, 
         \$18049%next\, \$18049%now\, \$v7176%next\, \$v7176%now\, 
         \$16194%next\, \$16194%now\, \$12719%next\, \$12719%now\, 
         \$17758%next\, \$17758%now\, \$17973%next\, \$17973%now\, 
         \$13939%next\, \$13939%now\, \$v7104%next\, \$v7104%now\, 
         \$17747%next\, \$17747%now\, \$12520_loop666_result%next\, 
         \$12520_loop666_result%now\, \$v6796%next\, \$v6796%now\, 
         \$12811%next\, \$12811%now\, \$v6536%next\, \$v6536%now\, 
         \$16510_forever6705925_arg%next\, \$16510_forever6705925_arg%now\, 
         \$16473%next\, \$16473%now\, \$18281%next\, \$18281%now\, 
         \$v7126%next\, \$v7126%now\, \$18735%next\, \$18735%now\, 
         \$v6253%next\, \$v6253%now\, \$v7061%next\, \$v7061%now\, 
         \$17482%next\, \$17482%now\, \$13535%next\, \$13535%now\, 
         \$19143%next\, \$19143%now\, \$v7102%next\, \$v7102%now\, 
         \$18122%next\, \$18122%now\, \$v6705%next\, \$v6705%now\, 
         \$16457%next\, \$16457%now\, \$13538%next\, \$13538%now\, 
         \$v7457%next\, \$v7457%now\, \$18922%next\, \$18922%now\, 
         \$v6759%next\, \$v6759%now\, \$17598%next\, \$17598%now\, 
         \$17972%next\, \$17972%now\, \$18842%next\, \$18842%now\, 
         \$18740%next\, \$18740%now\, \$17677%next\, \$17677%now\, 
         \$13021%next\, \$13021%now\, \$12713%next\, \$12713%now\, 
         \$v6531%next\, \$v6531%now\, \$14069%next\, \$14069%now\, 
         \$17388%next\, \$17388%now\, \$v5867%next\, \$v5867%now\, 
         \$v7051%next\, \$v7051%now\, \$13624%next\, \$13624%now\, 
         \$v7267%next\, \$v7267%now\, \$v6650%next\, \$v6650%now\, 
         \$14148%next\, \$14148%now\, \$17675%next\, \$17675%now\, 
         \$v7112%next\, \$v7112%now\, \$13383%next\, \$13383%now\, 
         \$v6433%next\, \$v6433%now\, \$v7095%next\, \$v7095%now\, 
         \$17320%next\, \$17320%now\, \$v7014%next\, \$v7014%now\, 
         \$14051%next\, \$14051%now\, \$13464%next\, \$13464%now\, 
         \$13236%next\, \$13236%now\, \$17395%next\, \$17395%now\, 
         \$v7296%next\, \$v7296%now\, \$v6784%next\, \$v6784%now\, 
         \$18674%next\, \$18674%now\, \$19136%next\, \$19136%now\, 
         \$v6436%next\, \$v6436%now\, \$13814%next\, \$13814%now\, 
         \$v5947%next\, \$v5947%now\, \$13539%next\, \$13539%now\, 
         \$12743%next\, \$12743%now\, \$v6133%next\, \$v6133%now\, 
         \$v5972%next\, \$v5972%now\, \$18046%next\, \$18046%now\, 
         \$17504%next\, \$17504%now\, \$18993%next\, \$18993%now\, 
         \$v6353%next\, \$v6353%now\, \$v6263%next\, \$v6263%now\, 
         \$v7115%next\, \$v7115%now\, \$18676%next\, \$18676%now\, 
         \$v5876%next\, \$v5876%now\, \$18844%next\, \$18844%now\, 
         \$v7194%next\, \$v7194%now\, \$v7289%next\, \$v7289%now\, 
         \$v7397%next\, \$v7397%now\, \$v6394%next\, \$v6394%now\, 
         \$13695%next\, \$13695%now\, \$17497%next\, \$17497%now\, 
         \$19242%next\, \$19242%now\, \$12814%next\, \$12814%now\, 
         \$17814%next\, \$17814%now\, \$v6409%next\, \$v6409%now\, 
         \$13227%next\, \$13227%now\, \$17673%next\, \$17673%now\, 
         \$16300%next\, \$16300%now\, \$v6752%next\, \$v6752%now\, 
         \$18196%next\, \$18196%now\, \$17347%next\, \$17347%now\, 
         \$19260%next\, \$19260%now\, \$v6335%next\, \$v6335%now\, 
         \$16811_compare6445898_result%next\, 
         \$16811_compare6445898_result%now\, \$14024%next\, \$14024%now\, 
         \$v6666%next\, \$v6666%now\, \$15679_res%next\, \$15679_res%now\, 
         \$v6956%next\, \$v6956%now\, \$v7083%next\, \$v7083%now\, 
         \$13691%next\, \$13691%now\, \$18921%next\, \$18921%now\, 
         \$18326%next\, \$18326%now\, \$v6606%next\, \$v6606%now\, 
         \$14033%next\, \$14033%now\, \$v6219%next\, \$v6219%now\, 
         \$18051%next\, \$18051%now\, \$12889%next\, \$12889%now\, 
         \$v6859%next\, \$v6859%now\, \$12847%next\, \$12847%now\, 
         \$v7101%next\, \$v7101%now\, \$17008%next\, \$17008%now\, 
         \$17595%next\, \$17595%now\, \$18918%next\, \$18918%now\, 
         \$18737%next\, \$18737%now\, \$12760%next\, \$12760%now\, 
         \$v6072%next\, \$v6072%now\, \$18119%next\, \$18119%now\, 
         \$v7197%next\, \$v7197%now\, \$17314%next\, \$17314%now\, 
         \$v6247%next\, \$v6247%now\, \$17759%next\, \$17759%now\, 
         \$16288%next\, \$16288%now\, \$13117%next\, \$13117%now\, 
         \$12696%next\, \$12696%now\, \$12705%next\, \$12705%now\, 
         \$17572%next\, \$17572%now\, \$14281%next\, \$14281%now\, 
         \$v6844%next\, \$v6844%now\, \$v7213%next\, \$v7213%now\, 
         \$12709%next\, \$12709%now\, \$17967%next\, \$17967%now\, 
         \$13626%next\, \$13626%now\, \$16403%next\, \$16403%now\, 
         \$15618%next\, \$15618%now\, \$v7273%next\, \$v7273%now\, 
         \$v7116%next\, \$v7116%now\, \$16507%next\, \$16507%now\, 
         \$v6917%next\, \$v6917%now\, \$15619%next\, \$15619%now\, 
         \$18191%next\, \$18191%now\, \$v6493%next\, \$v6493%now\, 
         \$13529%next\, \$13529%now\, \$v6243%next\, \$v6243%now\, 
         \$17532%next\, \$17532%now\, \$v7046%next\, \$v7046%now\, 
         \$v7449%next\, \$v7449%now\, \$18564%next\, \$18564%now\, 
         \$v7010%next\, \$v7010%now\, \$15860%next\, \$15860%now\, 
         \$13766%next\, \$13766%now\, \$18639%next\, \$18639%now\, 
         \$v5998%next\, \$v5998%now\, \$17968%next\, \$17968%now\, 
         \$v5967%next\, \$v5967%now\, \$15787_res%next\, \$15787_res%now\, 
         \$19214%next\, \$19214%now\, \$18673%next\, \$18673%now\, 
         \$17458_loop666_result%next\, \$17458_loop666_result%now\, 
         \$v7427%next\, \$v7427%now\, \$13688%next\, \$13688%now\, 
         \$12706%next\, \$12706%now\, \$17032%next\, \$17032%now\, 
         \$v6256%next\, \$v6256%now\, \$v6588%next\, \$v6588%now\, 
         \$12934%next\, \$12934%now\, \$v6236%next\, \$v6236%now\, 
         \$v6550%next\, \$v6550%now\, \$v6325%next\, \$v6325%now\, 
         \$v6714%next\, \$v6714%now\, \$13092%next\, \$13092%now\, 
         \$v5948%next\, \$v5948%now\, \$17393%next\, \$17393%now\, 
         \$v6283%next\, \$v6283%now\, \$13158%next\, \$13158%now\, 
         \$18998%next\, \$18998%now\, \$15715_res%next\, \$15715_res%now\, 
         \$v6889%next\, \$v6889%now\, \$v6180%next\, \$v6180%now\, 
         \$v7021%next\, \$v7021%now\, \$v5964%next\, \$v5964%now\, 
         \$v6190%next\, \$v6190%now\, \$17594%next\, \$17594%now\, 
         \$12720%next\, \$12720%now\, \$18044%next\, \$18044%now\, 
         \$v7350%next\, \$v7350%now\, \$18994%next\, \$18994%now\, 
         \$v6152%next\, \$v6152%now\, \$v6643%next\, \$v6643%now\, 
         \$v7260%next\, \$v7260%now\, \$19266%next\, \$19266%now\, 
         \$17048_w16565937_result%next\, \$17048_w16565937_result%now\, 
         \$v6379%next\, \$v6379%now\, \$v7056%next\, \$v7056%now\, 
         \$v6829%next\, \$v6829%now\, \$v7011%next\, \$v7011%now\, 
         \$v6880%next\, \$v6880%now\, \$v6938%next\, \$v6938%now\, 
         \rdy6504%next\, \rdy6504%now\, \$14273%next\, \$14273%now\, 
         \$12829%next\, \$12829%now\, \$13309%next\, \$13309%now\, 
         \$v6684%next\, \$v6684%now\, \$v6352%next\, \$v6352%now\, 
         \$v6031%next\, \$v6031%now\, \$v6075%next\, \$v6075%now\, 
         \$18913%next\, \$18913%now\, \$12710%next\, \$12710%now\, 
         \$v6176%next\, \$v6176%now\, \$v7093%next\, \$v7093%now\, 
         \$18668%next\, \$18668%now\, \$17592%next\, \$17592%now\, 
         \$13385%next\, \$13385%now\, \$18048%next\, \$18048%now\, 
         \$17883%next\, \$17883%now\, \$v7229%next\, \$v7229%now\, 
         \$v7459%next\, \$v7459%now\, \$18572%next\, \$18572%now\, 
         \$19268%next\, \$19268%now\, \$v7156%next\, \$v7156%now\, 
         \$v6899%next\, \$v6899%now\, \$16336%next\, \$16336%now\, 
         \$17173%next\, \$17173%now\, \$v7387%next\, \$v7387%now\, 
         \$v6223%next\, \$v6223%now\, \$v6790%next\, \$v6790%now\, 
         \$v6137%next\, \$v6137%now\, \$18660%next\, \$18660%now\, 
         \$18669%next\, \$18669%now\, \$v6521%next\, \$v6521%now\, 
         \$13818%next\, \$13818%now\, \$15613%next\, \$15613%now\, 
         \$13019%next\, \$13019%now\, \$17164%next\, \$17164%now\, 
         \$13149%next\, \$13149%now\, \$12830%next\, \$12830%now\, 
         \$v6623%next\, \$v6623%now\, \$16440%next\, \$16440%now\, 
         \$18478%next\, \$18478%now\, \$v6616%next\, \$v6616%now\, 
         \$19267%next\, \$19267%now\, \$v6354%next\, \$v6354%now\, 
         \$v7445%next\, \$v7445%now\, \$v6442%next\, \$v6442%now\, 
         \$17243%next\, \$17243%now\, \$v6155%next\, \$v6155%now\, 
         \$v6908%next\, \$v6908%now\, \$12717%next\, \$12717%now\, 
         \$v7167%next\, \$v7167%now\, \$17804%next\, \$17804%now\, 
         \$16626%next\, \$16626%now\, \$18476%next\, \$18476%now\, 
         \$v6902%next\, \$v6902%now\, \$15909%next\, \$15909%now\, 
         \$18470%next\, \$18470%now\, \$v6184%next\, \$v6184%now\, 
         \$v6547%next\, \$v6547%now\, \$18041%next\, \$18041%now\, 
         \$12942%next\, \$12942%now\, \$17502%next\, \$17502%now\, 
         \$v6036%next\, \$v6036%now\, \$v6660%next\, \$v6660%now\, 
         \$17066%next\, \$17066%now\, \$18732%next\, \$18732%now\, 
         \$v6535%next\, \$v6535%now\, \$v6553%next\, \$v6553%now\, 
         \$v6109%next\, \$v6109%now\, \$v6093%next\, \$v6093%now\, 
         \$12688%next\, \$12688%now\, \$16509%next\, \$16509%now\, 
         \$18738%next\, \$18738%now\, \$13316%next\, \$13316%now\, 
         \$18841%next\, \$18841%now\, \$v6766%next\, \$v6766%now\, 
         \$v7393%next\, \$v7393%now\, \$v5872%next\, \$v5872%now\, 
         \$v7081%next\, \$v7081%now\, \$v7020%next\, \$v7020%now\, 
         \$18546%next\, \$18546%now\, \$v6965%next\, \$v6965%now\, 
         \$v6319%next\, \$v6319%now\, \$v7044%next\, \$v7044%now\, 
         \$v6328%next\, \$v6328%now\, \$14008%next\, \$14008%now\, 
         \$18845%next\, \$18845%now\, \$v7375%next\, \$v7375%now\, 
         \$v6742%next\, \$v6742%now\, \$v7378%next\, \$v7378%now\, 
         \$13463%next\, \$13463%now\, \$v7426%next\, \$v7426%now\, 
         \$v6743%next\, \$v6743%now\, \$v6562%next\, \$v6562%now\, 
         \$v7188%next\, \$v7188%now\, \$v6692%next\, \$v6692%now\, 
         \$v6646%next\, \$v6646%now\, \$v7332%next\, \$v7332%now\, 
         \$v6758%next\, \$v6758%now\, \$18473%next\, \$18473%now\, 
         \$v6171%next\, \$v6171%now\, \$v6373%next\, \$v6373%now\, 
         \$v5995%next\, \$v5995%now\, \$15910%next\, \$15910%now\, 
         \$v6835%next\, \$v6835%now\, \$17513_forever6705889_arg%next\, 
         \$17513_forever6705889_arg%now\, \$v7100%next\, \$v7100%now\, 
         \$v6862%next\, \$v6862%now\, \$13540%next\, \$13540%now\, 
         \$18118%next\, \$18118%now\, \$v7110%next\, \$v7110%now\, 
         \$12704%next\, \$12704%now\, \$17671%next\, \$17671%now\, 
         \$v6585%next\, \$v6585%now\, \$v6543%next\, \$v6543%now\, 
         \$17892%next\, \$17892%now\, \$18184%next\, \$18184%now\, 
         \$18730%next\, \$18730%now\, \$v6765%next\, \$v6765%now\, 
         \$v6832%next\, \$v6832%now\, \$v7365%next\, \$v7365%now\, 
         \$13384%next\, \$13384%now\, \$v5986%next\, \$v5986%now\, 
         \$16321%next\, \$16321%now\, \$v6989%next\, \$v6989%now\, 
         \$v6920%next\, \$v6920%now\, \$17964%next\, \$17964%now\, 
         \rdy6469%next\, \rdy6469%now\, \$18189%next\, \$18189%now\, 
         \$15447_forever6705911_arg%next\, \$15447_forever6705911_arg%now\, 
         \$v6717%next\, \$v6717%now\, \$13234%next\, \$13234%now\, 
         \$v6042%next\, \$v6042%now\, \$v6654%next\, \$v6654%now\, 
         \$12701%next\, \$12701%now\, \$12694%next\, \$12694%now\, 
         \$19118%next\, \$19118%now\, \$17561%next\, \$17561%now\, 
         \$v6096%next\, \$v6096%now\, \$v6069%next\, \$v6069%now\, 
         \$13101%next\, \$13101%now\, \$18348%next\, \$18348%now\, 
         \$16317%next\, \$16317%now\, \$v7245%next\, \$v7245%now\, 
         \$18843%next\, \$18843%now\, \$13700%next\, \$13700%now\, 
         \$12938%next\, \$12938%now\, \$18806%next\, \$18806%now\, 
         \$v7135%next\, \$v7135%now\, \$16382%next\, \$16382%now\, 
         \$12903%next\, \$12903%now\, \$v6287%next\, \$v6287%now\, 
         \$13317%next\, \$13317%now\, \$18657%next\, \$18657%now\, 
         \$v7433%next\, \$v7433%now\, \$13940%next\, \$13940%now\, 
         \$13510%next\, \$13510%now\, \$v6421%next\, \$v6421%now\, 
         \$17805%next\, \$17805%now\, \$17500%next\, \$17500%now\, 
         \$v6424%next\, \$v6424%now\, \$12735%next\, \$12735%now\, 
         \$v6403%next\, \$v6403%now\, \$13822%next\, \$13822%now\, 
         \$v7203%next\, \$v7203%now\, \$v6097%next\, \$v6097%now\, 
         \$13100%next\, \$13100%now\, \$v6463%next\, \$v6463%now\, 
         \$17815%next\, \$17815%now\, \$14296%next\, \$14296%now\, 
         \$v7092%next\, \$v7092%now\, \$v6799%next\, \$v6799%now\, 
         \$v6080%next\, \$v6080%now\, \$v6563%next\, \$v6563%now\, 
         \$v6062%next\, \$v6062%now\, \$v6817%next\, \$v6817%now\, 
         \$13817%next\, \$13817%now\, \$v6670%next\, \$v6670%now\, 
         \$12886%next\, \$12886%now\, \$v7364%next\, \$v7364%now\, 
         \$v6232%next\, \$v6232%now\, \$13148%next\, \$13148%now\, 
         \$18280%next\, \$18280%now\, \$v6546%next\, \$v6546%now\, 
         \$v7206%next\, \$v7206%now\, \$v5999%next\, \$v5999%now\, 
         \$v6971%next\, \$v6971%now\, \$14311%next\, \$14311%now\, 
         \$17889%next\, \$17889%now\, \$v6207%next\, \$v6207%now\, 
         \$v6911%next\, \$v6911%now\, \$v6066%next\, \$v6066%now\, 
         \$14381%next\, \$14381%now\, \$18043%next\, \$18043%now\, 
         \$v6179%next\, \$v6179%now\, \$v6110%next\, \$v6110%now\, 
         \$18995%next\, \$18995%now\, \$13689%next\, \$13689%now\, 
         \$v6121%next\, \$v6121%now\, \$v6579%next\, \$v6579%now\, 
         \$17466%next\, \$17466%now\, \$v6003%next\, \$v6003%now\, 
         \$v6898%next\, \$v6898%now\, \$16986_compare6445898_result%next\, 
         \$16986_compare6445898_result%now\, \$17593%next\, \$17593%now\, 
         \$v6515%next\, \$v6515%now\, \$v6992%next\, \$v6992%now\, 
         \$v6624%next\, \$v6624%now\, \$18571%next\, \$18571%now\, 
         \$v7210%next\, \$v7210%now\, \$17812%next\, \$17812%now\, 
         \$18193%next\, \$18193%now\, \$18194%next\, \$18194%now\, 
         \$13129%next\, \$13129%now\, \$14135%next\, \$14135%now\, 
         \$12716%next\, \$12716%now\, \$17785%next\, \$17785%now\, 
         \$v6998%next\, \$v6998%now\, \$18187%next\, \$18187%now\, 
         \$17775%next\, \$17775%now\, \$v6724%next\, \$v6724%now\, 
         \$12736%next\, \$12736%now\, \$v7232%next\, \$v7232%now\, 
         \$12660%next\, \$12660%now\, \$12936%next\, \$12936%now\, 
         \$15828_compare6445897_result%next\, 
         \$15828_compare6445897_result%now\, \$17890%next\, \$17890%now\, 
         \$18475%next\, \$18475%now\, \$12913%next\, \$12913%now\, 
         \$v6388%next\, \$v6388%now\, \$v6400%next\, \$v6400%now\, 
         \$v7091%next\, \$v7091%now\, \$v7015%next\, \$v7015%now\, 
         \$16231%next\, \$16231%now\, \$17774%next\, \$17774%now\, 
         \$v6089%next\, \$v6089%now\, \$12695%next\, \$12695%now\, 
         \$v7054%next\, \$v7054%now\, \$18356%next\, \$18356%now\, 
         \$v7328%next\, \$v7328%now\, \$13694%next\, \$13694%now\, 
         \$17254%next\, \$17254%now\, \$19070%next\, \$19070%now\, 
         \$v6286%next\, \$v6286%now\, \$13238%next\, \$13238%now\, 
         \$v6847%next\, \$v6847%now\, \$19262%next\, \$19262%now\, 
         \$12914%next\, \$12914%now\, \$13794%next\, \$13794%now\, 
         \$17783%next\, \$17783%now\, \$12941%next\, \$12941%now\, 
         \$v6048%next\, \$v6048%now\, \$18679_forever6705881_arg%next\, 
         \$18679_forever6705881_arg%now\, \$17495%next\, \$17495%now\, 
         \$17590%next\, \$17590%now\, \$13387%next\, \$13387%now\, 
         \$13393%next\, \$13393%now\, \$17348%next\, \$17348%now\, 
         \$18677%next\, \$18677%now\, \$13389%next\, \$13389%now\, 
         \$14254%next\, \$14254%now\, \$18185%next\, \$18185%now\, 
         \$18472%next\, \$18472%now\, \$v6012%next\, \$v6012%now\, 
         \$v6162%next\, \$v6162%now\, \$v7458%next\, \$v7458%now\, 
         \$17455_loop666_result%next\, \$17455_loop666_result%now\, 
         \$v6595%next\, \$v6595%now\, \$v6947%next\, \$v6947%now\, 
         \$v6314%next\, \$v6314%now\, \$v5992%next\, \$v5992%now\, 
         \$v6183%next\, \$v6183%now\, \$18711%next\, \$18711%now\, 
         \$v5878%next\, \$v5878%now\, \$v7076%next\, \$v7076%now\, 
         \$15792_compare6445897_result%next\, 
         \$15792_compare6445897_result%now\, \$13312%next\, \$13312%now\, 
         \$12702%next\, \$12702%now\, \$v6364%next\, \$v6364%now\, 
         \$v6678%next\, \$v6678%now\, \$v6738%next\, \$v6738%now\, 
         \$v7030%next\, \$v7030%now\, \$18104%next\, \$18104%now\, 
         \$v6165%next\, \$v6165%now\, \$16767%next\, \$16767%now\, 
         \$16292%next\, \$16292%now\, \$v6751%next\, \$v6751%now\, 
         \$17463%next\, \$17463%now\, \$v7322%next\, \$v7322%now\, 
         \$13466%next\, \$13466%now\, \$v6853%next\, \$v6853%now\, 
         \$12904%next\, \$12904%now\, \$12734%next\, \$12734%now\, 
         \$v6229%next\, \$v6229%now\, \$13693%next\, \$13693%now\, 
         \$v7185%next\, \$v7185%now\, \$v5874%next\, \$v5874%now\, 
         \$v6301%next\, \$v6301%now\, \$18637%next\, \$18637%now\, 
         \$18999%next\, \$18999%now\, \$v7086%next\, \$v7086%now\, 
         \$v6773%next\, \$v6773%now\, \$v7219%next\, \$v7219%now\, 
         \$12857_forever6705883_arg%next\, \$12857_forever6705883_arg%now\, 
         \$18836%next\, \$18836%now\, \$16031%next\, \$16031%now\, 
         \$12878%next\, \$12878%now\, \$v7133%next\, \$v7133%now\, 
         \$16126%next\, \$16126%now\, \$17377%next\, \$17377%now\, 
         \$13928_w652_result%next\, \$13928_w652_result%now\, \$16035%next\, 
         \$16035%now\, \$18166%next\, \$18166%now\, \$v7416%next\, 
         \$v7416%now\, \$12939%next\, \$12939%now\, \$14042%next\, 
         \$14042%now\, \$13307%next\, \$13307%now\, \$17315%next\, 
         \$17315%now\, \$13946%next\, \$13946%now\, \$18818%next\, 
         \$18818%now\, \$v6175%next\, \$v6175%now\, \$v7121%next\, 
         \$v7121%now\, \$v6865%next\, \$v6865%now\, \$v6102%next\, 
         \$v6102%now\, \$v6609%next\, \$v6609%now\, \$14558%next\, 
         \$14558%now\, \$v7335%next\, \$v7335%now\, \$v6950%next\, 
         \$v6950%now\, \$v7453%next\, \$v7453%now\, \$v6701%next\, 
         \$v6701%now\, \$13153%next\, \$13153%now\, \$v6055%next\, 
         \$v6055%now\, \$18734%next\, \$18734%now\, 
         \$12806_loop666_result%next\, \$12806_loop666_result%now\, 
         \$v6681%next\, \$v6681%now\, \$v6271%next\, \$v6271%now\, 
         \$v7358%next\, \$v7358%now\, \$18479%next\, \$18479%now\, 
         \$13692%next\, \$13692%now\, \$v7023%next\, \$v7023%now\, 
         \$13103%next\, \$13103%now\, \$v6268%next\, \$v6268%now\, 
         \$v6307%next\, \$v6307%now\, \$v7016%next\, \$v7016%now\, 
         \$13957%next\, \$13957%now\, \$v6214%next\, \$v6214%now\, 
         \$17600%next\, \$17600%now\, \$v6657%next\, \$v6657%now\, 
         \$v6995%next\, \$v6995%now\, \$12943%next\, \$12943%now\, 
         \$v6117%next\, \$v6117%now\, \$v7368%next\, \$v7368%now\, 
         \$v7064%next\, \$v7064%now\, \$12843%next\, \$12843%now\, 
         \$14161%next\, \$14161%now\, \$13962%next\, \$13962%now\, 
         \$v7441%next\, \$v7441%now\, \$v6962%next\, \$v6962%now\, 
         \$v6277%next\, \$v6277%now\, \$v7455%next\, \$v7455%now\, 
         \$12741%next\, \$12741%now\, \$v6445%next\, \$v6445%now\, 
         \$17681%next\, \$17681%now\, \$17961%next\, \$17961%now\, 
         \$16805_b%next\, \$16805_b%now\, \$v6986%next\, \$v6986%now\, 
         \$v6935%next\, \$v6935%now\, \$v6750%next\, \$v6750%now\, 
         \$v7066%next\, \$v7066%now\, \$v6007%next\, \$v6007%now\, 
         \$v7140%next\, \$v7140%now\, \$16234%next\, \$16234%now\, 
         \$12679_loop666_result%next\, \$12679_loop666_result%now\, 
         \$17167%next\, \$17167%now\, \$12834%next\, \$12834%now\, 
         \$16192%next\, \$16192%now\, \$17349%next\, \$17349%now\, 
         \$13013%next\, \$13013%now\, \$18450%next\, \$18450%now\, 
         \$v5951%next\, \$v5951%now\, \$v5866%next\, \$v5866%now\, 
         \$v6203%next\, \$v6203%now\, \$v6868%next\, \$v6868%now\, 
         \$14222%next\, \$14222%now\, \$13530%next\, \$13530%now\, 
         \$v6709%next\, \$v6709%now\, \$v7090%next\, \$v7090%now\, 
         \$v7004%next\, \$v7004%now\, \$13127%next\, \$13127%now\, 
         \$v7179%next\, \$v7179%now\, \$15847%next\, \$15847%now\, 
         \$16606_b%next\, \$16606_b%now\, \$v5954%next\, \$v5954%now\, 
         \$v6342%next\, \$v6342%now\, \$v7299%next\, \$v7299%now\, 
         \$16165%next\, \$16165%now\, \$16078%next\, \$16078%now\, 
         \$13941%next\, \$13941%now\, \$17319%next\, \$17319%now\, 
         \$v7361%next\, \$v7361%now\, \$v6688%next\, \$v6688%now\, 
         \$16612_compare6445898_result%next\, 
         \$16612_compare6445898_result%now\, \$v6200%next\, \$v6200%now\, 
         \$v6367%next\, \$v6367%now\, \$17962%next\, \$17962%now\, 
         \$12691%next\, \$12691%now\, \$v7013%next\, \$v7013%now\, 
         \$v6651%next\, \$v6651%now\, \$v7372%next\, \$v7372%now\, 
         \$v6574%next\, \$v6574%now\, \$v6874%next\, \$v6874%now\, 
         \$16158_forever6705923_arg%next\, \$16158_forever6705923_arg%now\, 
         \$v6695%next\, \$v6695%now\, \$17394%next\, \$17394%now\, 
         \$v6826%next\, \$v6826%now\, \$12887%next\, \$12887%now\, 
         \$v7042%next\, \$v7042%now\, \$v7164%next\, \$v7164%now\, 
         \$17885%next\, \$17885%now\, \$18816%next\, \$18816%now\, 
         \$v7045%next\, \$v7045%now\, \$19263%next\, \$19263%now\, 
         \$16399%next\, \$16399%now\, \$v7248%next\, \$v7248%now\, 
         \$13623%next\, \$13623%now\, \$18570%next\, \$18570%now\, 
         \$v6856%next\, \$v6856%now\, \$v6710%next\, \$v6710%now\, 
         \$12848%next\, \$12848%now\, \$19071%next\, \$19071%now\, 
         \$19140%next\, \$19140%now\, \$15612%next\, \$15612%now\, 
         \$v6883%next\, \$v6883%now\, \$16875_b%next\, \$16875_b%now\, 
         \$17678%next\, \$17678%now\, \$v7034%next\, \$v7034%now\, 
         \$16677%next\, \$16677%now\, \$19144%next\, \$19144%now\, 
         \$13890%next\, \$13890%now\, \$18915%next\, \$18915%now\, 
         \$v6914%next\, \$v6914%now\, \$v6729%next\, \$v6729%now\, 
         \$17387%next\, \$17387%now\, \$v6892%next\, \$v6892%now\, 
         \$v6492%next\, \$v6492%now\, \$18045%next\, \$18045%now\, 
         \$v6136%next\, \$v6136%now\, \$12915%next\, \$12915%now\, 
         \$v6627%next\, \$v6627%now\, \$17591%next\, \$17591%now\, 
         \$18699%next\, \$18699%now\, \$12715%next\, \$12715%now\, 
         \$16365%next\, \$16365%now\, \$16574_compare6445898_result%next\, 
         \$16574_compare6445898_result%now\, \$17354%next\, \$17354%now\, 
         \$12945%next\, \$12945%now\, \$12712%next\, \$12712%now\, 
         \$17674%next\, \$17674%now\, \$13157%next\, \$13157%now\, 
         \$v6708%next\, \$v6708%now\, \$18346%next\, \$18346%now\, 
         \$16945_b%next\, \$16945_b%now\, \$17498%next\, \$17498%now\, 
         \$19001%next\, \$19001%now\, \$v6274%next\, \$v6274%now\, 
         \$17509_forever6705890_arg%next\, \$17509_forever6705890_arg%now\, 
         \$v6739%next\, \$v6739%now\, \$v7434%next\, \$v7434%now\, 
         \$13625%next\, \$13625%now\, \$12935%next\, \$12935%now\, 
         \$12692%next\, \$12692%now\, \$v6304%next\, \$v6304%now\, 
         \$13016%next\, \$13016%now\, \$18120%next\, \$18120%now\, 
         \$v7025%next\, \$v7025%now\, \$18279%next\, \$18279%now\, 
         \$v6953%next\, \$v6953%now\, \$v5957%next\, \$v5957%now\, 
         \$18733%next\, \$18733%now\, \$v6838%next\, \$v6838%now\, 
         \$18925%next\, \$18925%now\, \$v6746%next\, \$v6746%now\, 
         \$v6941%next\, \$v6941%now\, \$v7007%next\, \$v7007%now\, 
         \$17412%next\, \$17412%now\, \$19269%next\, \$19269%now\, 
         \$17559%next\, \$17559%now\, \$v6239%next\, \$v6239%now\, 
         \$16353%next\, \$16353%now\, \$13395%next\, \$13395%now\, 
         \$13823%next\, \$13823%now\, \$18709%next\, \$18709%now\, 
         \$v6397%next\, \$v6397%now\, \$v7035%next\, \$v7035%now\, 
         \$v7216%next\, \$v7216%now\, \$v6172%next\, \$v6172%now\, 
         \$18188%next\, \$18188%now\, \$12851%next\, \$12851%now\, 
         \$14431%next\, \$14431%now\, \$v6460%next\, \$v6460%now\, 
         \$v7279%next\, \$v7279%now\, \$18186%next\, \$18186%now\, 
         \$v6501%next\, \$v6501%now\, \$12685%next\, \$12685%now\, 
         \$18919%next\, \$18919%now\, \$v7293%next\, \$v7293%now\, 
         \$v6532%next\, \$v6532%now\, \$v6291%next\, \$v6291%now\, 
         \$19142%next\, \$19142%now\, \$17803%next\, \$17803%now\, 
         \$17963%next\, \$17963%now\, \$v6480%next\, \$v6480%now\, 
         \$13388%next\, \$13388%now\, \$17505_forever6705894_arg%next\, 
         \$17505_forever6705894_arg%now\, \$v6235%next\, \$v6235%now\, 
         \$14012%next\, \$14012%now\, \$13310%next\, \$13310%now\, 
         \$18563%next\, \$18563%now\, \$14122%next\, \$14122%now\, 
         \$v6058%next\, \$v6058%now\, \$v6633%next\, \$v6633%now\, 
         \$16327%next\, \$16327%now\, \$13606%next\, \$13606%now\, 
         \$18731%next\, \$18731%now\, \$v7085%next\, \$v7085%now\, 
         \$12544%next\, \$12544%now\, \$18278%next\, \$18278%now\, 
         \$v6518%next\, \$v6518%now\, \$v6298%next\, \$v6298%now\, 
         \$v6732%next\, \$v6732%now\, \$16881_compare6445898_result%next\, 
         \$16881_compare6445898_result%now\, \$12707%next\, \$12707%now\, 
         \$v7074%next\, \$v7074%now\, \$v7306%next\, \$v7306%now\, 
         \$17891%next\, \$17891%now\, \$v5944%next\, \$v5944%now\, 
         \$v5963%next\, \$v5963%now\, \$13950%next\, \$13950%now\, 
         \$17746%next\, \$17746%now\, \$v6596%next\, \$v6596%now\, 
         \$15874%next\, \$15874%now\, \$v6211%next\, \$v6211%now\, 
         \$13816%next\, \$13816%now\, \$v6591%next\, \$v6591%now\, 
         \$v6508%next\, \$v6508%now\, \$v7413%next\, \$v7413%now\, 
         \$v6667%next\, \$v6667%now\, \$v6489%next\, \$v6489%now\, 
         \$v6406%next\, \$v6406%now\, \$15893%next\, \$15893%now\, 
         \$19145%next\, \$19145%now\, \$17888%next\, \$17888%now\, 
         \$v7200%next\, \$v7200%now\, \$v7132%next\, \$v7132%now\, 
         \$v7406%next\, \$v7406%now\, \$v6218%next\, \$v6218%now\, 
         \$15823_res%next\, \$15823_res%now\, \$v6780%next\, \$v6780%now\, 
         \$v7144%next\, \$v7144%now\, \$18480%next\, \$18480%now\, 
         \$18698%next\, \$18698%now\, \$12877%next\, \$12877%now\, 
         \$18565%next\, \$18565%now\, \$v6559%next\, \$v6559%now\, 
         \$18815%next\, \$18815%now\, \$v6015%next\, \$v6015%now\, 
         \$13696%next\, \$13696%now\, \$17669%next\, \$17669%now\, 
         \$v6318%next\, \$v6318%now\, \$v6430%next\, \$v6430%now\, 
         \$v6599%next\, \$v6599%now\, \$17464%next\, \$17464%now\, 
         \$v6802%next\, \$v6802%now\, \$14555%next\, \$14555%now\, 
         \$17670%next\, \$17670%now\, \$13233%next\, \$13233%now\, 
         \$v6376%next\, \$v6376%now\, \$13235%next\, \$13235%now\, 
         \$13102%next\, \$13102%now\, \rdy5940%next\, \rdy5940%now\, 
         \$18355%next\, \$18355%now\, \$v6466%next\, \$v6466%now\, 
         \$13697%next\, \$13697%now\, \$v6021%next\, \$v6021%now\, 
         \$16115%next\, \$16115%now\, \$12937%next\, \$12937%now\, 
         \$13155%next\, \$13155%now\, \$12888%next\, \$12888%now\, 
         \$v7344%next\, \$v7344%now\, \$17773%next\, \$17773%now\, 
         \$12697%next\, \$12697%now\, \$v6146%next\, \$v6146%now\, 
         \$13237%next\, \$13237%now\, \$v7454%next\, \$v7454%now\, 
         \$v6496%next\, \$v6496%now\, \$v5869%next\, \$v5869%now\, 
         \$v6500%next\, \$v6500%now\, \$v6728%next\, \$v6728%now\, 
         \$17543%next\, \$17543%now\, \$18805%next\, \$18805%now\, 
         \$18837%next\, \$18837%now\, \$v6027%next\, \$v6027%now\, 
         \$18807%next\, \$18807%now\, \$12689%next\, \$12689%now\, 
         \$v7050%next\, \$v7050%now\, \$v7338%next\, \$v7338%now\, 
         \$v6721%next\, \$v6721%now\, \$v6823%next\, \$v6823%now\, 
         \$13532%next\, \$13532%now\, \$15756_compare6445897_result%next\, 
         \$15756_compare6445897_result%now\, \$17597%next\, \$17597%now\, 
         \$17484%next\, \$17484%now\, \$12714%next\, \$12714%now\, 
         \$18739%next\, \$18739%now\, \$v6370%next\, \$v6370%now\, 
         \$v6502%next\, \$v6502%now\, \$v7420%next\, \$v7420%now\, 
         \$13964%next\, \$13964%now\, \$18352%next\, \$18352%now\, 
         \$v6336%next\, \$v6336%now\, \$13154%next\, \$13154%now\, 
         \$17679%next\, \$17679%now\, \$18916%next\, \$18916%now\, 
         \$v6092%next\, \$v6092%now\, \$18917%next\, \$18917%now\, 
         \$18846%next\, \$18846%now\, \$v7381%next\, \$v7381%now\, 
         \$12944%next\, \$12944%now\, \$v6035%next\, \$v6035%now\, 
         \$12698%next\, \$12698%now\, \$17569%next\, \$17569%now\, 
         \$v6805%next\, \$v6805%now\, \$13151%next\, \$13151%now\, 
         \$17886%next\, \$17886%now\, \$18474%next\, \$18474%now\, 
         \$v6974%next\, \$v6974%now\, \$16748%next\, \$16748%now\, 
         \$v6427%next\, \$v6427%now\, \$v6619%next\, \$v6619%now\, 
         \$v7371%next\, \$v7371%now\, \$18655%next\, \$18655%now\, 
         \$16271%next\, \$16271%now\, \$16233%next\, \$16233%now\, 
         \$18050%next\, \$18050%now\, \$v7353%next\, \$v7353%now\, 
         \$15445%next\, \$15445%now\, \$17386%next\, \$17386%now\, 
         \$v6240%next\, \$v6240%now\, \$14326%next\, \$14326%now\, 
         \$v6385%next\, \$v6385%now\, \$17494%next\, \$17494%now\, 
         \$v7251%next\, \$v7251%now\, \$12853_forever6705887_arg%next\, 
         \$12853_forever6705887_arg%now\, \$v6382%next\, \$v6382%now\, 
         \$17121%next\, \$17121%now\, \$v6348%next\, \$v6348%now\, 
         \$17971%next\, \$17971%now\, \$13531%next\, \$13531%now\, 
         \$v6959%next\, \$v6959%now\, \$13824%next\, \$13824%now\, 
         \$18838%next\, \$18838%now\, \$v6391%next\, \$v6391%now\, 
         \$v7094%next\, \$v7094%now\, \$13945%next\, \$13945%now\, 
         \$19138%next\, \$19138%now\, \$v6575%next\, \$v6575%now\, 
         \$13156%next\, \$13156%now\, \$16141%next\, \$16141%now\, 
         \$v7236%next\, \$v7236%now\, \$15614_forever6705914_arg%next\, 
         \$15614_forever6705914_arg%now\, \$v7170%next\, \$v7170%now\, 
         \$v6206%next\, \$v6206%now\, \$13308%next\, \$13308%now\, 
         \$v6512%next\, \$v6512%now\, \$v7222%next\, \$v7222%now\, 
         \$18121%next\, \$18121%now\, \$17676%next\, \$17676%now\, 
         \$17570%next\, \$17570%now\, \$v7437%next\, \$v7437%now\, 
         \$17893%next\, \$17893%now\, \$19003%next\, \$19003%now\, 
         \$13090%next\, \$13090%now\, \$v7125%next\, \$v7125%now\, 
         \$12699%next\, \$12699%now\, \$v6567%next\, \$v6567%now\, 
         \$18835%next\, \$18835%now\, \$18997%next\, \$18997%now\, 
         \$17887%next\, \$17887%now\, \$v6473%next\, \$v6473%now\, 
         \$12852%next\, \$12852%now\, \$v7062%next\, \$v7062%now\, 
         \$12545_x%next\, \$12545_x%now\, \$v6451%next\, \$v6451%now\, 
         \$18354%next\, \$18354%now\, \$16182%next\, \$16182%now\, 
         \$v6725%next\, \$v6725%now\, \$v6127%next\, \$v6127%now\, 
         \$13670%next\, \$13670%now\, \$18192%next\, \$18192%now\, 
         \$18729%next\, \$18729%now\, \$v6642%next\, \$v6642%now\, 
         \$v7123%next\, \$v7123%now\, \$19272%next\, \$19272%now\, 
         \$v6197%next\, \$v6197%now\, \$v7263%next\, \$v7263%now\, 
         \$v6130%next\, \$v6130%now\, \$12673_rdy%next\, \$12673_rdy%now\, 
         \$18996%next\, \$18996%now\, \$13392%next\, \$13392%now\, 
         \$v7022%next\, \$v7022%now\, \$v6841%next\, \$v6841%now\, 
         \$17813%next\, \$17813%now\, \$v6570%next\, \$v6570%now\, 
         \$v6454%next\, \$v6454%now\, \$14060%next\, \$14060%now\ : value(0 to 0) := (others => '0');
  signal \$13926_make_block_n646_arg%next\, \$13926_make_block_n646_arg%now\ : value(0 to 171) := (others => '0');
  signal \$13924_apply638_arg%next\, \$13924_apply638_arg%now\ : value(0 to 165) := (others => '0');
  signal \$18793_copy_root_in_ram6635879_arg%next\, 
         \$18793_copy_root_in_ram6635879_arg%now\, 
         \$18686_copy_root_in_ram6635880_arg%next\, 
         \$18686_copy_root_in_ram6635880_arg%now\, 
         \$13078_copy_root_in_ram6635885_arg%next\, 
         \$13078_copy_root_in_ram6635885_arg%now\, 
         \$17520_copy_root_in_ram6635893_arg%next\, 
         \$17520_copy_root_in_ram6635893_arg%now\, \$12824%next\, 
         \$12824%now\, \$16662_fill6535928_arg%next\, 
         \$16662_fill6535928_arg%now\, \$12681_wait662_result%next\, 
         \$12681_wait662_result%now\, 
         \$17547_copy_root_in_ram6635891_arg%next\, 
         \$17547_copy_root_in_ram6635891_arg%now\, 
         \$17761_copy_root_in_ram6635891_arg%next\, 
         \$17761_copy_root_in_ram6635891_arg%now\, \$17476%next\, 
         \$17476%now\, \$12737%next\, \$12737%now\, 
         \$13105_copy_root_in_ram6635884_arg%next\, 
         \$13105_copy_root_in_ram6635884_arg%now\, 
         \$12864_copy_root_in_ram6635886_arg%next\, 
         \$12864_copy_root_in_ram6635886_arg%now\, \$17389%next\, 
         \$17389%now\, \$13922_wait662_result%next\, 
         \$13922_wait662_result%now\, \$17048_w16565937_arg%next\, 
         \$17048_w16565937_arg%now\, \$12522_wait662_result%next\, 
         \$12522_wait662_result%now\, 
         \$17734_copy_root_in_ram6635892_arg%next\, 
         \$17734_copy_root_in_ram6635892_arg%now\, 
         \$12891_copy_root_in_ram6635884_arg%next\, 
         \$12891_copy_root_in_ram6635884_arg%now\, \$18566%next\, 
         \$18566%now\, \$18650%next\, \$18650%now\, 
         \$16752_fill6545929_arg%next\, \$16752_fill6545929_arg%now\, 
         \$17018_w36575938_arg%next\, \$17018_w36575938_arg%now\ : value(0 to 79) := (others => '0');
  signal \$17444%next\, \$17444%now\, \$18611%next\, \$18611%now\, 
         \$18621%next\, \$18621%now\, \$17434%next\, \$17434%now\, 
         \$12792%next\, \$12792%now\, \$12782%next\, \$12782%now\ : value(0 to 128) := (others => '0');
  signal \$15625_binop_compare6455916_arg%next\, 
         \$15625_binop_compare6455916_arg%now\, \$16301%next\, \$16301%now\, 
         \$15044_binop_int6435906_arg%next\, 
         \$15044_binop_int6435906_arg%now\, \$16383%next\, \$16383%now\, 
         \$16337%next\, \$16337%now\, \$14724_binop_int6435902_arg%next\, 
         \$14724_binop_int6435902_arg%now\, \$16272%next\, \$16272%now\, 
         \$14964_binop_int6435905_arg%next\, 
         \$14964_binop_int6435905_arg%now\, 
         \$15451_binop_int6435912_arg%next\, 
         \$15451_binop_int6435912_arg%now\, 
         \$14884_binop_int6435904_arg%next\, 
         \$14884_binop_int6435904_arg%now\, 
         \$15364_binop_int6435910_arg%next\, 
         \$15364_binop_int6435910_arg%now\, 
         \$15204_binop_int6435908_arg%next\, 
         \$15204_binop_int6435908_arg%now\, 
         \$15284_binop_int6435909_arg%next\, 
         \$15284_binop_int6435909_arg%now\, 
         \$14644_binop_int6435901_arg%next\, 
         \$14644_binop_int6435901_arg%now\, 
         \$14804_binop_int6435903_arg%next\, 
         \$14804_binop_int6435903_arg%now\, 
         \$15124_binop_int6435907_arg%next\, 
         \$15124_binop_int6435907_arg%now\, 
         \$15733_binop_compare6455919_arg%next\, 
         \$15733_binop_compare6455919_arg%now\, 
         \$15805_binop_compare6455921_arg%next\, 
         \$15805_binop_compare6455921_arg%now\, \$16441%next\, \$16441%now\, 
         \$15697_binop_compare6455918_arg%next\, 
         \$15697_binop_compare6455918_arg%now\, 
         \$15769_binop_compare6455920_arg%next\, 
         \$15769_binop_compare6455920_arg%now\, 
         \$15661_binop_compare6455917_arg%next\, 
         \$15661_binop_compare6455917_arg%now\, 
         \$15531_binop_int6435913_arg%next\, 
         \$15531_binop_int6435913_arg%now\, 
         \$14564_binop_int6435900_arg%next\, 
         \$14564_binop_int6435900_arg%now\ : value(0 to 153) := (others => '0');
  signal \$12654%next\, \$12654%now\, \$13374_w%next\, \$13374_w%now\, 
         \$13628%next\, \$13628%now\, \$13093%next\, \$13093%now\, 
         \$15465_v%next\, \$15465_v%now\, \$13803_w%next\, \$13803_w%now\, 
         \$18340_hd%next\, \$18340_hd%now\, \$16437_v%next\, \$16437_v%now\, 
         \$14025_v%next\, \$14025_v%now\, \$v7087%next\, \$v7087%now\, 
         \$13120%next\, \$13120%now\, \$14493_v%next\, \$14493_v%now\, 
         \$v7141%next\, \$v7141%now\, \$14393_hd%next\, \$14393_hd%now\, 
         \$16041_v%next\, \$16041_v%now\, \$16335_v%next\, \$16335_v%now\, 
         \$14002_v%next\, \$14002_v%now\, \$13889%next\, \$13889%now\, 
         \$18545%next\, \$18545%now\, \$14081%next\, \$14081%now\, 
         \$17660_w%next\, \$17660_w%now\, \$13987_v%next\, \$13987_v%now\, 
         \$16313_v%next\, \$16313_v%now\, \$19132_hd%next\, \$19132_hd%now\, 
         \$17799_hd%next\, \$17799_hd%now\, \$v7067%next\, \$v7067%now\, 
         \$15138_v%next\, \$15138_v%now\, \$18284%next\, \$18284%now\, 
         \$14034_v%next\, \$14034_v%now\, \$18553%next\, \$18553%now\, 
         \$16725%next\, \$16725%now\, \$16381_v%next\, \$16381_v%now\, 
         \$14377_v%next\, \$14377_v%now\, \$16334_v%next\, \$16334_v%now\, 
         \$19076%next\, \$19076%now\, \$13972_v%next\, \$13972_v%now\, 
         \$13143_hd%next\, \$13143_hd%now\, \$19111%next\, \$19111%now\, 
         \$13684_hd%next\, \$13684_hd%now\, \$17562%next\, \$17562%now\, 
         \$17368_v%next\, \$17368_v%now\, \$18035_hd%next\, \$18035_hd%now\, 
         \$15747_v%next\, \$15747_v%now\, \$v7097%next\, \$v7097%now\, 
         \$15639_v%next\, \$15639_v%now\, \$v7149%next\, \$v7149%now\, 
         \$14103%next\, \$14103%now\, \$v7401%next\, \$v7401%now\, 
         \$v7037%next\, \$v7037%now\, \$14464_v%next\, \$14464_v%now\, 
         \$18180_hd%next\, \$18180_hd%now\, \$13787%next\, \$13787%now\, 
         \$v7157%next\, \$v7157%now\, \$13977_v%next\, \$13977_v%now\, 
         \$17952_w%next\, \$17952_w%now\, \$14185_next_env%next\, 
         \$14185_next_env%now\, \$16380_v%next\, \$16380_v%now\, 
         \$18030_w%next\, \$18030_w%now\, \$17183%next\, \$17183%now\, 
         \$18261%next\, \$18261%now\, \$14300_v%next\, \$14300_v%now\, 
         \$14512_v%next\, \$14512_v%now\, \$14898_v%next\, \$14898_v%now\, 
         \$14016_v%next\, \$14016_v%now\, \$v7047%next\, \$v7047%now\, 
         \$16074_v%next\, \$16074_v%now\, \$16709%next\, \$16709%now\, 
         \$v7127%next\, \$v7127%now\, \$13004_w%next\, \$13004_w%now\, 
         \$15711_v%next\, \$15711_v%now\, \$14423_v%next\, \$14423_v%now\, 
         \$14413_v%next\, \$14413_v%now\, \$18459_w%next\, \$18459_w%now\, 
         \$15545_v%next\, \$15545_v%now\, \$12929_hd%next\, \$12929_hd%now\, 
         \$13992_v%next\, \$13992_v%now\, \$18464_hd%next\, \$18464_hd%now\, 
         \$18701%next\, \$18701%now\, \$14446_v%next\, \$14446_v%now\, 
         \$18808%next\, \$18808%now\, \$19127_w%next\, \$19127_w%now\, 
         \$14578_v%next\, \$14578_v%now\, \$14043_v%next\, \$14043_v%now\, 
         \$15819_v%next\, \$15819_v%now\, \$17117_v%next\, \$17117_v%now\, 
         \$18335_w%next\, \$18335_w%now\, \$18175_w%next\, \$18175_w%now\, 
         \$17874_w%next\, \$17874_w%now\, \$17585_hd%next\, \$17585_hd%now\, 
         \$13605%next\, \$13605%now\, \$14165%next\, \$14165%now\, 
         \$14406_v%next\, \$14406_v%now\, \$19213%next\, \$19213%now\, 
         \$14738_v%next\, \$14738_v%now\, \$14070_v%next\, \$14070_v%now\, 
         \$16673_v%next\, \$16673_v%now\, \$16349_v%next\, \$16349_v%now\, 
         \$12553%next\, \$12553%now\, \$14139%next\, \$14139%now\, 
         \$17371_v%next\, \$17371_v%now\, \$15883%next\, \$15883%now\, 
         \$v7107%next\, \$v7107%now\, \$17749%next\, \$17749%now\, 
         \$17239_v%next\, \$17239_v%now\, \$13524_hd%next\, \$13524_hd%now\, 
         \$13223_hd%next\, \$13223_hd%now\, \$15861_v%next\, \$15861_v%now\, 
         \$v7117%next\, \$v7117%now\, \$16763_v%next\, \$16763_v%now\, 
         \$17535%next\, \$17535%now\, \$14463_v%next\, \$14463_v%now\, 
         \$15980_v%next\, \$15980_v%now\, \$14508_v%next\, \$14508_v%now\, 
         \$18443%next\, \$18443%now\, \$17374_v%next\, \$17374_v%now\, 
         \$18826_w%next\, \$18826_w%now\, \$17337%next\, \$17337%now\, 
         \$14092%next\, \$14092%now\, \$13009_hd%next\, \$13009_hd%now\, 
         \$14152%next\, \$14152%now\, \$12879%next\, \$12879%now\, 
         \$v7355%next\, \$v7355%now\, \$13765%next\, \$13765%now\, 
         \$v7399%next\, \$v7399%now\, \$12549%next\, \$12549%now\, 
         \$13379_hd%next\, \$13379_hd%now\, \$18124%next\, \$18124%now\, 
         \$14315_v%next\, \$14315_v%now\, \$18319%next\, \$18319%now\, 
         \$v7145%next\, \$v7145%now\, \$15897%next\, \$15897%now\, 
         \$16121_v%next\, \$16121_v%now\, \$13808_hd%next\, \$13808_hd%now\, 
         \$14221%next\, \$14221%now\, \$12924_w%next\, \$12924_w%now\, 
         \$17957_hd%next\, \$17957_hd%now\, \$12906%next\, \$12906%now\, 
         \$12546_dur%next\, \$12546_dur%now\, \$19251_w%next\, 
         \$19251_w%now\, \$19235%next\, \$19235%now\, \$13138_w%next\, 
         \$13138_w%now\, \$17879_hd%next\, \$17879_hd%now\, 
         \$14453_next_acc%next\, \$14453_next_acc%now\, \$17580_w%next\, 
         \$17580_w%now\, \$16630%next\, \$16630%now\, \$18724_hd%next\, 
         \$18724_hd%now\, \$16217_hd%next\, \$16217_hd%now\, \$15378_v%next\, 
         \$15378_v%now\, \$12538_cy%next\, \$12538_cy%now\, \$16379_v%next\, 
         \$16379_v%now\, \$v7398%next\, \$v7398%now\, \$14424_v%next\, 
         \$14424_v%now\, \$v7057%next\, \$v7057%now\, \$15981_v%next\, 
         \$15981_v%now\, \$16395_v%next\, \$16395_v%now\, \$18904_w%next\, 
         \$18904_w%now\, \$v7077%next\, \$v7077%now\, \$14285_v%next\, 
         \$14285_v%now\, \$14114%next\, \$14114%now\, \$16127_v%next\, 
         \$16127_v%now\, \$14658_v%next\, \$14658_v%now\, \$v7354%next\, 
         \$v7354%now\, \$16436_v%next\, \$16436_v%now\, \$14517_v%next\, 
         \$14517_v%now\, \$18982_w%next\, \$18982_w%now\, \$16439_v%next\, 
         \$16439_v%now\, \$14338_v%next\, \$14338_v%now\, \$15976_v%next\, 
         \$15976_v%now\, \$14818_v%next\, \$14818_v%now\, \$16042_v%next\, 
         \$16042_v%now\, \$v7400%next\, \$v7400%now\, \$13296_w%next\, 
         \$13296_w%now\, \$13301_hd%next\, \$13301_hd%now\, \$14330_v%next\, 
         \$14330_v%now\, \$15853_v%next\, \$15853_v%now\, \$v7017%next\, 
         \$v7017%now\, \$17250_v%next\, \$17250_v%now\, \$16713_v%next\, 
         \$16713_v%now\, \$17794_w%next\, \$17794_w%now\, \$13468%next\, 
         \$13468%now\, \$18831_hd%next\, \$18831_hd%now\, \$16438_v%next\, 
         \$16438_v%now\, \$15218_v%next\, \$15218_v%now\, \$18909_hd%next\, 
         \$18909_hd%now\, \$15298_v%next\, \$15298_v%now\, \$16037_v%next\, 
         \$16037_v%now\, \$15783_v%next\, \$15783_v%now\, \$14351_v%next\, 
         \$14351_v%now\, \$14177_hd%next\, \$14177_hd%now\, \$v7403%next\, 
         \$v7403%now\, \$15961%next\, \$15961%now\, \$18159%next\, 
         \$18159%now\, \$17665_hd%next\, \$17665_hd%now\, \$16169_v%next\, 
         \$16169_v%now\, \$17776%next\, \$17776%now\, \$13519_w%next\, 
         \$13519_w%now\, \$v7402%next\, \$v7402%now\, \$15932%next\, 
         \$15932%now\, \$13218_w%next\, \$13218_w%now\, \$13663%next\, 
         \$13663%now\, \$13679_w%next\, \$13679_w%now\, \$v7027%next\, 
         \$v7027%now\, \$16284_v%next\, \$16284_v%now\, \$14364_v%next\, 
         \$14364_v%now\, \$19337%next\, \$19337%now\, \$19256_hd%next\, 
         \$19256_hd%now\, \$13967_v%next\, \$13967_v%now\, \$v7161%next\, 
         \$v7161%now\, \$15058_v%next\, \$15058_v%now\, \$16729_v%next\, 
         \$16729_v%now\, \$14061_v%next\, \$14061_v%now\, \$14978_v%next\, 
         \$14978_v%now\, \$13997_v%next\, \$13997_v%now\, \$16299_v%next\, 
         \$16299_v%now\, \$v7137%next\, \$v7137%now\, \$16527_f0%next\, 
         \$16527_f0%now\, \$18987_hd%next\, \$18987_hd%now\, \$18719_w%next\, 
         \$18719_w%now\, \$13982_v%next\, \$13982_v%now\, \$16178_v%next\, 
         \$16178_v%now\, \$v7153%next\, \$v7153%now\, \$16453_v%next\, 
         \$16453_v%now\, \$14126%next\, \$14126%now\, \$13503%next\, 
         \$13503%now\, \$14052_v%next\, \$14052_v%now\, \$15675_v%next\, 
         \$15675_v%now\, \$18421%next\, \$18421%now\, \$14516_v%next\, 
         \$14516_v%now\ : value(0 to 31) := (others => '0');
  signal \$15364_binop_int6435910_result%next\, 
         \$15364_binop_int6435910_result%now\, 
         \$16551_compbranch6505926_result%next\, 
         \$16551_compbranch6505926_result%now\, 
         \$15733_binop_compare6455919_result%next\, 
         \$15733_binop_compare6455919_result%now\, 
         \$16858_compbranch6505932_result%next\, 
         \$16858_compbranch6505932_result%now\, 
         \$15124_binop_int6435907_result%next\, 
         \$15124_binop_int6435907_result%now\, 
         \$14884_binop_int6435904_result%next\, 
         \$14884_binop_int6435904_result%now\, 
         \$15769_binop_compare6455920_result%next\, 
         \$15769_binop_compare6455920_result%now\, 
         \$15531_binop_int6435913_result%next\, 
         \$15531_binop_int6435913_result%now\, 
         \$14964_binop_int6435905_result%next\, 
         \$14964_binop_int6435905_result%now\, 
         \$15805_binop_compare6455921_result%next\, 
         \$15805_binop_compare6455921_result%now\, 
         \$15451_binop_int6435912_result%next\, 
         \$15451_binop_int6435912_result%now\, 
         \$16788_compbranch6505930_result%next\, 
         \$16788_compbranch6505930_result%now\, 
         \$16963_compbranch6505935_result%next\, 
         \$16963_compbranch6505935_result%now\, 
         \$16589_compbranch6505927_result%next\, 
         \$16589_compbranch6505927_result%now\, 
         \$13925_offsetclosure_n639_result%next\, 
         \$13925_offsetclosure_n639_result%now\, 
         \$15044_binop_int6435906_result%next\, 
         \$15044_binop_int6435906_result%now\, \$13924_apply638_result%next\, 
         \$13924_apply638_result%now\, \$13926_make_block_n646_result%next\, 
         \$13926_make_block_n646_result%now\, 
         \$15661_binop_compare6455917_result%next\, 
         \$15661_binop_compare6455917_result%now\, 
         \$15284_binop_int6435909_result%next\, 
         \$15284_binop_int6435909_result%now\, 
         \$14804_binop_int6435903_result%next\, 
         \$14804_binop_int6435903_result%now\, 
         \$15204_binop_int6435908_result%next\, 
         \$15204_binop_int6435908_result%now\, 
         \$16928_compbranch6505934_result%next\, 
         \$16928_compbranch6505934_result%now\, 
         \$16823_compbranch6505931_result%next\, 
         \$16823_compbranch6505931_result%now\, 
         \$15625_binop_compare6455916_result%next\, 
         \$15625_binop_compare6455916_result%now\, 
         \$15697_binop_compare6455918_result%next\, 
         \$15697_binop_compare6455918_result%now\, \result6468%next\, 
         \result6468%now\, \$14644_binop_int6435901_result%next\, 
         \$14644_binop_int6435901_result%now\, 
         \$13927_branch_if648_result%next\, \$13927_branch_if648_result%now\, 
         \$16893_compbranch6505933_result%next\, 
         \$16893_compbranch6505933_result%now\, 
         \$14564_binop_int6435900_result%next\, 
         \$14564_binop_int6435900_result%now\, 
         \$14724_binop_int6435902_result%next\, 
         \$14724_binop_int6435902_result%now\ : value(0 to 121) := (others => '0');
  
  begin
    process (clk)
            begin
            if rising_edge(clk) then
                 if \$ram_write_request\ = '1' then
                    ram(\$ram_ptr_write\) <= \$ram_write\;
                 end if;
                 \$ram_value\ <= ram(\$ram_ptr\);
            end if;
        end process;
    
    process (clk)
            begin
            if rising_edge(clk) then
                 if \$global_end_write_request\ = '1' then
                    global_end(\$global_end_ptr_write\) <= \$global_end_write\;
                 end if;
                 \$global_end_value\ <= global_end(\$global_end_ptr\);
            end if;
        end process;
    
    process (clk)
            begin
            if rising_edge(clk) then
                 if \$code_write_request\ = '1' then
                    code(\$code_ptr_write\) <= \$code_write\;
                 end if;
                 \$code_value\ <= code(\$code_ptr\);
            end if;
        end process;
    
    process (reset,clk)
      begin
      if reset = '1' then
        \$12559%now\ <= (others => '0');
        \$14060%now\ <= (others => '0');
        \$v6454%now\ <= (others => '0');
        \$14516_v%now\ <= (others => '0');
        \$15069_modulo6685895_arg%now\ <= (others => '0');
        \$18421%now\ <= (others => '0');
        \$v6570%now\ <= (others => '0');
        \$14564_binop_int6435900_arg%now\ <= (others => '0');
        \$17813%now\ <= (others => '0');
        \$v6841%now\ <= (others => '0');
        \$14666_r%now\ <= (others => '0');
        \$v7022%now\ <= (others => '0');
        \$14589_modulo6685895_result%now\ <= (others => '0');
        \$13392%now\ <= (others => '0');
        \$18996%now\ <= (others => '0');
        \$12673_rdy%now\ <= (others => '0');
        \$v6130%now\ <= (others => '0');
        \$v7263%now\ <= (others => '0');
        \$14917_modulo6685888_arg%now\ <= (others => '0');
        \$v6197%now\ <= (others => '0');
        \$19272%now\ <= (others => '0');
        \$v7123%now\ <= (others => '0');
        \$v6642%now\ <= (others => '0');
        \$18729%now\ <= (others => '0');
        \$18192%now\ <= (others => '0');
        \$13670%now\ <= (others => '0');
        \$v6127%now\ <= (others => '0');
        \$15675_v%now\ <= (others => '0');
        \$15077_modulo6685888_result%now\ <= (others => '0');
        \$v6725%now\ <= (others => '0');
        \$16182%now\ <= (others => '0');
        \$14052_v%now\ <= (others => '0');
        \$18354%now\ <= (others => '0');
        \$14749_modulo6685895_result%now\ <= (others => '0');
        \$v6451%now\ <= (others => '0');
        \$12545_x%now\ <= (others => '0');
        \$v7062%now\ <= (others => '0');
        \$17496_next%now\ <= (others => '0');
        \$12852%now\ <= (others => '0');
        \$13503%now\ <= (others => '0');
        \$v6473%now\ <= (others => '0');
        \$15531_binop_int6435913_arg%now\ <= (others => '0');
        \$17887%now\ <= (others => '0');
        \$18997%now\ <= (others => '0');
        \$18835%now\ <= (others => '0');
        \$v6567%now\ <= (others => '0');
        \$v7313%now\ <= (others => '0');
        \$14724_binop_int6435902_result%now\ <= (others => '0');
        \$12699%now\ <= (others => '0');
        \$v7125%now\ <= (others => '0');
        \$14989_modulo6685895_arg%now\ <= (others => '0');
        \$13090%now\ <= (others => '0');
        \$19003%now\ <= (others => '0');
        \$12522_wait662_arg%now\ <= (others => '0');
        \$16811_compare6445898_arg%now\ <= (others => '0');
        \$17893%now\ <= (others => '0');
        \$15661_binop_compare6455917_arg%now\ <= (others => '0');
        \$14126%now\ <= (others => '0');
        \$v7437%now\ <= (others => '0');
        \$17570%now\ <= (others => '0');
        \$16453_v%now\ <= (others => '0');
        \$17676%now\ <= (others => '0');
        \$18121%now\ <= (others => '0');
        \$v7222%now\ <= (others => '0');
        \$v6512%now\ <= (others => '0');
        \$13308%now\ <= (others => '0');
        \$17018_w36575938_arg%now\ <= (others => '0');
        \$v6206%now\ <= (others => '0');
        \$15484_modulo6685888_result%now\ <= (others => '0');
        \$v7170%now\ <= (others => '0');
        \$15614_forever6705914_arg%now\ <= (others => '0');
        \$16858_compbranch6505932_arg%now\ <= (others => '0');
        \$v7236%now\ <= (others => '0');
        \$v7153%now\ <= (others => '0');
        \$16893_compbranch6505933_id%now\ <= (others => '0');
        \$14597_modulo6685888_arg%now\ <= (others => '0');
        \$16141%now\ <= (others => '0');
        \$v6105%now\ <= (others => '0');
        \$v7446%now\ <= (others => '0');
        \$13156%now\ <= (others => '0');
        \$v6575%now\ <= (others => '0');
        \$19138%now\ <= (others => '0');
        \$16178_v%now\ <= (others => '0');
        \$13945%now\ <= (others => '0');
        \$v7094%now\ <= (others => '0');
        \$v6391%now\ <= (others => '0');
        \$18838%now\ <= (others => '0');
        \$13824%now\ <= (others => '0');
        \$v6959%now\ <= (others => '0');
        \$13531%now\ <= (others => '0');
        \$16788_compbranch6505930_arg%now\ <= (others => '0');
        \$17971%now\ <= (others => '0');
        \$v6348%now\ <= (others => '0');
        \$17121%now\ <= (others => '0');
        \$16752_fill6545929_arg%now\ <= (others => '0');
        \$v6382%now\ <= (others => '0');
        \$12853_forever6705887_arg%now\ <= (others => '0');
        \$v7251%now\ <= (others => '0');
        \$15769_binop_compare6455920_arg%now\ <= (others => '0');
        \$17494%now\ <= (others => '0');
        \$v6385%now\ <= (others => '0');
        \$14326%now\ <= (others => '0');
        \$v6240%now\ <= (others => '0');
        \$19080_next%now\ <= (others => '0');
        \$17386%now\ <= (others => '0');
        \$13982_v%now\ <= (others => '0');
        \$17459_loop665_arg%now\ <= (others => '0');
        \$18719_w%now\ <= (others => '0');
        \$15445%now\ <= (others => '0');
        \$v7353%now\ <= (others => '0');
        \$16752_fill6545929_result%now\ <= (others => '0');
        \$14997_modulo6685888_id%now\ <= (others => '0');
        \$18050%now\ <= (others => '0');
        \$12883%now\ <= (others => '0');
        \$16823_compbranch6505931_arg%now\ <= (others => '0');
        \$16233%now\ <= (others => '0');
        \$16271%now\ <= (others => '0');
        \$12682_make_block579_arg%now\ <= (others => '0');
        \$18655%now\ <= (others => '0');
        \$v7371%now\ <= (others => '0');
        \$18987_hd%now\ <= (others => '0');
        \$v6619%now\ <= (others => '0');
        \$v6427%now\ <= (others => '0');
        \$16748%now\ <= (others => '0');
        \$v6974%now\ <= (others => '0');
        \$18474%now\ <= (others => '0');
        \$17886%now\ <= (others => '0');
        \$15756_compare6445897_arg%now\ <= (others => '0');
        \$13151%now\ <= (others => '0');
        \$v6805%now\ <= (others => '0');
        \$17569%now\ <= (others => '0');
        \$12698%now\ <= (others => '0');
        \$15389_modulo6685895_arg%now\ <= (others => '0');
        \$v6035%now\ <= (others => '0');
        \$15553_r%now\ <= (others => '0');
        \$15237_modulo6685888_result%now\ <= (others => '0');
        \$12944%now\ <= (others => '0');
        \$14613_modulo6685896_result%now\ <= (others => '0');
        \$v7381%now\ <= (others => '0');
        \$18846%now\ <= (others => '0');
        \$18917%now\ <= (others => '0');
        \$v6092%now\ <= (others => '0');
        \$18916%now\ <= (others => '0');
        \$15261_modulo6685888_id%now\ <= (others => '0');
        \$17679%now\ <= (others => '0');
        \$13154%now\ <= (others => '0');
        \$v6336%now\ <= (others => '0');
        \$16527_f0%now\ <= (others => '0');
        \$18352%now\ <= (others => '0');
        \$13964%now\ <= (others => '0');
        \$v7420%now\ <= (others => '0');
        \$13632_next%now\ <= (others => '0');
        \$v6502%now\ <= (others => '0');
        \$v6370%now\ <= (others => '0');
        \$18739%now\ <= (others => '0');
        \$12714%now\ <= (others => '0');
        \$17484%now\ <= (others => '0');
        \$17597%now\ <= (others => '0');
        \$15756_compare6445897_result%now\ <= (others => '0');
        \$v7137%now\ <= (others => '0');
        \$13532%now\ <= (others => '0');
        \$v6823%now\ <= (others => '0');
        \$14781_modulo6685888_result%now\ <= (others => '0');
        \$v6721%now\ <= (others => '0');
        \$17734_copy_root_in_ram6635892_id%now\ <= (others => '0');
        \$v7338%now\ <= (others => '0');
        \$14749_modulo6685895_arg%now\ <= (others => '0');
        \$v7050%now\ <= (others => '0');
        \$16299_v%now\ <= (others => '0');
        \$12689%now\ <= (others => '0');
        \$18807%now\ <= (others => '0');
        \$13920_loop666_arg%now\ <= (others => '0');
        \$17455_loop666_id%now\ <= (others => '0');
        \$v6027%now\ <= (others => '0');
        \$18650%now\ <= (others => '0');
        \$18837%now\ <= (others => '0');
        \$16951_compare6445898_arg%now\ <= (others => '0');
        \$14861_modulo6685888_result%now\ <= (others => '0');
        \$18805%now\ <= (others => '0');
        \$17543%now\ <= (others => '0');
        \$13997_v%now\ <= (others => '0');
        \$16574_compare6445898_id%now\ <= (others => '0');
        \$v6728%now\ <= (others => '0');
        \$v6500%now\ <= (others => '0');
        \$v5869%now\ <= (others => '0');
        \$v6496%now\ <= (others => '0');
        \$14978_v%now\ <= (others => '0');
        \$v7454%now\ <= (others => '0');
        \$13237%now\ <= (others => '0');
        \$v6146%now\ <= (others => '0');
        \$15330_r%now\ <= (others => '0');
        \$12839%now\ <= (others => '0');
        \$14061_v%now\ <= (others => '0');
        \$14701_modulo6685888_arg%now\ <= (others => '0');
        \$12697%now\ <= (others => '0');
        \$17773%now\ <= (others => '0');
        \$v7344%now\ <= (others => '0');
        \$12888%now\ <= (others => '0');
        \$13155%now\ <= (others => '0');
        \$12937%now\ <= (others => '0');
        \$16115%now\ <= (others => '0');
        \$12805_aux664_result%now\ <= (others => '0');
        \$v6021%now\ <= (others => '0');
        \$13697%now\ <= (others => '0');
        \$v6466%now\ <= (others => '0');
        \$18355%now\ <= (others => '0');
        \rdy5940%now\ <= (others => '0');
        \$13102%now\ <= (others => '0');
        \$13235%now\ <= (others => '0');
        \$15044_binop_int6435906_id%now\ <= (others => '0');
        \$16729_v%now\ <= (others => '0');
        \$v6376%now\ <= (others => '0');
        \$13233%now\ <= (others => '0');
        \$17670%now\ <= (others => '0');
        \$14555%now\ <= (others => '0');
        \$14564_binop_int6435900_result%now\ <= (others => '0');
        \$v6802%now\ <= (others => '0');
        \$15058_v%now\ <= (others => '0');
        \$17464%now\ <= (others => '0');
        \$v6599%now\ <= (others => '0');
        \$v6430%now\ <= (others => '0');
        \$v6318%now\ <= (others => '0');
        \$v7161%now\ <= (others => '0');
        \$17669%now\ <= (others => '0');
        \$16963_compbranch6505935_id%now\ <= (others => '0');
        \$13967_v%now\ <= (others => '0');
        \$13696%now\ <= (others => '0');
        \$v6015%now\ <= (others => '0');
        \$15476_modulo6685895_arg%now\ <= (others => '0');
        \$17470%now\ <= (others => '0');
        \$12520_loop666_id%now\ <= (others => '0');
        \$18815%now\ <= (others => '0');
        \$v6559%now\ <= (others => '0');
        \$18565%now\ <= (others => '0');
        \$16551_compbranch6505926_id%now\ <= (others => '0');
        \$15397_modulo6685888_result%now\ <= (others => '0');
        \$12877%now\ <= (others => '0');
        \$18698%now\ <= (others => '0');
        \$18480%now\ <= (others => '0');
        \$v7300%now\ <= (others => '0');
        \$15389_modulo6685895_result%now\ <= (others => '0');
        \$v7144%now\ <= (others => '0');
        \$v6780%now\ <= (others => '0');
        \$19256_hd%now\ <= (others => '0');
        \$15823_res%now\ <= (others => '0');
        \$15124_binop_int6435907_id%now\ <= (others => '0');
        \$v6218%now\ <= (others => '0');
        \$v7406%now\ <= (others => '0');
        \$16963_compbranch6505935_arg%now\ <= (others => '0');
        \$v7132%now\ <= (others => '0');
        \$v7200%now\ <= (others => '0');
        \$18633_loop665_id%now\ <= (others => '0');
        \$17888%now\ <= (others => '0');
        \$19145%now\ <= (others => '0');
        \$15625_binop_compare6455916_id%now\ <= (others => '0');
        \$19337%now\ <= (others => '0');
        \$15893%now\ <= (others => '0');
        \$14364_v%now\ <= (others => '0');
        \$16893_compbranch6505933_result%now\ <= (others => '0');
        \$v6406%now\ <= (others => '0');
        \$v6489%now\ <= (others => '0');
        \$14837_modulo6685888_result%now\ <= (others => '0');
        \$14677_modulo6685888_arg%now\ <= (others => '0');
        \$v6667%now\ <= (others => '0');
        \$v7413%now\ <= (others => '0');
        \$v6508%now\ <= (others => '0');
        \$v6591%now\ <= (others => '0');
        \$16284_v%now\ <= (others => '0');
        \$12808_aux664_result%now\ <= (others => '0');
        \$13816%now\ <= (others => '0');
        \$v6211%now\ <= (others => '0');
        \$15874%now\ <= (others => '0');
        \$14829_modulo6685895_id%now\ <= (others => '0');
        \$v7027%now\ <= (others => '0');
        \$v6596%now\ <= (others => '0');
        \$17746%now\ <= (others => '0');
        \$13950%now\ <= (others => '0');
        \$v5963%now\ <= (others => '0');
        \$v5944%now\ <= (others => '0');
        \$14597_modulo6685888_result%now\ <= (others => '0');
        \$14582_res%now\ <= (others => '0');
        \$17891%now\ <= (others => '0');
        \$15397_modulo6685888_arg%now\ <= (others => '0');
        \$13927_branch_if648_result%now\ <= (others => '0');
        \$v7306%now\ <= (others => '0');
        \$v7074%now\ <= (others => '0');
        \$15021_modulo6685888_result%now\ <= (others => '0');
        \$12707%now\ <= (others => '0');
        \$16881_compare6445898_result%now\ <= (others => '0');
        \$13679_w%now\ <= (others => '0');
        \$13663%now\ <= (others => '0');
        \$18447%now\ <= (others => '0');
        \$v6732%now\ <= (others => '0');
        \$v6298%now\ <= (others => '0');
        \$v6518%now\ <= (others => '0');
        \$18278%now\ <= (others => '0');
        \$12544%now\ <= (others => '0');
        \$13218_w%now\ <= (others => '0');
        \$15932%now\ <= (others => '0');
        \$v7402%now\ <= (others => '0');
        \$v7085%now\ <= (others => '0');
        \$18731%now\ <= (others => '0');
        \$13519_w%now\ <= (others => '0');
        \$13606%now\ <= (others => '0');
        \$17776%now\ <= (others => '0');
        \$18644%now\ <= (others => '0');
        \$16327%now\ <= (others => '0');
        \$16169_v%now\ <= (others => '0');
        \$16551_compbranch6505926_arg%now\ <= (others => '0');
        \$15229_modulo6685895_arg%now\ <= (others => '0');
        \$17457_aux664_result%now\ <= (others => '0');
        \$v6633%now\ <= (others => '0');
        \$17665_hd%now\ <= (others => '0');
        \$18159%now\ <= (others => '0');
        \$v6058%now\ <= (others => '0');
        \$14122%now\ <= (others => '0');
        \$18563%now\ <= (others => '0');
        \$13310%now\ <= (others => '0');
        \$14012%now\ <= (others => '0');
        \$14677_modulo6685888_id%now\ <= (others => '0');
        \$14181_sp%now\ <= (others => '0');
        \$v6235%now\ <= (others => '0');
        \$15961%now\ <= (others => '0');
        \$15476_modulo6685895_result%now\ <= (others => '0');
        \$15237_modulo6685888_id%now\ <= (others => '0');
        \$17505_forever6705894_arg%now\ <= (others => '0');
        \$13388%now\ <= (others => '0');
        \$v6480%now\ <= (others => '0');
        \$17001%now\ <= (others => '0');
        \$17963%now\ <= (others => '0');
        \$17803%now\ <= (others => '0');
        \$19142%now\ <= (others => '0');
        \$18679_forever6705881_id%now\ <= (others => '0');
        \$v6291%now\ <= (others => '0');
        \$v6532%now\ <= (others => '0');
        \$v7293%now\ <= (others => '0');
        \$18919%now\ <= (others => '0');
        \$12685%now\ <= (others => '0');
        \$v6501%now\ <= (others => '0');
        \$17238_sp%now\ <= (others => '0');
        \$18186%now\ <= (others => '0');
        \$v7279%now\ <= (others => '0');
        \$v6460%now\ <= (others => '0');
        \$14431%now\ <= (others => '0');
        \$13667%now\ <= (others => '0');
        \$17455_loop666_arg%now\ <= (others => '0');
        \$12851%now\ <= (others => '0');
        \$18188%now\ <= (others => '0');
        \$v6172%now\ <= (others => '0');
        \$v7403%now\ <= (others => '0');
        \$v7216%now\ <= (others => '0');
        \$v7035%now\ <= (others => '0');
        \$v6397%now\ <= (others => '0');
        \$18709%now\ <= (others => '0');
        \$15720_compare6445897_id%now\ <= (others => '0');
        \$13823%now\ <= (others => '0');
        \$14177_hd%now\ <= (others => '0');
        \result6503%now\ <= (others => '0');
        \$13395%now\ <= (others => '0');
        \$16353%now\ <= (others => '0');
        \$v6239%now\ <= (others => '0');
        \$17559%now\ <= (others => '0');
        \$14351_v%now\ <= (others => '0');
        \$12808_aux664_id%now\ <= (others => '0');
        \$19269%now\ <= (others => '0');
        \$17412%now\ <= (others => '0');
        \$v7007%now\ <= (others => '0');
        \$v6941%now\ <= (others => '0');
        \$v6746%now\ <= (others => '0');
        \$18925%now\ <= (others => '0');
        \$v6838%now\ <= (others => '0');
        \$18733%now\ <= (others => '0');
        \$v5957%now\ <= (others => '0');
        \$v6953%now\ <= (others => '0');
        \$15783_v%now\ <= (others => '0');
        \$18279%now\ <= (others => '0');
        \$14207_loop_push6495899_result%now\ <= (others => '0');
        \$v6108%now\ <= (others => '0');
        \$v7025%now\ <= (others => '0');
        \$18120%now\ <= (others => '0');
        \$18566%now\ <= (others => '0');
        \$13016%now\ <= (others => '0');
        \$v6304%now\ <= (others => '0');
        \$12692%now\ <= (others => '0');
        \$16037_v%now\ <= (others => '0');
        \$12935%now\ <= (others => '0');
        \$13625%now\ <= (others => '0');
        \$v7434%now\ <= (others => '0');
        \$v6739%now\ <= (others => '0');
        \$17509_forever6705890_arg%now\ <= (others => '0');
        \$v6274%now\ <= (others => '0');
        \$19001%now\ <= (others => '0');
        \$v7290%now\ <= (others => '0');
        \$17498%now\ <= (others => '0');
        \$16945_b%now\ <= (others => '0');
        \$15298_v%now\ <= (others => '0');
        \$18346%now\ <= (others => '0');
        \$16589_compbranch6505927_id%now\ <= (others => '0');
        \$v6708%now\ <= (others => '0');
        \$13157%now\ <= (others => '0');
        \$18909_hd%now\ <= (others => '0');
        \$17674%now\ <= (others => '0');
        \$12712%now\ <= (others => '0');
        \$12945%now\ <= (others => '0');
        \$17354%now\ <= (others => '0');
        \$16574_compare6445898_result%now\ <= (others => '0');
        \$16365%now\ <= (others => '0');
        \$12715%now\ <= (others => '0');
        \$16510_forever6705925_id%now\ <= (others => '0');
        \$15218_v%now\ <= (others => '0');
        \$18699%now\ <= (others => '0');
        \$17591%now\ <= (others => '0');
        \$v6627%now\ <= (others => '0');
        \$12915%now\ <= (others => '0');
        \$v6136%now\ <= (others => '0');
        \$18045%now\ <= (others => '0');
        \$17460_aux664_id%now\ <= (others => '0');
        \$12807_loop665_id%now\ <= (others => '0');
        \$15069_modulo6685895_id%now\ <= (others => '0');
        \$v6492%now\ <= (others => '0');
        \$17487%now\ <= (others => '0');
        \$v6892%now\ <= (others => '0');
        \$17387%now\ <= (others => '0');
        \$15386_r%now\ <= (others => '0');
        \$v6729%now\ <= (others => '0');
        \$v6914%now\ <= (others => '0');
        \$18915%now\ <= (others => '0');
        \$17105_w06555936_id%now\ <= (others => '0');
        \$16589_compbranch6505927_arg%now\ <= (others => '0');
        \$13890%now\ <= (others => '0');
        \$19144%now\ <= (others => '0');
        \$16677%now\ <= (others => '0');
        \$v7034%now\ <= (others => '0');
        \$17678%now\ <= (others => '0');
        \$16875_b%now\ <= (others => '0');
        \$13927_branch_if648_arg%now\ <= (others => '0');
        \$v6883%now\ <= (others => '0');
        \$16438_v%now\ <= (others => '0');
        \$15612%now\ <= (others => '0');
        \$14773_modulo6685896_arg%now\ <= (others => '0');
        \$19140%now\ <= (others => '0');
        \$19071%now\ <= (others => '0');
        \$12848%now\ <= (others => '0');
        \$18831_hd%now\ <= (others => '0');
        \$v6710%now\ <= (others => '0');
        \$13468%now\ <= (others => '0');
        \$v6856%now\ <= (others => '0');
        \$15317_modulo6685888_result%now\ <= (others => '0');
        \$18570%now\ <= (others => '0');
        \$13623%now\ <= (others => '0');
        \$18128_next%now\ <= (others => '0');
        \$v7248%now\ <= (others => '0');
        \$14644_binop_int6435901_result%now\ <= (others => '0');
        \$12679_loop666_id%now\ <= (others => '0');
        \$16399%now\ <= (others => '0');
        \$19263%now\ <= (others => '0');
        \$14749_modulo6685895_id%now\ <= (others => '0');
        \$17794_w%now\ <= (others => '0');
        \result6468%now\ <= (others => '0');
        \$v7045%now\ <= (others => '0');
        \$18816%now\ <= (others => '0');
        \$17885%now\ <= (others => '0');
        \$v7164%now\ <= (others => '0');
        \$15101_modulo6685888_result%now\ <= (others => '0');
        \$v7042%now\ <= (others => '0');
        \$15500_modulo6685896_arg%now\ <= (others => '0');
        \$15333_modulo6685896_result%now\ <= (others => '0');
        \$17761_copy_root_in_ram6635891_result%now\ <= (others => '0');
        \$15720_compare6445897_arg%now\ <= (others => '0');
        \$16713_v%now\ <= (others => '0');
        \$15697_binop_compare6455918_arg%now\ <= (others => '0');
        \$17250_v%now\ <= (others => '0');
        \$12887%now\ <= (others => '0');
        \$v6826%now\ <= (others => '0');
        \$17394%now\ <= (others => '0');
        \$v6695%now\ <= (others => '0');
        \$17333_sp%now\ <= (others => '0');
        \$v7017%now\ <= (others => '0');
        \$16158_forever6705923_arg%now\ <= (others => '0');
        \$v6874%now\ <= (others => '0');
        \$v6574%now\ <= (others => '0');
        \$15853_v%now\ <= (others => '0');
        \$v7372%now\ <= (others => '0');
        \$v6651%now\ <= (others => '0');
        \$v7013%now\ <= (others => '0');
        \$15181_modulo6685888_result%now\ <= (others => '0');
        \$12691%now\ <= (others => '0');
        \$17962%now\ <= (others => '0');
        \$v6367%now\ <= (others => '0');
        \$v6200%now\ <= (others => '0');
        \$16612_compare6445898_result%now\ <= (others => '0');
        \$v6688%now\ <= (others => '0');
        \$14330_v%now\ <= (others => '0');
        \$v7361%now\ <= (others => '0');
        \$17319%now\ <= (others => '0');
        \$13941%now\ <= (others => '0');
        \$16078%now\ <= (others => '0');
        \$16165%now\ <= (others => '0');
        \$v7299%now\ <= (others => '0');
        \$17012_sp%now\ <= (others => '0');
        \$15261_modulo6685888_arg%now\ <= (others => '0');
        \$v6342%now\ <= (others => '0');
        \$v5954%now\ <= (others => '0');
        \$16606_b%now\ <= (others => '0');
        \$14986_r%now\ <= (others => '0');
        \$13301_hd%now\ <= (others => '0');
        \$15847%now\ <= (others => '0');
        \$v7179%now\ <= (others => '0');
        \$15021_modulo6685888_arg%now\ <= (others => '0');
        \$13127%now\ <= (others => '0');
        \$v7004%now\ <= (others => '0');
        \$v7090%now\ <= (others => '0');
        \$v6709%now\ <= (others => '0');
        \$17321%now\ <= (others => '0');
        \$13530%now\ <= (others => '0');
        \$14222%now\ <= (others => '0');
        \$v6868%now\ <= (others => '0');
        \$v6203%now\ <= (others => '0');
        \$v5866%now\ <= (others => '0');
        \$v5951%now\ <= (others => '0');
        \$18450%now\ <= (others => '0');
        \$13296_w%now\ <= (others => '0');
        \$14724_binop_int6435902_id%now\ <= (others => '0');
        \$v7400%now\ <= (others => '0');
        \$13013%now\ <= (others => '0');
        \$17349%now\ <= (others => '0');
        \$16192%now\ <= (others => '0');
        \$12834%now\ <= (others => '0');
        \$16441%now\ <= (others => '0');
        \$17167%now\ <= (others => '0');
        \$16042_v%now\ <= (others => '0');
        \$15697_binop_compare6455918_result%now\ <= (others => '0');
        \$12679_loop666_result%now\ <= (others => '0');
        \$16234%now\ <= (others => '0');
        \$15625_binop_compare6455916_result%now\ <= (others => '0');
        \$v7140%now\ <= (others => '0');
        \$18163%now\ <= (others => '0');
        \$v6007%now\ <= (others => '0');
        \$14933_modulo6685896_result%now\ <= (others => '0');
        \$v7066%now\ <= (others => '0');
        \$14818_v%now\ <= (others => '0');
        \$v6750%now\ <= (others => '0');
        \$15976_v%now\ <= (others => '0');
        \$v6935%now\ <= (others => '0');
        \$14338_v%now\ <= (others => '0');
        \$v6986%now\ <= (others => '0');
        \$16805_b%now\ <= (others => '0');
        \$17961%now\ <= (others => '0');
        \$16439_v%now\ <= (others => '0');
        \$14933_modulo6685896_id%now\ <= (others => '0');
        \$17681%now\ <= (others => '0');
        \$12910%now\ <= (others => '0');
        \$v6445%now\ <= (others => '0');
        \$12741%now\ <= (others => '0');
        \$v7455%now\ <= (others => '0');
        \$v6277%now\ <= (others => '0');
        \$v6962%now\ <= (others => '0');
        \$v7441%now\ <= (others => '0');
        \$13962%now\ <= (others => '0');
        \$15010_r%now\ <= (others => '0');
        \$14829_modulo6685895_result%now\ <= (others => '0');
        \$12521_loop665_arg%now\ <= (others => '0');
        \$14161%now\ <= (others => '0');
        \$15805_binop_compare6455921_arg%now\ <= (others => '0');
        \$12843%now\ <= (others => '0');
        \$15413_modulo6685896_result%now\ <= (others => '0');
        \$v7064%now\ <= (others => '0');
        \$15484_modulo6685888_arg%now\ <= (others => '0');
        \$v7368%now\ <= (others => '0');
        \$v6117%now\ <= (others => '0');
        \$18634_aux664_result%now\ <= (others => '0');
        \$12943%now\ <= (others => '0');
        \$v6995%now\ <= (others => '0');
        \$v6657%now\ <= (others => '0');
        \$17600%now\ <= (others => '0');
        \$v6214%now\ <= (others => '0');
        \$13957%now\ <= (others => '0');
        \$v7016%now\ <= (others => '0');
        \$v6307%now\ <= (others => '0');
        \$v6268%now\ <= (others => '0');
        \$18982_w%now\ <= (others => '0');
        \$13103%now\ <= (others => '0');
        \$14517_v%now\ <= (others => '0');
        \$v7023%now\ <= (others => '0');
        \$13692%now\ <= (others => '0');
        \$18479%now\ <= (others => '0');
        \$v7358%now\ <= (others => '0');
        \$v6271%now\ <= (others => '0');
        \$v6681%now\ <= (others => '0');
        \$12806_loop666_result%now\ <= (others => '0');
        \$12680_loop665_result%now\ <= (others => '0');
        \$18734%now\ <= (others => '0');
        \$15484_modulo6685888_id%now\ <= (others => '0');
        \$v6055%now\ <= (others => '0');
        \$14746_r%now\ <= (others => '0');
        \$17327%now\ <= (others => '0');
        \$13153%now\ <= (others => '0');
        \$v6701%now\ <= (others => '0');
        \$v7453%now\ <= (others => '0');
        \$v6950%now\ <= (others => '0');
        \$15733_binop_compare6455919_arg%now\ <= (others => '0');
        \$16436_v%now\ <= (others => '0');
        \$v7335%now\ <= (others => '0');
        \$14837_modulo6685888_arg%now\ <= (others => '0');
        \$14558%now\ <= (others => '0');
        \$v6609%now\ <= (others => '0');
        \$v6102%now\ <= (others => '0');
        \$v6865%now\ <= (others => '0');
        \$v7121%now\ <= (others => '0');
        \$v6175%now\ <= (others => '0');
        \$17520_copy_root_in_ram6635893_id%now\ <= (others => '0');
        \$18818%now\ <= (others => '0');
        \$17018_w36575938_id%now\ <= (others => '0');
        \$13946%now\ <= (others => '0');
        \$v7354%now\ <= (others => '0');
        \$17315%now\ <= (others => '0');
        \$15204_binop_int6435908_id%now\ <= (others => '0');
        \$14658_v%now\ <= (others => '0');
        \$13307%now\ <= (others => '0');
        \$14042%now\ <= (others => '0');
        \$12939%now\ <= (others => '0');
        \$12891_copy_root_in_ram6635884_arg%now\ <= (others => '0');
        \$v7416%now\ <= (others => '0');
        \$18166%now\ <= (others => '0');
        \$15556_modulo6685895_result%now\ <= (others => '0');
        \$16035%now\ <= (others => '0');
        \$14853_modulo6685896_arg%now\ <= (others => '0');
        \$15124_binop_int6435907_arg%now\ <= (others => '0');
        \$13928_w652_result%now\ <= (others => '0');
        \$15317_modulo6685888_arg%now\ <= (others => '0');
        \$17377%now\ <= (others => '0');
        \$16126%now\ <= (others => '0');
        \$v7133%now\ <= (others => '0');
        \$16127_v%now\ <= (others => '0');
        \$12878%now\ <= (others => '0');
        \$16031%now\ <= (others => '0');
        \$18836%now\ <= (others => '0');
        \$12857_forever6705883_arg%now\ <= (others => '0');
        \$v7219%now\ <= (others => '0');
        \$v6773%now\ <= (others => '0');
        \$14114%now\ <= (others => '0');
        \$v7086%now\ <= (others => '0');
        \$18999%now\ <= (others => '0');
        \$18637%now\ <= (others => '0');
        \$v6301%now\ <= (others => '0');
        \$17734_copy_root_in_ram6635892_arg%now\ <= (others => '0');
        \$v5874%now\ <= (others => '0');
        \$v7185%now\ <= (others => '0');
        \$13693%now\ <= (others => '0');
        \$v6229%now\ <= (others => '0');
        \$14285_v%now\ <= (others => '0');
        \$12734%now\ <= (others => '0');
        \$15341_modulo6685888_arg%now\ <= (others => '0');
        \$12904%now\ <= (others => '0');
        \$v7077%now\ <= (others => '0');
        \$17513_forever6705889_id%now\ <= (others => '0');
        \$v6853%now\ <= (others => '0');
        \$13466%now\ <= (others => '0');
        \$v7322%now\ <= (others => '0');
        \$14804_binop_int6435903_arg%now\ <= (others => '0');
        \$17463%now\ <= (others => '0');
        \$19115%now\ <= (others => '0');
        \$18904_w%now\ <= (others => '0');
        \$12818%now\ <= (others => '0');
        \$v6751%now\ <= (others => '0');
        \$16292%now\ <= (others => '0');
        \$12844_next%now\ <= (others => '0');
        \$16395_v%now\ <= (others => '0');
        \$14964_binop_int6435905_id%now\ <= (others => '0');
        \$16767%now\ <= (others => '0');
        \$15093_modulo6685896_arg%now\ <= (others => '0');
        \$v6103%now\ <= (others => '0');
        \$15648_compare6445897_id%now\ <= (others => '0');
        \$v6165%now\ <= (others => '0');
        \$18104%now\ <= (others => '0');
        \$v7030%now\ <= (others => '0');
        \$14613_modulo6685896_id%now\ <= (others => '0');
        \$v6738%now\ <= (others => '0');
        \$v6678%now\ <= (others => '0');
        \$17491%now\ <= (others => '0');
        \$13078_copy_root_in_ram6635885_id%now\ <= (others => '0');
        \$15981_v%now\ <= (others => '0');
        \$12560%now\ <= (others => '0');
        \$v7057%now\ <= (others => '0');
        \$v6364%now\ <= (others => '0');
        \$12702%now\ <= (others => '0');
        \$13312%now\ <= (others => '0');
        \$12520_loop666_arg%now\ <= (others => '0');
        \$15792_compare6445897_result%now\ <= (others => '0');
        \$15341_modulo6685888_result%now\ <= (others => '0');
        \$v7076%now\ <= (others => '0');
        \$14669_modulo6685895_id%now\ <= (others => '0');
        \$v5878%now\ <= (others => '0');
        \$18711%now\ <= (others => '0');
        \$15828_compare6445897_id%now\ <= (others => '0');
        \$15237_modulo6685888_arg%now\ <= (others => '0');
        \$v6183%now\ <= (others => '0');
        \$v5992%now\ <= (others => '0');
        \$v6314%now\ <= (others => '0');
        \$12522_wait662_result%now\ <= (others => '0');
        \$v6947%now\ <= (others => '0');
        \$v6595%now\ <= (others => '0');
        \$17455_loop666_result%now\ <= (others => '0');
        \$v7458%now\ <= (others => '0');
        \$v6162%now\ <= (others => '0');
        \$12838_next%now\ <= (others => '0');
        \$v6012%now\ <= (others => '0');
        \$18472%now\ <= (others => '0');
        \$16036_sp%now\ <= (others => '0');
        \$18185%now\ <= (others => '0');
        \$14424_v%now\ <= (others => '0');
        \$14254%now\ <= (others => '0');
        \$13389%now\ <= (others => '0');
        \$18677%now\ <= (others => '0');
        \$17348%now\ <= (others => '0');
        \$13393%now\ <= (others => '0');
        \$15769_binop_compare6455920_id%now\ <= (others => '0');
        \$13387%now\ <= (others => '0');
        \$17590%now\ <= (others => '0');
        \$v7398%now\ <= (others => '0');
        \$16823_compbranch6505931_id%now\ <= (others => '0');
        \$17495%now\ <= (others => '0');
        \$16379_v%now\ <= (others => '0');
        \$16881_compare6445898_arg%now\ <= (others => '0');
        \$18679_forever6705881_arg%now\ <= (others => '0');
        \$v6048%now\ <= (others => '0');
        \$14677_modulo6685888_result%now\ <= (others => '0');
        \$18288_next%now\ <= (others => '0');
        \$12538_cy%now\ <= (others => '0');
        \$15378_v%now\ <= (others => '0');
        \$12941%now\ <= (others => '0');
        \$17783%now\ <= (others => '0');
        \$13794%now\ <= (others => '0');
        \$14693_modulo6685896_arg%now\ <= (others => '0');
        \$12914%now\ <= (others => '0');
        \$19262%now\ <= (others => '0');
        \$v6847%now\ <= (others => '0');
        \$15382_res%now\ <= (others => '0');
        \$12521_loop665_result%now\ <= (others => '0');
        \$13238%now\ <= (others => '0');
        \$v6286%now\ <= (others => '0');
        \$19070%now\ <= (others => '0');
        \$17254%now\ <= (others => '0');
        \$13694%now\ <= (others => '0');
        \$14941_modulo6685888_arg%now\ <= (others => '0');
        \$v7328%now\ <= (others => '0');
        \$18356%now\ <= (others => '0');
        \$v7054%now\ <= (others => '0');
        \$17761_copy_root_in_ram6635891_id%now\ <= (others => '0');
        \$12695%now\ <= (others => '0');
        \$v6089%now\ <= (others => '0');
        \$17774%now\ <= (others => '0');
        \$16231%now\ <= (others => '0');
        \$v7015%now\ <= (others => '0');
        \$16202_ofs%now\ <= (others => '0');
        \$v7091%now\ <= (others => '0');
        \$16217_hd%now\ <= (others => '0');
        \$v6400%now\ <= (others => '0');
        \$v6388%now\ <= (others => '0');
        \$16024%now\ <= (others => '0');
        \$12913%now\ <= (others => '0');
        \$17048_w16565937_arg%now\ <= (others => '0');
        \$15476_modulo6685895_id%now\ <= (others => '0');
        \$16823_compbranch6505931_result%now\ <= (others => '0');
        \$16928_compbranch6505934_result%now\ <= (others => '0');
        \$18475%now\ <= (others => '0');
        \$17890%now\ <= (others => '0');
        \$15580_modulo6685896_id%now\ <= (others => '0');
        \$15828_compare6445897_result%now\ <= (others => '0');
        \$12936%now\ <= (others => '0');
        \$17165%now\ <= (others => '0');
        \$12660%now\ <= (others => '0');
        \$v7232%now\ <= (others => '0');
        \$12736%now\ <= (others => '0');
        \$v6724%now\ <= (others => '0');
        \$18724_hd%now\ <= (others => '0');
        \$17775%now\ <= (others => '0');
        \$16630%now\ <= (others => '0');
        \$15341_modulo6685888_id%now\ <= (others => '0');
        \$18187%now\ <= (others => '0');
        \$v6998%now\ <= (others => '0');
        \$17580_w%now\ <= (others => '0');
        \$17785%now\ <= (others => '0');
        \$12716%now\ <= (others => '0');
        \$15253_modulo6685896_id%now\ <= (others => '0');
        \$14135%now\ <= (others => '0');
        \$15828_compare6445897_arg%now\ <= (others => '0');
        \$13129%now\ <= (others => '0');
        \$18194%now\ <= (others => '0');
        \$18193%now\ <= (others => '0');
        \$16916_compare6445898_arg%now\ <= (others => '0');
        \$17812%now\ <= (others => '0');
        \$12806_loop666_id%now\ <= (others => '0');
        \$15204_binop_int6435908_result%now\ <= (others => '0');
        \$v7210%now\ <= (others => '0');
        \$17457_aux664_arg%now\ <= (others => '0');
        \$14453_next_acc%now\ <= (others => '0');
        \$18571%now\ <= (others => '0');
        \$15309_modulo6685895_result%now\ <= (others => '0');
        \$17879_hd%now\ <= (others => '0');
        \$13138_w%now\ <= (others => '0');
        \$v6624%now\ <= (others => '0');
        \$v6992%now\ <= (others => '0');
        \$14644_binop_int6435901_arg%now\ <= (others => '0');
        \$v6515%now\ <= (others => '0');
        \$13507%now\ <= (others => '0');
        \$19235%now\ <= (others => '0');
        \$17593%now\ <= (others => '0');
        \$17460_aux664_result%now\ <= (others => '0');
        \$v7283%now\ <= (others => '0');
        \$16986_compare6445898_result%now\ <= (others => '0');
        \$14930_r%now\ <= (others => '0');
        \$v6898%now\ <= (others => '0');
        \$v6003%now\ <= (others => '0');
        \$17466%now\ <= (others => '0');
        \$v6579%now\ <= (others => '0');
        \$v6121%now\ <= (others => '0');
        \$14621_modulo6685888_result%now\ <= (others => '0');
        \$13689%now\ <= (others => '0');
        \$14804_binop_int6435903_result%now\ <= (others => '0');
        \$12782%now\ <= (others => '0');
        \$18995%now\ <= (others => '0');
        \$v6110%now\ <= (others => '0');
        \$v6179%now\ <= (others => '0');
        \$18043%now\ <= (others => '0');
        \$19251_w%now\ <= (others => '0');
        \$14381%now\ <= (others => '0');
        \$v6066%now\ <= (others => '0');
        \$12546_dur%now\ <= (others => '0');
        \$v6911%now\ <= (others => '0');
        \$v6207%now\ <= (others => '0');
        \$15253_modulo6685896_result%now\ <= (others => '0');
        \$17889%now\ <= (others => '0');
        \$14311%now\ <= (others => '0');
        \$v6971%now\ <= (others => '0');
        \$v5999%now\ <= (others => '0');
        \$12906%now\ <= (others => '0');
        \$v7206%now\ <= (others => '0');
        \$14917_modulo6685888_id%now\ <= (others => '0');
        \$18661%now\ <= (others => '0');
        \$17957_hd%now\ <= (others => '0');
        \$12924_w%now\ <= (others => '0');
        \$v6546%now\ <= (others => '0');
        \$18280%now\ <= (others => '0');
        \$13148%now\ <= (others => '0');
        \$v6232%now\ <= (others => '0');
        \$18633_loop665_arg%now\ <= (others => '0');
        \$14757_modulo6685888_result%now\ <= (others => '0');
        \$13922_wait662_result%now\ <= (others => '0');
        \$v7364%now\ <= (others => '0');
        \$15580_modulo6685896_result%now\ <= (others => '0');
        \$15421_modulo6685888_id%now\ <= (others => '0');
        \$14610_r%now\ <= (others => '0');
        \$16916_compare6445898_id%now\ <= (others => '0');
        \$12886%now\ <= (others => '0');
        \$16195_forever6705924_id%now\ <= (others => '0');
        \$v6670%now\ <= (others => '0');
        \$13817%now\ <= (others => '0');
        \$v6817%now\ <= (others => '0');
        \$14221%now\ <= (others => '0');
        \$v6062%now\ <= (others => '0');
        \$17389%now\ <= (others => '0');
        \$v6563%now\ <= (others => '0');
        \$v6080%now\ <= (others => '0');
        \$v6799%now\ <= (others => '0');
        \$v7092%now\ <= (others => '0');
        \$14296%now\ <= (others => '0');
        \$17815%now\ <= (others => '0');
        \$v6463%now\ <= (others => '0');
        \$13100%now\ <= (others => '0');
        \$v6097%now\ <= (others => '0');
        \$v7203%now\ <= (others => '0');
        \$13808_hd%now\ <= (others => '0');
        \$13822%now\ <= (others => '0');
        \$16121_v%now\ <= (others => '0');
        \$v6403%now\ <= (others => '0');
        \$17000_sp%now\ <= (others => '0');
        \$12735%now\ <= (others => '0');
        \$v6424%now\ <= (others => '0');
        \$15261_modulo6685888_result%now\ <= (others => '0');
        \$17500%now\ <= (others => '0');
        \$17805%now\ <= (others => '0');
        \$v6421%now\ <= (others => '0');
        \$13510%now\ <= (others => '0');
        \$13940%now\ <= (others => '0');
        \$v7433%now\ <= (others => '0');
        \$15309_modulo6685895_arg%now\ <= (others => '0');
        \$18657%now\ <= (others => '0');
        \$16574_compare6445898_arg%now\ <= (others => '0');
        \$13317%now\ <= (others => '0');
        \$v6287%now\ <= (others => '0');
        \$12903%now\ <= (others => '0');
        \$16382%now\ <= (others => '0');
        \$15897%now\ <= (others => '0');
        \$14941_modulo6685888_result%now\ <= (others => '0');
        \$14909_modulo6685895_result%now\ <= (others => '0');
        \$v7135%now\ <= (others => '0');
        \$18806%now\ <= (others => '0');
        \$17458_loop666_arg%now\ <= (others => '0');
        \$12938%now\ <= (others => '0');
        \$15531_binop_int6435913_id%now\ <= (others => '0');
        \$15284_binop_int6435909_id%now\ <= (others => '0');
        \$13700%now\ <= (others => '0');
        \$18843%now\ <= (others => '0');
        \$15364_binop_int6435910_id%now\ <= (others => '0');
        \$12523_make_block579_arg%now\ <= (others => '0');
        \$v7245%now\ <= (others => '0');
        \$16317%now\ <= (others => '0');
        \$18348%now\ <= (others => '0');
        \$13101%now\ <= (others => '0');
        \$v6069%now\ <= (others => '0');
        \$16063_w6515922_result%now\ <= (others => '0');
        \$v6096%now\ <= (others => '0');
        \$12864_copy_root_in_ram6635886_arg%now\ <= (others => '0');
        \$14669_modulo6685895_arg%now\ <= (others => '0');
        \$17561%now\ <= (others => '0');
        \$19118%now\ <= (others => '0');
        \$14837_modulo6685888_id%now\ <= (others => '0');
        \$12694%now\ <= (others => '0');
        \$15284_binop_int6435909_arg%now\ <= (others => '0');
        \$12701%now\ <= (others => '0');
        \$v7450%now\ <= (others => '0');
        \$16158_forever6705923_id%now\ <= (others => '0');
        \$15101_modulo6685888_id%now\ <= (others => '0');
        \$v7145%now\ <= (others => '0');
        \$v6654%now\ <= (others => '0');
        \$v6042%now\ <= (others => '0');
        \$13234%now\ <= (others => '0');
        \$v6717%now\ <= (others => '0');
        \$15580_modulo6685896_arg%now\ <= (others => '0');
        \$15500_modulo6685896_result%now\ <= (others => '0');
        \$15447_forever6705911_arg%now\ <= (others => '0');
        \$18189%now\ <= (others => '0');
        \rdy6469%now\ <= (others => '0');
        \$17964%now\ <= (others => '0');
        \$18319%now\ <= (others => '0');
        \$v6920%now\ <= (others => '0');
        \$v6989%now\ <= (others => '0');
        \$14315_v%now\ <= (others => '0');
        \$18124%now\ <= (others => '0');
        \$16321%now\ <= (others => '0');
        \$v5986%now\ <= (others => '0');
        \$13384%now\ <= (others => '0');
        \$13379_hd%now\ <= (others => '0');
        \$15421_modulo6685888_arg%now\ <= (others => '0');
        \$v7365%now\ <= (others => '0');
        \$13922_wait662_id%now\ <= (others => '0');
        \$12549%now\ <= (others => '0');
        \$v6832%now\ <= (others => '0');
        \$v6765%now\ <= (others => '0');
        \$v6104%now\ <= (others => '0');
        \$18730%now\ <= (others => '0');
        \$18184%now\ <= (others => '0');
        \$17892%now\ <= (others => '0');
        \$v6543%now\ <= (others => '0');
        \$v6585%now\ <= (others => '0');
        \$17671%now\ <= (others => '0');
        \$v6106%now\ <= (others => '0');
        \$12704%now\ <= (others => '0');
        \$v7399%now\ <= (others => '0');
        \$v7110%now\ <= (others => '0');
        \$18118%now\ <= (others => '0');
        \$13540%now\ <= (others => '0');
        \$v6862%now\ <= (others => '0');
        \$15508_modulo6685888_result%now\ <= (others => '0');
        \$v7100%now\ <= (others => '0');
        \$17513_forever6705889_arg%now\ <= (others => '0');
        \$v6835%now\ <= (others => '0');
        \$16203%now\ <= (others => '0');
        \$15229_modulo6685895_result%now\ <= (others => '0');
        \$15910%now\ <= (others => '0');
        \$17456_loop665_result%now\ <= (others => '0');
        \$v5995%now\ <= (others => '0');
        \$13765%now\ <= (others => '0');
        \$12807_loop665_result%now\ <= (others => '0');
        \$v6373%now\ <= (others => '0');
        \$v6171%now\ <= (others => '0');
        \$18473%now\ <= (others => '0');
        \$v6758%now\ <= (others => '0');
        \$v7332%now\ <= (others => '0');
        \$v6646%now\ <= (others => '0');
        \$v6692%now\ <= (others => '0');
        \$v7188%now\ <= (others => '0');
        \$16063_w6515922_id%now\ <= (others => '0');
        \$v6562%now\ <= (others => '0');
        \$v6743%now\ <= (others => '0');
        \$v7426%now\ <= (others => '0');
        \$13463%now\ <= (others => '0');
        \$18686_copy_root_in_ram6635880_id%now\ <= (others => '0');
        \$v7378%now\ <= (others => '0');
        \$v6742%now\ <= (others => '0');
        \$14989_modulo6685895_result%now\ <= (others => '0');
        \$v7375%now\ <= (others => '0');
        \$15204_binop_int6435908_arg%now\ <= (others => '0');
        \$18845%now\ <= (others => '0');
        \$14008%now\ <= (others => '0');
        \$v6328%now\ <= (others => '0');
        \$v7355%now\ <= (others => '0');
        \$v7044%now\ <= (others => '0');
        \$v6319%now\ <= (others => '0');
        \$15364_binop_int6435910_arg%now\ <= (others => '0');
        \$v6965%now\ <= (others => '0');
        \$12879%now\ <= (others => '0');
        \$15284_binop_int6435909_result%now\ <= (others => '0');
        \$12804_loop665_result%now\ <= (others => '0');
        \$18546%now\ <= (others => '0');
        \$v7020%now\ <= (others => '0');
        \$15564_modulo6685888_result%now\ <= (others => '0');
        \$v7081%now\ <= (others => '0');
        \$v5872%now\ <= (others => '0');
        \$v7393%now\ <= (others => '0');
        \$14152%now\ <= (others => '0');
        \$v6766%now\ <= (others => '0');
        \$18841%now\ <= (others => '0');
        \$15661_binop_compare6455917_result%now\ <= (others => '0');
        \$13316%now\ <= (others => '0');
        \$13009_hd%now\ <= (others => '0');
        \$14909_modulo6685895_arg%now\ <= (others => '0');
        \$12682_make_block579_result%now\ <= (others => '0');
        \$18738%now\ <= (others => '0');
        \$16509%now\ <= (others => '0');
        \$12688%now\ <= (others => '0');
        \$15577_r%now\ <= (others => '0');
        \$v6093%now\ <= (others => '0');
        \$v6109%now\ <= (others => '0');
        \$15564_modulo6685888_arg%now\ <= (others => '0');
        \$16928_compbranch6505934_id%now\ <= (others => '0');
        \$14884_binop_int6435904_arg%now\ <= (others => '0');
        \$v6553%now\ <= (others => '0');
        \$14092%now\ <= (others => '0');
        \$v6535%now\ <= (others => '0');
        \$18732%now\ <= (others => '0');
        \$17066%now\ <= (others => '0');
        \$15389_modulo6685895_id%now\ <= (others => '0');
        \$v6660%now\ <= (others => '0');
        \$17337%now\ <= (others => '0');
        \$18826_w%now\ <= (others => '0');
        \$v6036%now\ <= (others => '0');
        \$17374_v%now\ <= (others => '0');
        \$17502%now\ <= (others => '0');
        \$12942%now\ <= (others => '0');
        \$14773_modulo6685896_id%now\ <= (others => '0');
        \$14757_modulo6685888_id%now\ <= (others => '0');
        \$18041%now\ <= (others => '0');
        \$v6547%now\ <= (others => '0');
        \$v6184%now\ <= (others => '0');
        \$12864_copy_root_in_ram6635886_id%now\ <= (others => '0');
        \$18470%now\ <= (others => '0');
        \$12835%now\ <= (others => '0');
        \$15909%now\ <= (others => '0');
        \$v6902%now\ <= (others => '0');
        \$17009_sp%now\ <= (others => '0');
        \$18476%now\ <= (others => '0');
        \$16626%now\ <= (others => '0');
        \$17804%now\ <= (others => '0');
        \$18443%now\ <= (others => '0');
        \$14701_modulo6685888_result%now\ <= (others => '0');
        \$v7167%now\ <= (others => '0');
        \$14902_res%now\ <= (others => '0');
        \$12717%now\ <= (others => '0');
        \$v6908%now\ <= (others => '0');
        \$13917%now\ <= (others => '0');
        \$16749_sp%now\ <= (others => '0');
        \$v6155%now\ <= (others => '0');
        \$17243%now\ <= (others => '0');
        \$v6442%now\ <= (others => '0');
        \$13923_make_block579_result%now\ <= (others => '0');
        \$v7445%now\ <= (others => '0');
        \$v6354%now\ <= (others => '0');
        \$14508_v%now\ <= (others => '0');
        \$15157_modulo6685888_arg%now\ <= (others => '0');
        \$19267%now\ <= (others => '0');
        \$16846_compare6445898_id%now\ <= (others => '0');
        \$15170_r%now\ <= (others => '0');
        \$v6616%now\ <= (others => '0');
        \$13926_make_block_n646_id%now\ <= (others => '0');
        \$18478%now\ <= (others => '0');
        \$16440%now\ <= (others => '0');
        \$15451_binop_int6435912_arg%now\ <= (others => '0');
        \$15980_v%now\ <= (others => '0');
        \$v6623%now\ <= (others => '0');
        \$14909_modulo6685895_id%now\ <= (others => '0');
        \$12830%now\ <= (others => '0');
        \$13149%now\ <= (others => '0');
        \$17164%now\ <= (others => '0');
        \$14463_v%now\ <= (others => '0');
        \$13019%now\ <= (others => '0');
        \$15613%now\ <= (others => '0');
        \$17535%now\ <= (others => '0');
        \$13818%now\ <= (others => '0');
        \$v6521%now\ <= (others => '0');
        \$16763_v%now\ <= (others => '0');
        \$18669%now\ <= (others => '0');
        \$18660%now\ <= (others => '0');
        \$v6137%now\ <= (others => '0');
        \$v6790%now\ <= (others => '0');
        \$v7117%now\ <= (others => '0');
        \$v6223%now\ <= (others => '0');
        \$13105_copy_root_in_ram6635884_arg%now\ <= (others => '0');
        \$v7387%now\ <= (others => '0');
        \$17547_copy_root_in_ram6635891_id%now\ <= (others => '0');
        \$15157_modulo6685888_id%now\ <= (others => '0');
        \$18632_loop666_arg%now\ <= (others => '0');
        \$17173%now\ <= (others => '0');
        \$15447_forever6705911_id%now\ <= (others => '0');
        \$15861_v%now\ <= (others => '0');
        \$13223_hd%now\ <= (others => '0');
        \$13524_hd%now\ <= (others => '0');
        \$16336%now\ <= (others => '0');
        \$v6899%now\ <= (others => '0');
        \$v7156%now\ <= (others => '0');
        \$15302_res%now\ <= (others => '0');
        \$19268%now\ <= (others => '0');
        \$18572%now\ <= (others => '0');
        \$v7459%now\ <= (others => '0');
        \$v7229%now\ <= (others => '0');
        \$17883%now\ <= (others => '0');
        \$18048%now\ <= (others => '0');
        \$13385%now\ <= (others => '0');
        \$17239_v%now\ <= (others => '0');
        \$14773_modulo6685896_result%now\ <= (others => '0');
        \$17592%now\ <= (others => '0');
        \$13926_make_block_n646_result%now\ <= (others => '0');
        \$17749%now\ <= (others => '0');
        \$18668%now\ <= (others => '0');
        \$v7093%now\ <= (others => '0');
        \$v6176%now\ <= (others => '0');
        \$12710%now\ <= (others => '0');
        \$18913%now\ <= (others => '0');
        \$v7107%now\ <= (others => '0');
        \$v6075%now\ <= (others => '0');
        \$v6031%now\ <= (others => '0');
        \$14861_modulo6685888_arg%now\ <= (others => '0');
        \$v6352%now\ <= (others => '0');
        \$13924_apply638_result%now\ <= (others => '0');
        \$15883%now\ <= (others => '0');
        \$v6684%now\ <= (others => '0');
        \$13309%now\ <= (others => '0');
        \$12829%now\ <= (others => '0');
        \$14273%now\ <= (others => '0');
        \rdy6504%now\ <= (others => '0');
        \$v6938%now\ <= (others => '0');
        \$17371_v%now\ <= (others => '0');
        \$v6880%now\ <= (others => '0');
        \$v7011%now\ <= (others => '0');
        \$17232%now\ <= (others => '0');
        \$12864_copy_root_in_ram6635886_result%now\ <= (others => '0');
        \$v6829%now\ <= (others => '0');
        \$v7056%now\ <= (others => '0');
        \$14139%now\ <= (others => '0');
        \$v6379%now\ <= (others => '0');
        \$17332_sp%now\ <= (others => '0');
        \$17048_w16565937_result%now\ <= (others => '0');
        \$19266%now\ <= (others => '0');
        \$15588_modulo6685888_result%now\ <= (others => '0');
        \$v7260%now\ <= (others => '0');
        \$14621_modulo6685888_arg%now\ <= (others => '0');
        \$13924_apply638_arg%now\ <= (others => '0');
        \$v6643%now\ <= (others => '0');
        \$v6152%now\ <= (others => '0');
        \$18994%now\ <= (others => '0');
        \$15250_r%now\ <= (others => '0');
        \$15044_binop_int6435906_result%now\ <= (others => '0');
        \$16650_sp%now\ <= (others => '0');
        \$v7350%now\ <= (others => '0');
        \$18633_loop665_result%now\ <= (others => '0');
        \$12553%now\ <= (others => '0');
        \$18044%now\ <= (others => '0');
        \$12720%now\ <= (others => '0');
        \$17594%now\ <= (others => '0');
        \$v6190%now\ <= (others => '0');
        \$v5964%now\ <= (others => '0');
        \$13926_make_block_n646_arg%now\ <= (others => '0');
        \$15077_modulo6685888_id%now\ <= (others => '0');
        \$v7021%now\ <= (others => '0');
        \$17018_w36575938_result%now\ <= (others => '0');
        \$v6180%now\ <= (others => '0');
        \$v6889%now\ <= (others => '0');
        \$15715_res%now\ <= (others => '0');
        \$16349_v%now\ <= (others => '0');
        \$14964_binop_int6435905_arg%now\ <= (others => '0');
        \$18998%now\ <= (others => '0');
        \$13158%now\ <= (others => '0');
        \$v6283%now\ <= (others => '0');
        \$17393%now\ <= (others => '0');
        \$v5948%now\ <= (others => '0');
        \$13092%now\ <= (others => '0');
        \$v6714%now\ <= (others => '0');
        \$v6325%now\ <= (others => '0');
        \$14997_modulo6685888_result%now\ <= (others => '0');
        \$v6550%now\ <= (others => '0');
        \$v6236%now\ <= (others => '0');
        \$12934%now\ <= (others => '0');
        \$v6588%now\ <= (others => '0');
        \$v6256%now\ <= (others => '0');
        \$17458_loop666_id%now\ <= (others => '0');
        \$17032%now\ <= (others => '0');
        \$12706%now\ <= (others => '0');
        \$16673_v%now\ <= (others => '0');
        \$13688%now\ <= (others => '0');
        \$v7427%now\ <= (others => '0');
        \$17458_loop666_result%now\ <= (others => '0');
        \$12681_wait662_arg%now\ <= (others => '0');
        \$18673%now\ <= (others => '0');
        \$17324%now\ <= (others => '0');
        \$14070_v%now\ <= (others => '0');
        \$12737%now\ <= (others => '0');
        \$19214%now\ <= (others => '0');
        \$15787_res%now\ <= (others => '0');
        \$14589_modulo6685895_arg%now\ <= (others => '0');
        \$v5967%now\ <= (others => '0');
        \$17968%now\ <= (others => '0');
        \$14738_v%now\ <= (others => '0');
        \$v5998%now\ <= (others => '0');
        \$18639%now\ <= (others => '0');
        \$13766%now\ <= (others => '0');
        \$15413_modulo6685896_arg%now\ <= (others => '0');
        \$15860%now\ <= (others => '0');
        \$v7010%now\ <= (others => '0');
        \$18564%now\ <= (others => '0');
        \$v7449%now\ <= (others => '0');
        \$v7046%now\ <= (others => '0');
        \$17532%now\ <= (others => '0');
        \$v6243%now\ <= (others => '0');
        \$19213%now\ <= (others => '0');
        \$13529%now\ <= (others => '0');
        \$v6493%now\ <= (others => '0');
        \$15421_modulo6685888_result%now\ <= (others => '0');
        \$18191%now\ <= (others => '0');
        \$14564_binop_int6435900_id%now\ <= (others => '0');
        \$12679_loop666_arg%now\ <= (others => '0');
        \$14406_v%now\ <= (others => '0');
        \$15619%now\ <= (others => '0');
        \$v6917%now\ <= (others => '0');
        \$16507%now\ <= (others => '0');
        \$v7116%now\ <= (others => '0');
        \$v7273%now\ <= (others => '0');
        \$14165%now\ <= (others => '0');
        \$13920_loop666_id%now\ <= (others => '0');
        \$15618%now\ <= (others => '0');
        \$16403%now\ <= (others => '0');
        \$17476%now\ <= (others => '0');
        \$13626%now\ <= (others => '0');
        \$17967%now\ <= (others => '0');
        \$12709%now\ <= (others => '0');
        \$v7213%now\ <= (others => '0');
        \$14861_modulo6685888_id%now\ <= (others => '0');
        \$v6844%now\ <= (others => '0');
        \$12804_loop665_arg%now\ <= (others => '0');
        \$14281%now\ <= (others => '0');
        \$16272%now\ <= (others => '0');
        \$17572%now\ <= (others => '0');
        \$12705%now\ <= (others => '0');
        \$12696%now\ <= (others => '0');
        \$13117%now\ <= (others => '0');
        \$13605%now\ <= (others => '0');
        \$16288%now\ <= (others => '0');
        \$12853_forever6705887_id%now\ <= (others => '0');
        \$17734_copy_root_in_ram6635892_result%now\ <= (others => '0');
        \$17759%now\ <= (others => '0');
        \$v6247%now\ <= (others => '0');
        \$16986_compare6445898_id%now\ <= (others => '0');
        \$17314%now\ <= (others => '0');
        \$v7197%now\ <= (others => '0');
        \$12680_loop665_arg%now\ <= (others => '0');
        \$18119%now\ <= (others => '0');
        \$v6072%now\ <= (others => '0');
        \$12760%now\ <= (others => '0');
        \$12548_dis%now\ <= (others => '0');
        \$15077_modulo6685888_arg%now\ <= (others => '0');
        \$14853_modulo6685896_result%now\ <= (others => '0');
        \$18737%now\ <= (others => '0');
        \$18918%now\ <= (others => '0');
        \$17237_sp%now\ <= (others => '0');
        \$15173_modulo6685896_arg%now\ <= (others => '0');
        \$17595%now\ <= (others => '0');
        \$17008%now\ <= (others => '0');
        \$17761_copy_root_in_ram6635891_arg%now\ <= (others => '0');
        \$v7101%now\ <= (others => '0');
        \$12847%now\ <= (others => '0');
        \$v6859%now\ <= (others => '0');
        \$12889%now\ <= (others => '0');
        \$18051%now\ <= (others => '0');
        \$v6219%now\ <= (others => '0');
        \$14826_r%now\ <= (others => '0');
        \$14033%now\ <= (others => '0');
        \$v6606%now\ <= (others => '0');
        \$18326%now\ <= (others => '0');
        \$18921%now\ <= (others => '0');
        \$13691%now\ <= (others => '0');
        \$v7083%now\ <= (others => '0');
        \$v6956%now\ <= (others => '0');
        \$15679_res%now\ <= (others => '0');
        \$v6666%now\ <= (others => '0');
        \$19239%now\ <= (others => '0');
        \$14024%now\ <= (others => '0');
        \$v7442%now\ <= (others => '0');
        \$16811_compare6445898_result%now\ <= (others => '0');
        \$14781_modulo6685888_arg%now\ <= (others => '0');
        \$v6335%now\ <= (others => '0');
        \$19260%now\ <= (others => '0');
        \$17347%now\ <= (others => '0');
        \$15333_modulo6685896_id%now\ <= (others => '0');
        \$18196%now\ <= (others => '0');
        \$v6752%now\ <= (others => '0');
        \$16300%now\ <= (others => '0');
        \$17673%now\ <= (others => '0');
        \$13227%now\ <= (others => '0');
        \$16612_compare6445898_arg%now\ <= (others => '0');
        \$13925_offsetclosure_n639_result%now\ <= (others => '0');
        \$v6409%now\ <= (others => '0');
        \$17814%now\ <= (others => '0');
        \$17585_hd%now\ <= (others => '0');
        \$17509_forever6705890_id%now\ <= (others => '0');
        \$17566%now\ <= (others => '0');
        \$12814%now\ <= (others => '0');
        \$19242%now\ <= (others => '0');
        \$17497%now\ <= (others => '0');
        \$13695%now\ <= (others => '0');
        \$v6394%now\ <= (others => '0');
        \$v7397%now\ <= (others => '0');
        \$v7289%now\ <= (others => '0');
        \$v7194%now\ <= (others => '0');
        \$17874_w%now\ <= (others => '0');
        \$18844%now\ <= (others => '0');
        \$15181_modulo6685888_arg%now\ <= (others => '0');
        \$18175_w%now\ <= (others => '0');
        \$v5876%now\ <= (others => '0');
        \$18676%now\ <= (others => '0');
        \$17539%now\ <= (others => '0');
        \$v7115%now\ <= (others => '0');
        \$v6263%now\ <= (others => '0');
        \$v6353%now\ <= (others => '0');
        \$18335_w%now\ <= (others => '0');
        \$18993%now\ <= (others => '0');
        \$13928_w652_id%now\ <= (others => '0');
        \$17504%now\ <= (others => '0');
        \$18046%now\ <= (others => '0');
        \$12670%now\ <= (others => '0');
        \$v5972%now\ <= (others => '0');
        \$v6133%now\ <= (others => '0');
        \$12743%now\ <= (others => '0');
        \$13539%now\ <= (others => '0');
        \$v5947%now\ <= (others => '0');
        \$17117_v%now\ <= (others => '0');
        \$15173_modulo6685896_result%now\ <= (others => '0');
        \$15819_v%now\ <= (others => '0');
        \$17547_copy_root_in_ram6635891_arg%now\ <= (others => '0');
        \$12681_wait662_id%now\ <= (others => '0');
        \$14043_v%now\ <= (others => '0');
        \$13814%now\ <= (others => '0');
        \$12803_loop666_arg%now\ <= (others => '0');
        \$v6436%now\ <= (others => '0');
        \$19136%now\ <= (others => '0');
        \$18674%now\ <= (others => '0');
        \$v6784%now\ <= (others => '0');
        \$v7296%now\ <= (others => '0');
        \$17395%now\ <= (others => '0');
        \$13236%now\ <= (others => '0');
        \$13464%now\ <= (others => '0');
        \$14051%now\ <= (others => '0');
        \$v7014%now\ <= (others => '0');
        \$17320%now\ <= (others => '0');
        \$v7095%now\ <= (others => '0');
        \$v6433%now\ <= (others => '0');
        \$12681_wait662_result%now\ <= (others => '0');
        \$13383%now\ <= (others => '0');
        \$14578_v%now\ <= (others => '0');
        \$v7112%now\ <= (others => '0');
        \$17675%now\ <= (others => '0');
        \$19127_w%now\ <= (others => '0');
        \$18808%now\ <= (others => '0');
        \$14148%now\ <= (others => '0');
        \$18705%now\ <= (others => '0');
        \$14804_binop_int6435903_id%now\ <= (others => '0');
        \$v6650%now\ <= (others => '0');
        \$v7267%now\ <= (others => '0');
        \$13624%now\ <= (others => '0');
        \$15588_modulo6685888_arg%now\ <= (others => '0');
        \$v7051%now\ <= (others => '0');
        \$v5867%now\ <= (others => '0');
        \$17388%now\ <= (others => '0');
        \$15173_modulo6685896_id%now\ <= (others => '0');
        \$16589_compbranch6505927_result%now\ <= (others => '0');
        \$14069%now\ <= (others => '0');
        \$v6531%now\ <= (others => '0');
        \$12713%now\ <= (others => '0');
        \$13021%now\ <= (others => '0');
        \$18666_next%now\ <= (others => '0');
        \$14446_v%now\ <= (others => '0');
        \$17677%now\ <= (others => '0');
        \$18740%now\ <= (others => '0');
        \$18842%now\ <= (others => '0');
        \$17972%now\ <= (others => '0');
        \$14989_modulo6685895_id%now\ <= (others => '0');
        \$17598%now\ <= (others => '0');
        \$12522_wait662_id%now\ <= (others => '0');
        \$18701%now\ <= (others => '0');
        \$16662_fill6535928_arg%now\ <= (others => '0');
        \$17490_next%now\ <= (others => '0');
        \$v6759%now\ <= (others => '0');
        \$16928_compbranch6505934_arg%now\ <= (others => '0');
        \$18922%now\ <= (others => '0');
        \$18464_hd%now\ <= (others => '0');
        \$16963_compbranch6505935_result%now\ <= (others => '0');
        \$13992_v%now\ <= (others => '0');
        \$15508_modulo6685888_arg%now\ <= (others => '0');
        \$12929_hd%now\ <= (others => '0');
        \$v7457%now\ <= (others => '0');
        \$13538%now\ <= (others => '0');
        \$16457%now\ <= (others => '0');
        \$15306_r%now\ <= (others => '0');
        \$v6705%now\ <= (others => '0');
        \$18122%now\ <= (others => '0');
        \$v7102%now\ <= (others => '0');
        \$19143%now\ <= (others => '0');
        \$18670_next%now\ <= (others => '0');
        \$18634_aux664_arg%now\ <= (others => '0');
        \$18793_copy_root_in_ram6635879_id%now\ <= (others => '0');
        \$15149_modulo6685895_id%now\ <= (others => '0');
        \$16788_compbranch6505930_result%now\ <= (others => '0');
        \$13535%now\ <= (others => '0');
        \$15545_v%now\ <= (others => '0');
        \$17482%now\ <= (others => '0');
        \$v7061%now\ <= (others => '0');
        \$v6253%now\ <= (others => '0');
        \$13897%now\ <= (others => '0');
        \$18735%now\ <= (others => '0');
        \$v7126%now\ <= (others => '0');
        \$18281%now\ <= (others => '0');
        \$16473%now\ <= (others => '0');
        \$14917_modulo6685888_result%now\ <= (others => '0');
        \$16741%now\ <= (others => '0');
        \$16510_forever6705925_arg%now\ <= (others => '0');
        \$v6536%now\ <= (others => '0');
        \$12811%now\ <= (others => '0');
        \$v6796%now\ <= (others => '0');
        \$18459_w%now\ <= (others => '0');
        \$14413_v%now\ <= (others => '0');
        \$12520_loop666_result%now\ <= (others => '0');
        \$16612_compare6445898_id%now\ <= (others => '0');
        \$17747%now\ <= (others => '0');
        \$v7104%now\ <= (others => '0');
        \$13939%now\ <= (others => '0');
        \$15661_binop_compare6455917_id%now\ <= (others => '0');
        \$17973%now\ <= (others => '0');
        \$12804_loop665_id%now\ <= (others => '0');
        \$17758%now\ <= (others => '0');
        \$12719%now\ <= (others => '0');
        \$15397_modulo6685888_id%now\ <= (others => '0');
        \$17105_w06555936_arg%now\ <= (others => '0');
        \$12792%now\ <= (others => '0');
        \$16194%now\ <= (others => '0');
        \$v7176%now\ <= (others => '0');
        \$14829_modulo6685895_arg%now\ <= (others => '0');
        \$18049%now\ <= (others => '0');
        \$13536%now\ <= (others => '0');
        \$12842%now\ <= (others => '0');
        \$v7182%now\ <= (others => '0');
        \$v6511%now\ <= (others => '0');
        \$14693_modulo6685896_id%now\ <= (others => '0');
        \$13023%now\ <= (others => '0');
        \$v6098%now\ <= (others => '0');
        \$15792_compare6445897_arg%now\ <= (others => '0');
        \$v6905%now\ <= (others => '0');
        \$13313%now\ <= (others => '0');
        \$14552%now\ <= (others => '0');
        \$16840_b%now\ <= (others => '0');
        \$16568_b%now\ <= (others => '0');
        \$14423_v%now\ <= (others => '0');
        \$v6527%now\ <= (others => '0');
        \$18262%now\ <= (others => '0');
        \$13078_copy_root_in_ram6635885_result%now\ <= (others => '0');
        \$18351%now\ <= (others => '0');
        \$16232%now\ <= (others => '0');
        \$16133%now\ <= (others => '0');
        \$15711_v%now\ <= (others => '0');
        \$15614_forever6705914_id%now\ <= (others => '0');
        \$13004_w%now\ <= (others => '0');
        \$12803_loop666_id%now\ <= (others => '0');
        \$12744%now\ <= (others => '0');
        \$13311%now\ <= (others => '0');
        \$18664_next%now\ <= (others => '0');
        \$19264%now\ <= (others => '0');
        \$13472_next%now\ <= (others => '0');
        \$16858_compbranch6505932_id%now\ <= (others => '0');
        \$v7096%now\ <= (others => '0');
        \$17966%now\ <= (others => '0');
        \$v6787%now\ <= (others => '0');
        \$17459_loop665_result%now\ <= (others => '0');
        \$v7120%now\ <= (others => '0');
        \$17310%now\ <= (others => '0');
        \$17492_next%now\ <= (others => '0');
        \$v6045%now\ <= (others => '0');
        \$17748%now\ <= (others => '0');
        \$18638%now\ <= (others => '0');
        \$15792_compare6445897_id%now\ <= (others => '0');
        \$13963%now\ <= (others => '0');
        \$v6140%now\ <= (others => '0');
        \$12933%now\ <= (others => '0');
        \$18640%now\ <= (others => '0');
        \$13528%now\ <= (others => '0');
        \$v7254%now\ <= (others => '0');
        \$16881_compare6445898_id%now\ <= (others => '0');
        \$17460_aux664_arg%now\ <= (others => '0');
        \$12523_make_block579_result%now\ <= (others => '0');
        \$13922_wait662_arg%now\ <= (others => '0');
        \$v6156%now\ <= (others => '0');
        \$v6814%now\ <= (others => '0');
        \$v7419%now\ <= (others => '0');
        \$15451_binop_int6435912_result%now\ <= (others => '0');
        \$v6322%now\ <= (others => '0');
        \$17331_sp%now\ <= (others => '0');
        \$17894%now\ <= (others => '0');
        \$v6002%now\ <= (others => '0');
        \$v6476%now\ <= (others => '0');
        \$13239%now\ <= (others => '0');
        \$12708%now\ <= (others => '0');
        \$18812%now\ <= (others => '0');
        \$v6187%now\ <= (others => '0');
        \$v7072%now\ <= (others => '0');
        \rdy6148%now\ <= (others => '0');
        \$18047%now\ <= (others => '0');
        \$14644_binop_int6435901_id%now\ <= (others => '0');
        \$14597_modulo6685888_id%now\ <= (others => '0');
        \$v7103%now\ <= (others => '0');
        \$19261%now\ <= (others => '0');
        \$16893_compbranch6505933_arg%now\ <= (others => '0');
        \$13390%now\ <= (others => '0');
        \$16534%now\ <= (others => '0');
        \$v7191%now\ <= (others => '0');
        \$19002%now\ <= (others => '0');
        \$v7041%now\ <= (others => '0');
        \$v6968%now\ <= (others => '0');
        \$v7127%now\ <= (others => '0');
        \$17520_copy_root_in_ram6635893_result%now\ <= (others => '0');
        \$v6332%now\ <= (others => '0');
        \$13229%now\ <= (others => '0');
        \$v6159%now\ <= (others => '0');
        \$15684_compare6445897_id%now\ <= (others => '0');
        \$v7114%now\ <= (others => '0');
        \$17544%now\ <= (others => '0');
        \$v6704%now\ <= (others => '0');
        \$18040%now\ <= (others => '0');
        \$17786%now\ <= (others => '0');
        \$v7233%now\ <= (others => '0');
        \$14207_loop_push6495899_arg%now\ <= (others => '0');
        \$16709%now\ <= (others => '0');
        \$v7113%now\ <= (others => '0');
        \$14724_binop_int6435902_arg%now\ <= (others => '0');
        \$13232%now\ <= (others => '0');
        \$16986_compare6445898_arg%now\ <= (others => '0');
        \$v6054%now\ <= (others => '0');
        \$16074_v%now\ <= (others => '0');
        \$v6781%now\ <= (others => '0');
        \$v7047%now\ <= (others => '0');
        \$17503%now\ <= (others => '0');
        \$13147%now\ <= (others => '0');
        \$v6259%now\ <= (others => '0');
        \$v6144%now\ <= (others => '0');
        \$13018%now\ <= (others => '0');
        \$v6603%now\ <= (others => '0');
        \$14016_v%now\ <= (others => '0');
        \$16752_fill6545929_id%now\ <= (others => '0');
        \$v5973%now\ <= (others => '0');
        \$13815%now\ <= (others => '0');
        \$v7033%now\ <= (others => '0');
        \$v5983%now\ <= (others => '0');
        \$19271%now\ <= (others => '0');
        \$v6735%now\ <= (others => '0');
        \$v6769%now\ <= (others => '0');
        \$v7242%now\ <= (others => '0');
        \$16508%now\ <= (others => '0');
        \$12808_aux664_arg%now\ <= (others => '0');
        \$18708%now\ <= (others => '0');
        \$18991%now\ <= (others => '0');
        \$14471%now\ <= (others => '0');
        \$v7070%now\ <= (others => '0');
        \$12547%now\ <= (others => '0');
        \$v7031%now\ <= (others => '0');
        \$v6315%now\ <= (others => '0');
        \$12674%now\ <= (others => '0');
        \$12846%now\ <= (others => '0');
        \$17010%now\ <= (others => '0');
        \$17560%now\ <= (others => '0');
        \$16156%now\ <= (others => '0');
        \$15021_modulo6685888_id%now\ <= (others => '0');
        \$13925_offsetclosure_n639_arg%now\ <= (others => '0');
        \$14898_v%now\ <= (others => '0');
        \$14693_modulo6685896_result%now\ <= (others => '0');
        \$15497_r%now\ <= (others => '0');
        \$13105_copy_root_in_ram6635884_id%now\ <= (others => '0');
        \$17434%now\ <= (others => '0');
        \$16515%now\ <= (others => '0');
        \$14512_v%now\ <= (others => '0');
        \$14300_v%now\ <= (others => '0');
        \$18261%now\ <= (others => '0');
        \$17207_arg%now\ <= (others => '0');
        \$13315%now\ <= (others => '0');
        \$18992%now\ <= (others => '0');
        \$18344%now\ <= (others => '0');
        \$17183%now\ <= (others => '0');
        \$v7032%now\ <= (others => '0');
        \result6112%now\ <= (others => '0');
        \$v5960%now\ <= (others => '0');
        \$v7084%now\ <= (others => '0');
        \$v6639%now\ <= (others => '0');
        \$v7060%now\ <= (others => '0');
        \$18030_w%now\ <= (others => '0');
        \$18190%now\ <= (others => '0');
        \$16380_v%now\ <= (others => '0');
        \$v6295%now\ <= (others => '0');
        \$18924%now\ <= (others => '0');
        \$12659%now\ <= (others => '0');
        \$v6111%now\ <= (others => '0');
        \$v6011%now\ <= (others => '0');
        \$12891_copy_root_in_ram6635884_result%now\ <= (others => '0');
        \$18621%now\ <= (others => '0');
        \$14185_next_env%now\ <= (others => '0');
        \$17166%now\ <= (others => '0');
        \$v6059%now\ <= (others => '0');
        \$12703%now\ <= (others => '0');
        \$v6358%now\ <= (others => '0');
        \$12832%now\ <= (others => '0');
        \$15684_compare6445897_result%now\ <= (others => '0');
        \$v7111%now\ <= (others => '0');
        \$17895%now\ <= (others => '0');
        \$13812%now\ <= (others => '0');
        \$18632_loop666_id%now\ <= (others => '0');
        \$17952_w%now\ <= (others => '0');
        \$13820%now\ <= (others => '0');
        \$13533%now\ <= (others => '0');
        \$15805_binop_compare6455921_result%now\ <= (others => '0');
        \$15413_modulo6685896_id%now\ <= (others => '0');
        \$13977_v%now\ <= (others => '0');
        \$v6294%now\ <= (others => '0');
        \$12857_forever6705883_id%now\ <= (others => '0');
        \$v7438%now\ <= (others => '0');
        \$v7082%now\ <= (others => '0');
        \$v6415%now\ <= (others => '0');
        \$v5982%now\ <= (others => '0');
        \$19265%now\ <= (others => '0');
        \$17011%now\ <= (others => '0');
        \$v7012%now\ <= (others => '0');
        \$17505_forever6705894_id%now\ <= (others => '0');
        \$v7282%now\ <= (others => '0');
        \$12813%now\ <= (others => '0');
        \$17499%now\ <= (others => '0');
        \$v6457%now\ <= (others => '0');
        \$13150%now\ <= (others => '0');
        \$17808%now\ <= (others => '0');
        \$v6820%now\ <= (others => '0');
        \$17970%now\ <= (others => '0');
        \$12803_loop666_result%now\ <= (others => '0');
        \$v7276%now\ <= (others => '0');
        \$14964_binop_int6435905_result%now\ <= (others => '0');
        \$v7134%now\ <= (others => '0');
        \$17809%now\ <= (others => '0');
        \$16404%now\ <= (others => '0');
        \$v7157%now\ <= (others => '0');
        \$17969%now\ <= (others => '0');
        \$v6280%now\ <= (others => '0');
        \$12845%now\ <= (others => '0');
        \$v6361%now\ <= (others => '0');
        \$12561%now\ <= (others => '0');
        \$17545%now\ <= (others => '0');
        \$18634_aux664_id%now\ <= (others => '0');
        \$15410_r%now\ <= (others => '0');
        \$v6582%now\ <= (others => '0');
        \$v6600%now\ <= (others => '0');
        \$15062_res%now\ <= (others => '0');
        \$v6264%now\ <= (others => '0');
        \$14342%now\ <= (others => '0');
        \$v6691%now\ <= (others => '0');
        \$12562%now\ <= (others => '0');
        \result5939%now\ <= (others => '0');
        \$12657%now\ <= (others => '0');
        \$v7130%now\ <= (others => '0');
        \$16193%now\ <= (others => '0');
        \$16916_compare6445898_result%now\ <= (others => '0');
        \$18839%now\ <= (others => '0');
        \$13787%now\ <= (others => '0');
        \$v7303%now\ <= (others => '0');
        \$19146%now\ <= (others => '0');
        \$15684_compare6445897_arg%now\ <= (others => '0');
        \$15142_res%now\ <= (others => '0');
        \$12905%now\ <= (others => '0');
        \$v6267%now\ <= (others => '0');
        \$18658%now\ <= (others => '0');
        \$13386%now\ <= (others => '0');
        \$17465%now\ <= (others => '0');
        \$v6477%now\ <= (others => '0');
        \$13025%now\ <= (others => '0');
        \$18678%now\ <= (others => '0');
        \$16461%now\ <= (others => '0');
        \$v6774%now\ <= (others => '0');
        \$18180_hd%now\ <= (others => '0');
        \$v6811%now\ <= (others => '0');
        \$13791%now\ <= (others => '0');
        \$14464_v%now\ <= (others => '0');
        \$15851_argument1%now\ <= (others => '0');
        \$13022%now\ <= (others => '0');
        \$15101_modulo6685888_arg%now\ <= (others => '0');
        \$13124%now\ <= (others => '0');
        \$v6762%now\ <= (others => '0');
        \$v6720%now\ <= (others => '0');
        \$v6528%now\ <= (others => '0');
        \$v6083%now\ <= (others => '0');
        \$16724%now\ <= (others => '0');
        \$v6524%now\ <= (others => '0');
        \$v6448%now\ <= (others => '0');
        \$17184%now\ <= (others => '0');
        \$13228%now\ <= (others => '0');
        \$19139%now\ <= (others => '0');
        \$v7036%now\ <= (others => '0');
        \$v6755%now\ <= (others => '0');
        \$17533%now\ <= (others => '0');
        \result5974%now\ <= (others => '0');
        \$v7037%now\ <= (others => '0');
        \$18589%now\ <= (others => '0');
        \$14669_modulo6685895_result%now\ <= (others => '0');
        \$13813%now\ <= (others => '0');
        \$17105_w06555936_result%now\ <= (others => '0');
        \$13921_loop665_arg%now\ <= (others => '0');
        \$17599%now\ <= (others => '0');
        \$13921_loop665_result%now\ <= (others => '0');
        \$v7401%now\ <= (others => '0');
        \$v6980%now\ <= (others => '0');
        \$16337%now\ <= (others => '0');
        \$17534%now\ <= (others => '0');
        \$12558%now\ <= (others => '0');
        \$v6926%now\ <= (others => '0');
        \$16811_compare6445898_id%now\ <= (others => '0');
        \$v5989%now\ <= (others => '0');
        \$14103%now\ <= (others => '0');
        \$15556_modulo6685895_arg%now\ <= (others => '0');
        \$19147%now\ <= (others => '0');
        \$16383%now\ <= (others => '0');
        \$v7149%now\ <= (others => '0');
        \$13314%now\ <= (others => '0');
        \$15639_v%now\ <= (others => '0');
        \$16624_argument2%now\ <= (others => '0');
        \$15069_modulo6685895_result%now\ <= (others => '0');
        \$16662_fill6535928_id%now\ <= (others => '0');
        \rdy6113%now\ <= (others => '0');
        \$17542%now\ <= (others => '0');
        \$v6345%now\ <= (others => '0');
        \$v6194%now\ <= (others => '0');
        \$v6571%now\ <= (others => '0');
        \$15531_binop_int6435913_result%now\ <= (others => '0');
        \$v6439%now\ <= (others => '0');
        \$v6079%now\ <= (others => '0');
        \$15621_forever6705915_arg%now\ <= (others => '0');
        \$17884%now\ <= (others => '0');
        \$v7097%now\ <= (others => '0');
        \$13927_branch_if648_id%now\ <= (others => '0');
        \$14982_res%now\ <= (others => '0');
        \$18353%now\ <= (others => '0');
        \$v7347%now\ <= (others => '0');
        \$16846_compare6445898_arg%now\ <= (others => '0');
        \$v6895%now\ <= (others => '0');
        \$16195_forever6705924_arg%now\ <= (others => '0');
        \$17589%now\ <= (others => '0');
        \$13017%now\ <= (others => '0');
        \$15747_v%now\ <= (others => '0');
        \$16662_fill6535928_result%now\ <= (others => '0');
        \$18345%now\ <= (others => '0');
        \$v7122%now\ <= (others => '0');
        \$17048_w16565937_id%now\ <= (others => '0');
        \$18686_copy_root_in_ram6635880_result%now\ <= (others => '0');
        \$15093_modulo6685896_id%now\ <= (others => '0');
        \$18736%now\ <= (others => '0');
        \$18671%now\ <= (others => '0');
        \$15500_modulo6685896_id%now\ <= (others => '0');
        \$v7226%now\ <= (others => '0');
        \$17459_loop665_id%now\ <= (others => '0');
        \$15333_modulo6685896_arg%now\ <= (others => '0');
        \$17807%now\ <= (others => '0');
        \$v6220%now\ <= (others => '0');
        \$13821%now\ <= (others => '0');
        \$18035_hd%now\ <= (others => '0');
        \$v6290%now\ <= (others => '0');
        \$17172%now\ <= (others => '0');
        \$13394%now\ <= (others => '0');
        \$19338%now\ <= (others => '0');
        \$17368_v%now\ <= (others => '0');
        \$v5871%now\ <= (others => '0');
        \$13958%now\ <= (others => '0');
        \$12824%now\ <= (others => '0');
        \$17562%now\ <= (others => '0');
        \$16322%now\ <= (others => '0');
        \$v7105%now\ <= (others => '0');
        \$13698%now\ <= (others => '0');
        \$17520_copy_root_in_ram6635893_arg%now\ <= (others => '0');
        \$15556_modulo6685895_id%now\ <= (others => '0');
        \$13105_copy_root_in_ram6635884_result%now\ <= (others => '0');
        \$12891_copy_root_in_ram6635884_id%now\ <= (others => '0');
        \$12806_loop666_arg%now\ <= (others => '0');
        \$v6566%now\ <= (others => '0');
        \$15181_modulo6685888_id%now\ <= (others => '0');
        \$v7080%now\ <= (others => '0');
        \$v6675%now\ <= (others => '0');
        \$v6576%now\ <= (others => '0');
        \$16998_argument3%now\ <= (others => '0');
        \$v7423%now\ <= (others => '0');
        \$18728%now\ <= (others => '0');
        \$16157%now\ <= (others => '0');
        \$13684_hd%now\ <= (others => '0');
        \$19111%now\ <= (others => '0');
        \$v6647%now\ <= (others => '0');
        \$13091%now\ <= (others => '0');
        \$13143_hd%now\ <= (others => '0');
        \$18793_copy_root_in_ram6635879_result%now\ <= (others => '0');
        \$15769_binop_compare6455920_result%now\ <= (others => '0');
        \$16462%now\ <= (others => '0');
        \$14265%now\ <= (others => '0');
        \$12916%now\ <= (others => '0');
        \$v6244%now\ <= (others => '0');
        \$12742%now\ <= (others => '0');
        \$13119%now\ <= (others => '0');
        \$13972_v%now\ <= (others => '0');
        \$14884_binop_int6435904_result%now\ <= (others => '0');
        \$13951%now\ <= (others => '0');
        \$v7024%now\ <= (others => '0');
        \$13923_make_block579_arg%now\ <= (others => '0');
        \$15648_compare6445897_result%now\ <= (others => '0');
        \$17330_sp%now\ <= (others => '0');
        \$v6620%now\ <= (others => '0');
        \$17353%now\ <= (others => '0');
        \$v6983%now\ <= (others => '0');
        \$v7257%now\ <= (others => '0');
        \$v6663%now\ <= (others => '0');
        \$13118%now\ <= (others => '0');
        \$v6032%now\ <= (others => '0');
        \$18672%now\ <= (others => '0');
        \$19074%now\ <= (others => '0');
        \$15309_modulo6685895_id%now\ <= (others => '0');
        \$v6260%now\ <= (others => '0');
        \$19076%now\ <= (others => '0');
        \rdy5975%now\ <= (others => '0');
        \$15124_binop_int6435907_result%now\ <= (others => '0');
        \$16334_v%now\ <= (others => '0');
        \$v7270%now\ <= (others => '0');
        \$18042%now\ <= (others => '0');
        \$18611%now\ <= (others => '0');
        \$14377_v%now\ <= (others => '0');
        \$16381_v%now\ <= (others => '0');
        \$v6076%now\ <= (others => '0');
        \$15908%now\ <= (others => '0');
        \$12563%now\ <= (others => '0');
        \$v7026%now\ <= (others => '0');
        \$v6698%now\ <= (others => '0');
        \$15013_modulo6685896_result%now\ <= (others => '0');
        \$12805_aux664_arg%now\ <= (others => '0');
        \$v7075%now\ <= (others => '0');
        \$13024%now\ <= (others => '0');
        \$13965%now\ <= (others => '0');
        \$18573%now\ <= (others => '0');
        \$v6124%now\ <= (others => '0');
        \$17481%now\ <= (others => '0');
        \$v6215%now\ <= (others => '0');
        \$15720_compare6445897_result%now\ <= (others => '0');
        \$v7160%now\ <= (others => '0');
        \$v6497%now\ <= (others => '0');
        \$15044_binop_int6435906_arg%now\ <= (others => '0');
        \$13097%now\ <= (others => '0');
        \$17456_loop665_arg%now\ <= (others => '0');
        \$13952%now\ <= (others => '0');
        \$15093_modulo6685896_result%now\ <= (others => '0');
        \$13924_apply638_id%now\ <= (others => '0');
        \$v6556%now\ <= (others => '0');
        \$14701_modulo6685888_id%now\ <= (others => '0');
        \$12687%now\ <= (others => '0');
        \$15473_r%now\ <= (others => '0');
        \$17061%now\ <= (others => '0');
        \$16725%now\ <= (others => '0');
        \$v6412%now\ <= (others => '0');
        \$v7407%now\ <= (others => '0');
        \$v6747%now\ <= (others => '0');
        \$12831%now\ <= (others => '0');
        \$16651%now\ <= (others => '0');
        \$14781_modulo6685888_id%now\ <= (others => '0');
        \$16658%now\ <= (others => '0');
        \$v7136%now\ <= (others => '0');
        \$14589_modulo6685895_id%now\ <= (others => '0');
        \$v5968%now\ <= (others => '0');
        \$v6339%now\ <= (others => '0');
        \$16788_compbranch6505930_id%now\ <= (others => '0');
        \$17486%now\ <= (others => '0');
        \$v6331%now\ <= (others => '0');
        \$18553%now\ <= (others => '0');
        \$14034_v%now\ <= (others => '0');
        \$v7410%now\ <= (others => '0');
        \$v7131%now\ <= (others => '0');
        \$18284%now\ <= (others => '0');
        \$v7390%now\ <= (others => '0');
        \$13306%now\ <= (others => '0');
        \$v6539%now\ <= (others => '0');
        \$v7341%now\ <= (others => '0');
        \$15090_r%now\ <= (others => '0');
        \$14906_r%now\ <= (others => '0');
        \$13462%now\ <= (others => '0');
        \$19270%now\ <= (others => '0');
        \$v6850%now\ <= (others => '0');
        \$v7430%now\ <= (others => '0');
        \$v6671%now\ <= (others => '0');
        \$15149_modulo6685895_result%now\ <= (others => '0');
        \$15756_compare6445897_id%now\ <= (others => '0');
        \$v6418%now\ <= (others => '0');
        \$v6250%now\ <= (others => '0');
        \$v6051%now\ <= (others => '0');
        \$15621_forever6705915_id%now\ <= (others => '0');
        \$v6886%now\ <= (others => '0');
        \$16858_compbranch6505932_result%now\ <= (others => '0');
        \$15222_res%now\ <= (others => '0');
        \$v6770%now\ <= (others => '0');
        \$v7040%now\ <= (others => '0');
        \$16301%now\ <= (others => '0');
        \$13911%now\ <= (others => '0');
        \$17680%now\ <= (others => '0');
        \$v6191%now\ <= (others => '0');
        \$15138_v%now\ <= (others => '0');
        \$v6486%now\ <= (others => '0');
        \$13152%now\ <= (others => '0');
        \$16155%now\ <= (others => '0');
        \$14933_modulo6685896_arg%now\ <= (others => '0');
        \$12693%now\ <= (others => '0');
        \$v7106%now\ <= (others => '0');
        \$v7067%now\ <= (others => '0');
        \$13920_loop666_result%now\ <= (others => '0');
        \$16293%now\ <= (others => '0');
        \$13159%now\ <= (others => '0');
        \$13953%now\ <= (others => '0');
        \$15625_binop_compare6455916_arg%now\ <= (others => '0');
        \$13015%now\ <= (others => '0');
        \$17799_hd%now\ <= (others => '0');
        \$v6039%now\ <= (others => '0');
        \$15611%now\ <= (others => '0');
        \$v6808%now\ <= (others => '0');
        \$17444%now\ <= (others => '0');
        \$14853_modulo6685896_id%now\ <= (others => '0');
        \$18665%now\ <= (others => '0');
        \$19132_hd%now\ <= (others => '0');
        \$16313_v%now\ <= (others => '0');
        \$14757_modulo6685888_arg%now\ <= (others => '0');
        \$18710%now\ <= (others => '0');
        \$v5979%now\ <= (others => '0');
        \$v6006%now\ <= (others => '0');
        \$14621_modulo6685888_id%now\ <= (others => '0');
        \$14941_modulo6685888_id%now\ <= (others => '0');
        \$19073%now\ <= (others => '0');
        \$15733_binop_compare6455919_id%now\ <= (others => '0');
        \$15620%now\ <= (others => '0');
        \$17596%now\ <= (others => '0');
        \$16413%now\ <= (others => '0');
        \$19141%now\ <= (others => '0');
        \$17753%now\ <= (others => '0');
        \$16706%now\ <= (others => '0');
        \$16296%now\ <= (others => '0');
        \$v7001%now\ <= (others => '0');
        \$18468%now\ <= (others => '0');
        \$19000%now\ <= (others => '0');
        \$v5877%now\ <= (others => '0');
        \$16951_compare6445898_id%now\ <= (others => '0');
        \$13231%now\ <= (others => '0');
        \$v6024%now\ <= (others => '0');
        \$13130%now\ <= (others => '0');
        \$15469_res%now\ <= (others => '0');
        \$18471%now\ <= (others => '0');
        \$v6793%now\ <= (others => '0');
        \$v7266%now\ <= (others => '0');
        \$18350%now\ <= (others => '0');
        \$16357%now\ <= (others => '0');
        \$15149_modulo6685895_arg%now\ <= (others => '0');
        \$13987_v%now\ <= (others => '0');
        \$v7055%now\ <= (others => '0');
        \$17483%now\ <= (others => '0');
        \$14260%now\ <= (others => '0');
        \$15588_modulo6685888_id%now\ <= (others => '0');
        \$v7309%now\ <= (others => '0');
        \$15643_res%now\ <= (others => '0');
        \$13078_copy_root_in_ram6635885_arg%now\ <= (others => '0');
        \$18914%now\ <= (others => '0');
        \$17660_w%now\ <= (others => '0');
        \$16846_compare6445898_result%now\ <= (others => '0');
        \$18817%now\ <= (others => '0');
        \$v6871%now\ <= (others => '0');
        \$17672%now\ <= (others => '0');
        \$19148%now\ <= (others => '0');
        \$v7329%now\ <= (others => '0');
        \$19072%now\ <= (others => '0');
        \$15733_binop_compare6455919_result%now\ <= (others => '0');
        \$14081%now\ <= (others => '0');
        \$18545%now\ <= (others => '0');
        \$13889%now\ <= (others => '0');
        \$14015%now\ <= (others => '0');
        \$12840_next%now\ <= (others => '0');
        \$18686_copy_root_in_ram6635880_arg%now\ <= (others => '0');
        \$14742_res%now\ <= (others => '0');
        \$14586_r%now\ <= (others => '0');
        \$18195%now\ <= (others => '0');
        \$v6540%now\ <= (others => '0');
        \$18793_copy_root_in_ram6635879_arg%now\ <= (others => '0');
        \$15317_modulo6685888_id%now\ <= (others => '0');
        \$16551_compbranch6505926_result%now\ <= (others => '0');
        \$17811%now\ <= (others => '0');
        \$16980_b%now\ <= (others => '0');
        \$18349%now\ <= (others => '0');
        \$15451_binop_int6435912_id%now\ <= (others => '0');
        \$14002_v%now\ <= (others => '0');
        \$14997_modulo6685888_arg%now\ <= (others => '0');
        \$16335_v%now\ <= (others => '0');
        \$13014%now\ <= (others => '0');
        \$v6977%now\ <= (others => '0');
        \$18039%now\ <= (others => '0');
        \$13448%now\ <= (others => '0');
        \$17571%now\ <= (others => '0');
        \$17757%now\ <= (others => '0');
        \$v6018%now\ <= (others => '0');
        \$16358%now\ <= (others => '0');
        \$v7052%now\ <= (others => '0');
        \$17352%now\ <= (others => '0');
        \$17756%now\ <= (others => '0');
        \$v6141%now\ <= (others => '0');
        \$13391%now\ <= (others => '0');
        \$v6086%now\ <= (others => '0');
        \$v6145%now\ <= (others => '0');
        \$15066_r%now\ <= (others => '0');
        \result6147%now\ <= (others => '0');
        \$15446%now\ <= (others => '0');
        \$v6877%now\ <= (others => '0');
        \$16041_v%now\ <= (others => '0');
        \$16063_w6515922_arg%now\ <= (others => '0');
        \$12700%now\ <= (others => '0');
        \$16951_compare6445898_result%now\ <= (others => '0');
        \$v6210%now\ <= (others => '0');
        \$15564_modulo6685888_id%now\ <= (others => '0');
        \$12721%now\ <= (others => '0');
        \$18920%now\ <= (others => '0');
        \$14393_hd%now\ <= (others => '0');
        \$18282%now\ <= (others => '0');
        \$v7141%now\ <= (others => '0');
        \$15157_modulo6685888_result%now\ <= (others => '0');
        \$14850_r%now\ <= (others => '0');
        \$17601%now\ <= (others => '0');
        \$v6310%now\ <= (others => '0');
        \$14493_v%now\ <= (others => '0');
        \$12711%now\ <= (others => '0');
        \$v5864%now\ <= (others => '0');
        \$v6483%now\ <= (others => '0');
        \$13819%now\ <= (others => '0');
        \$v7325%now\ <= (others => '0');
        \$13120%now\ <= (others => '0');
        \$v7087%now\ <= (others => '0');
        \$v6615%now\ <= (others => '0');
        \$15146_r%now\ <= (others => '0');
        \$v7394%now\ <= (others => '0');
        \$18347%now\ <= (others => '0');
        \$18700%now\ <= (others => '0');
        \$v6777%now\ <= (others => '0');
        \$12940%now\ <= (others => '0');
        \$v7173%now\ <= (others => '0');
        \$17062%now\ <= (others => '0');
        \$v7073%now\ <= (others => '0');
        \$14025_v%now\ <= (others => '0');
        \$14561%now\ <= (others => '0');
        \$16437_v%now\ <= (others => '0');
        \$15549_res%now\ <= (others => '0');
        \$15253_modulo6685896_arg%now\ <= (others => '0');
        \$15013_modulo6685896_arg%now\ <= (others => '0');
        \$14822_res%now\ <= (others => '0');
        \$18847%now\ <= (others => '0');
        \$18840%now\ <= (others => '0');
        \$18340_hd%now\ <= (others => '0');
        \$v7148%now\ <= (others => '0');
        \$14884_binop_int6435904_id%now\ <= (others => '0');
        \$18632_loop666_result%now\ <= (others => '0');
        \$15226_r%now\ <= (others => '0');
        \$18422%now\ <= (others => '0');
        \$15444%now\ <= (others => '0');
        \$19137%now\ <= (others => '0');
        \$18923%now\ <= (others => '0');
        \$17161%now\ <= (others => '0');
        \$12662%now\ <= (others => '0');
        \$v7065%now\ <= (others => '0');
        \$14662_res%now\ <= (others => '0');
        \$v6226%now\ <= (others => '0');
        \$v7319%now\ <= (others => '0');
        \$17396%now\ <= (others => '0');
        \$17806%now\ <= (others => '0');
        \$v6612%now\ <= (others => '0');
        \$15805_binop_compare6455921_id%now\ <= (others => '0');
        \$13305%now\ <= (others => '0');
        \$13230%now\ <= (others => '0');
        \$19056%now\ <= (others => '0');
        \$18469%now\ <= (others => '0');
        \$v7286%now\ <= (others => '0');
        \$13534%now\ <= (others => '0');
        \$v7152%now\ <= (others => '0');
        \$v6929%now\ <= (others => '0');
        \$16910_b%now\ <= (others => '0');
        \$v7043%now\ <= (others => '0');
        \$12850%now\ <= (others => '0');
        \$17456_loop665_id%now\ <= (others => '0');
        \$18477%now\ <= (others => '0');
        \$v7225%now\ <= (others => '0');
        \$v6923%now\ <= (others => '0');
        \$v6674%now\ <= (others => '0');
        \$13699%now\ <= (others => '0');
        \$v6944%now\ <= (others => '0');
        \$13923_make_block579_id%now\ <= (others => '0');
        \$14207_loop_push6495899_id%now\ <= (others => '0');
        \$15648_compare6445897_arg%now\ <= (others => '0');
        \$13803_w%now\ <= (others => '0');
        \$17780%now\ <= (others => '0');
        \$12876%now\ <= (others => '0');
        \$18656%now\ <= (others => '0');
        \$v6687%now\ <= (others => '0');
        \$v6107%now\ <= (others => '0');
        \$12661%now\ <= (others => '0');
        \$v6630%now\ <= (others => '0');
        \$15697_binop_compare6455918_id%now\ <= (others => '0');
        \$v7124%now\ <= (others => '0');
        \$v7384%now\ <= (others => '0');
        \$v7063%now\ <= (others => '0');
        \$13928_w652_arg%now\ <= (others => '0');
        \$15465_v%now\ <= (others => '0');
        \$13622%now\ <= (others => '0');
        \$14355%now\ <= (others => '0');
        \$v7312%now\ <= (others => '0');
        \$v6636%now\ <= (others => '0');
        \$14770_r%now\ <= (others => '0');
        \$v6063%now\ <= (others => '0');
        \$15013_modulo6685896_id%now\ <= (others => '0');
        \$14690_r%now\ <= (others => '0');
        \$12807_loop665_arg%now\ <= (others => '0');
        \$v6120%now\ <= (others => '0');
        \$17810%now\ <= (others => '0');
        \$v6168%now\ <= (others => '0');
        \$v7053%now\ <= (others => '0');
        \$v7239%now\ <= (others => '0');
        \$17236%now\ <= (others => '0');
        \$v7209%now\ <= (others => '0');
        \$13128%now\ <= (others => '0');
        \$15229_modulo6685895_id%now\ <= (others => '0');
        \$v7316%now\ <= (others => '0');
        \$12690%now\ <= (others => '0');
        \$13925_offsetclosure_n639_id%now\ <= (others => '0');
        \$13020%now\ <= (others => '0');
        \$v6932%now\ <= (others => '0');
        \$12539%now\ <= (others => '0');
        \$v6592%now\ <= (others => '0');
        \$v6010%now\ <= (others => '0');
        \$13093%now\ <= (others => '0');
        \$18323%now\ <= (others => '0');
        \$17965%now\ <= (others => '0');
        \$v5971%now\ <= (others => '0');
        \$16659_sp%now\ <= (others => '0');
        \$17547_copy_root_in_ram6635891_result%now\ <= (others => '0');
        \$13690%now\ <= (others => '0');
        \$13628%now\ <= (others => '0');
        \$v6349%now\ <= (others => '0');
        \$13465%now\ <= (others => '0');
        \$12812%now\ <= (others => '0');
        \$v6028%now\ <= (others => '0');
        \$13374_w%now\ <= (others => '0');
        \$14368%now\ <= (others => '0');
        \$12718%now\ <= (others => '0');
        \$17784%now\ <= (others => '0');
        \$15508_modulo6685888_id%now\ <= (others => '0');
        \$15364_binop_int6435910_result%now\ <= (others => '0');
        \$14613_modulo6685896_arg%now\ <= (others => '0');
        \$15751_res%now\ <= (others => '0');
        \$13537%now\ <= (others => '0');
        \$12654%now\ <= (others => '0');
        \$v7071%now\ <= (others => '0');
        \$v6311%now\ <= (others => '0');
        \$ram_lock%now\ <= (others => '0');
        \$global_end_lock%now\ <= (others => '0');
        \$code_lock%now\ <= (others => '0');
        \state%now\ <= idle5941;
        \state_var7464%now\ <= idle5976;
        \state_var7463%now\ <= idle6149;
        \state_var7462%now\ <= idle6114;
        \state_var7461%now\ <= idle6505;
        \state_var7460%now\ <= idle6470;
      elsif (rising_edge(clk)) then
        \$12559%now\ <= \$12559%next\;
        \$14060%now\ <= \$14060%next\;
        \$v6454%now\ <= \$v6454%next\;
        \$14516_v%now\ <= \$14516_v%next\;
        \$15069_modulo6685895_arg%now\ <= \$15069_modulo6685895_arg%next\;
        \$18421%now\ <= \$18421%next\;
        \$v6570%now\ <= \$v6570%next\;
        \$14564_binop_int6435900_arg%now\ <= \$14564_binop_int6435900_arg%next\;
        \$17813%now\ <= \$17813%next\;
        \$v6841%now\ <= \$v6841%next\;
        \$14666_r%now\ <= \$14666_r%next\;
        \$v7022%now\ <= \$v7022%next\;
        \$14589_modulo6685895_result%now\ <= \$14589_modulo6685895_result%next\;
        \$13392%now\ <= \$13392%next\;
        \$18996%now\ <= \$18996%next\;
        \$12673_rdy%now\ <= \$12673_rdy%next\;
        \$v6130%now\ <= \$v6130%next\;
        \$v7263%now\ <= \$v7263%next\;
        \$14917_modulo6685888_arg%now\ <= \$14917_modulo6685888_arg%next\;
        \$v6197%now\ <= \$v6197%next\;
        \$19272%now\ <= \$19272%next\;
        \$v7123%now\ <= \$v7123%next\;
        \$v6642%now\ <= \$v6642%next\;
        \$18729%now\ <= \$18729%next\;
        \$18192%now\ <= \$18192%next\;
        \$13670%now\ <= \$13670%next\;
        \$v6127%now\ <= \$v6127%next\;
        \$15675_v%now\ <= \$15675_v%next\;
        \$15077_modulo6685888_result%now\ <= \$15077_modulo6685888_result%next\;
        \$v6725%now\ <= \$v6725%next\;
        \$16182%now\ <= \$16182%next\;
        \$14052_v%now\ <= \$14052_v%next\;
        \$18354%now\ <= \$18354%next\;
        \$14749_modulo6685895_result%now\ <= \$14749_modulo6685895_result%next\;
        \$v6451%now\ <= \$v6451%next\;
        \$12545_x%now\ <= \$12545_x%next\;
        \$v7062%now\ <= \$v7062%next\;
        \$17496_next%now\ <= \$17496_next%next\;
        \$12852%now\ <= \$12852%next\;
        \$13503%now\ <= \$13503%next\;
        \$v6473%now\ <= \$v6473%next\;
        \$15531_binop_int6435913_arg%now\ <= \$15531_binop_int6435913_arg%next\;
        \$17887%now\ <= \$17887%next\;
        \$18997%now\ <= \$18997%next\;
        \$18835%now\ <= \$18835%next\;
        \$v6567%now\ <= \$v6567%next\;
        \$v7313%now\ <= \$v7313%next\;
        \$14724_binop_int6435902_result%now\ <= \$14724_binop_int6435902_result%next\;
        \$12699%now\ <= \$12699%next\;
        \$v7125%now\ <= \$v7125%next\;
        \$14989_modulo6685895_arg%now\ <= \$14989_modulo6685895_arg%next\;
        \$13090%now\ <= \$13090%next\;
        \$19003%now\ <= \$19003%next\;
        \$12522_wait662_arg%now\ <= \$12522_wait662_arg%next\;
        \$16811_compare6445898_arg%now\ <= \$16811_compare6445898_arg%next\;
        \$17893%now\ <= \$17893%next\;
        \$15661_binop_compare6455917_arg%now\ <= \$15661_binop_compare6455917_arg%next\;
        \$14126%now\ <= \$14126%next\;
        \$v7437%now\ <= \$v7437%next\;
        \$17570%now\ <= \$17570%next\;
        \$16453_v%now\ <= \$16453_v%next\;
        \$17676%now\ <= \$17676%next\;
        \$18121%now\ <= \$18121%next\;
        \$v7222%now\ <= \$v7222%next\;
        \$v6512%now\ <= \$v6512%next\;
        \$13308%now\ <= \$13308%next\;
        \$17018_w36575938_arg%now\ <= \$17018_w36575938_arg%next\;
        \$v6206%now\ <= \$v6206%next\;
        \$15484_modulo6685888_result%now\ <= \$15484_modulo6685888_result%next\;
        \$v7170%now\ <= \$v7170%next\;
        \$15614_forever6705914_arg%now\ <= \$15614_forever6705914_arg%next\;
        \$16858_compbranch6505932_arg%now\ <= \$16858_compbranch6505932_arg%next\;
        \$v7236%now\ <= \$v7236%next\;
        \$v7153%now\ <= \$v7153%next\;
        \$16893_compbranch6505933_id%now\ <= \$16893_compbranch6505933_id%next\;
        \$14597_modulo6685888_arg%now\ <= \$14597_modulo6685888_arg%next\;
        \$16141%now\ <= \$16141%next\;
        \$v6105%now\ <= \$v6105%next\;
        \$v7446%now\ <= \$v7446%next\;
        \$13156%now\ <= \$13156%next\;
        \$v6575%now\ <= \$v6575%next\;
        \$19138%now\ <= \$19138%next\;
        \$16178_v%now\ <= \$16178_v%next\;
        \$13945%now\ <= \$13945%next\;
        \$v7094%now\ <= \$v7094%next\;
        \$v6391%now\ <= \$v6391%next\;
        \$18838%now\ <= \$18838%next\;
        \$13824%now\ <= \$13824%next\;
        \$v6959%now\ <= \$v6959%next\;
        \$13531%now\ <= \$13531%next\;
        \$16788_compbranch6505930_arg%now\ <= \$16788_compbranch6505930_arg%next\;
        \$17971%now\ <= \$17971%next\;
        \$v6348%now\ <= \$v6348%next\;
        \$17121%now\ <= \$17121%next\;
        \$16752_fill6545929_arg%now\ <= \$16752_fill6545929_arg%next\;
        \$v6382%now\ <= \$v6382%next\;
        \$12853_forever6705887_arg%now\ <= \$12853_forever6705887_arg%next\;
        \$v7251%now\ <= \$v7251%next\;
        \$15769_binop_compare6455920_arg%now\ <= \$15769_binop_compare6455920_arg%next\;
        \$17494%now\ <= \$17494%next\;
        \$v6385%now\ <= \$v6385%next\;
        \$14326%now\ <= \$14326%next\;
        \$v6240%now\ <= \$v6240%next\;
        \$19080_next%now\ <= \$19080_next%next\;
        \$17386%now\ <= \$17386%next\;
        \$13982_v%now\ <= \$13982_v%next\;
        \$17459_loop665_arg%now\ <= \$17459_loop665_arg%next\;
        \$18719_w%now\ <= \$18719_w%next\;
        \$15445%now\ <= \$15445%next\;
        \$v7353%now\ <= \$v7353%next\;
        \$16752_fill6545929_result%now\ <= \$16752_fill6545929_result%next\;
        \$14997_modulo6685888_id%now\ <= \$14997_modulo6685888_id%next\;
        \$18050%now\ <= \$18050%next\;
        \$12883%now\ <= \$12883%next\;
        \$16823_compbranch6505931_arg%now\ <= \$16823_compbranch6505931_arg%next\;
        \$16233%now\ <= \$16233%next\;
        \$16271%now\ <= \$16271%next\;
        \$12682_make_block579_arg%now\ <= \$12682_make_block579_arg%next\;
        \$18655%now\ <= \$18655%next\;
        \$v7371%now\ <= \$v7371%next\;
        \$18987_hd%now\ <= \$18987_hd%next\;
        \$v6619%now\ <= \$v6619%next\;
        \$v6427%now\ <= \$v6427%next\;
        \$16748%now\ <= \$16748%next\;
        \$v6974%now\ <= \$v6974%next\;
        \$18474%now\ <= \$18474%next\;
        \$17886%now\ <= \$17886%next\;
        \$15756_compare6445897_arg%now\ <= \$15756_compare6445897_arg%next\;
        \$13151%now\ <= \$13151%next\;
        \$v6805%now\ <= \$v6805%next\;
        \$17569%now\ <= \$17569%next\;
        \$12698%now\ <= \$12698%next\;
        \$15389_modulo6685895_arg%now\ <= \$15389_modulo6685895_arg%next\;
        \$v6035%now\ <= \$v6035%next\;
        \$15553_r%now\ <= \$15553_r%next\;
        \$15237_modulo6685888_result%now\ <= \$15237_modulo6685888_result%next\;
        \$12944%now\ <= \$12944%next\;
        \$14613_modulo6685896_result%now\ <= \$14613_modulo6685896_result%next\;
        \$v7381%now\ <= \$v7381%next\;
        \$18846%now\ <= \$18846%next\;
        \$18917%now\ <= \$18917%next\;
        \$v6092%now\ <= \$v6092%next\;
        \$18916%now\ <= \$18916%next\;
        \$15261_modulo6685888_id%now\ <= \$15261_modulo6685888_id%next\;
        \$17679%now\ <= \$17679%next\;
        \$13154%now\ <= \$13154%next\;
        \$v6336%now\ <= \$v6336%next\;
        \$16527_f0%now\ <= \$16527_f0%next\;
        \$18352%now\ <= \$18352%next\;
        \$13964%now\ <= \$13964%next\;
        \$v7420%now\ <= \$v7420%next\;
        \$13632_next%now\ <= \$13632_next%next\;
        \$v6502%now\ <= \$v6502%next\;
        \$v6370%now\ <= \$v6370%next\;
        \$18739%now\ <= \$18739%next\;
        \$12714%now\ <= \$12714%next\;
        \$17484%now\ <= \$17484%next\;
        \$17597%now\ <= \$17597%next\;
        \$15756_compare6445897_result%now\ <= \$15756_compare6445897_result%next\;
        \$v7137%now\ <= \$v7137%next\;
        \$13532%now\ <= \$13532%next\;
        \$v6823%now\ <= \$v6823%next\;
        \$14781_modulo6685888_result%now\ <= \$14781_modulo6685888_result%next\;
        \$v6721%now\ <= \$v6721%next\;
        \$17734_copy_root_in_ram6635892_id%now\ <= \$17734_copy_root_in_ram6635892_id%next\;
        \$v7338%now\ <= \$v7338%next\;
        \$14749_modulo6685895_arg%now\ <= \$14749_modulo6685895_arg%next\;
        \$v7050%now\ <= \$v7050%next\;
        \$16299_v%now\ <= \$16299_v%next\;
        \$12689%now\ <= \$12689%next\;
        \$18807%now\ <= \$18807%next\;
        \$13920_loop666_arg%now\ <= \$13920_loop666_arg%next\;
        \$17455_loop666_id%now\ <= \$17455_loop666_id%next\;
        \$v6027%now\ <= \$v6027%next\;
        \$18650%now\ <= \$18650%next\;
        \$18837%now\ <= \$18837%next\;
        \$16951_compare6445898_arg%now\ <= \$16951_compare6445898_arg%next\;
        \$14861_modulo6685888_result%now\ <= \$14861_modulo6685888_result%next\;
        \$18805%now\ <= \$18805%next\;
        \$17543%now\ <= \$17543%next\;
        \$13997_v%now\ <= \$13997_v%next\;
        \$16574_compare6445898_id%now\ <= \$16574_compare6445898_id%next\;
        \$v6728%now\ <= \$v6728%next\;
        \$v6500%now\ <= \$v6500%next\;
        \$v5869%now\ <= \$v5869%next\;
        \$v6496%now\ <= \$v6496%next\;
        \$14978_v%now\ <= \$14978_v%next\;
        \$v7454%now\ <= \$v7454%next\;
        \$13237%now\ <= \$13237%next\;
        \$v6146%now\ <= \$v6146%next\;
        \$15330_r%now\ <= \$15330_r%next\;
        \$12839%now\ <= \$12839%next\;
        \$14061_v%now\ <= \$14061_v%next\;
        \$14701_modulo6685888_arg%now\ <= \$14701_modulo6685888_arg%next\;
        \$12697%now\ <= \$12697%next\;
        \$17773%now\ <= \$17773%next\;
        \$v7344%now\ <= \$v7344%next\;
        \$12888%now\ <= \$12888%next\;
        \$13155%now\ <= \$13155%next\;
        \$12937%now\ <= \$12937%next\;
        \$16115%now\ <= \$16115%next\;
        \$12805_aux664_result%now\ <= \$12805_aux664_result%next\;
        \$v6021%now\ <= \$v6021%next\;
        \$13697%now\ <= \$13697%next\;
        \$v6466%now\ <= \$v6466%next\;
        \$18355%now\ <= \$18355%next\;
        \rdy5940%now\ <= \rdy5940%next\;
        \$13102%now\ <= \$13102%next\;
        \$13235%now\ <= \$13235%next\;
        \$15044_binop_int6435906_id%now\ <= \$15044_binop_int6435906_id%next\;
        \$16729_v%now\ <= \$16729_v%next\;
        \$v6376%now\ <= \$v6376%next\;
        \$13233%now\ <= \$13233%next\;
        \$17670%now\ <= \$17670%next\;
        \$14555%now\ <= \$14555%next\;
        \$14564_binop_int6435900_result%now\ <= \$14564_binop_int6435900_result%next\;
        \$v6802%now\ <= \$v6802%next\;
        \$15058_v%now\ <= \$15058_v%next\;
        \$17464%now\ <= \$17464%next\;
        \$v6599%now\ <= \$v6599%next\;
        \$v6430%now\ <= \$v6430%next\;
        \$v6318%now\ <= \$v6318%next\;
        \$v7161%now\ <= \$v7161%next\;
        \$17669%now\ <= \$17669%next\;
        \$16963_compbranch6505935_id%now\ <= \$16963_compbranch6505935_id%next\;
        \$13967_v%now\ <= \$13967_v%next\;
        \$13696%now\ <= \$13696%next\;
        \$v6015%now\ <= \$v6015%next\;
        \$15476_modulo6685895_arg%now\ <= \$15476_modulo6685895_arg%next\;
        \$17470%now\ <= \$17470%next\;
        \$12520_loop666_id%now\ <= \$12520_loop666_id%next\;
        \$18815%now\ <= \$18815%next\;
        \$v6559%now\ <= \$v6559%next\;
        \$18565%now\ <= \$18565%next\;
        \$16551_compbranch6505926_id%now\ <= \$16551_compbranch6505926_id%next\;
        \$15397_modulo6685888_result%now\ <= \$15397_modulo6685888_result%next\;
        \$12877%now\ <= \$12877%next\;
        \$18698%now\ <= \$18698%next\;
        \$18480%now\ <= \$18480%next\;
        \$v7300%now\ <= \$v7300%next\;
        \$15389_modulo6685895_result%now\ <= \$15389_modulo6685895_result%next\;
        \$v7144%now\ <= \$v7144%next\;
        \$v6780%now\ <= \$v6780%next\;
        \$19256_hd%now\ <= \$19256_hd%next\;
        \$15823_res%now\ <= \$15823_res%next\;
        \$15124_binop_int6435907_id%now\ <= \$15124_binop_int6435907_id%next\;
        \$v6218%now\ <= \$v6218%next\;
        \$v7406%now\ <= \$v7406%next\;
        \$16963_compbranch6505935_arg%now\ <= \$16963_compbranch6505935_arg%next\;
        \$v7132%now\ <= \$v7132%next\;
        \$v7200%now\ <= \$v7200%next\;
        \$18633_loop665_id%now\ <= \$18633_loop665_id%next\;
        \$17888%now\ <= \$17888%next\;
        \$19145%now\ <= \$19145%next\;
        \$15625_binop_compare6455916_id%now\ <= \$15625_binop_compare6455916_id%next\;
        \$19337%now\ <= \$19337%next\;
        \$15893%now\ <= \$15893%next\;
        \$14364_v%now\ <= \$14364_v%next\;
        \$16893_compbranch6505933_result%now\ <= \$16893_compbranch6505933_result%next\;
        \$v6406%now\ <= \$v6406%next\;
        \$v6489%now\ <= \$v6489%next\;
        \$14837_modulo6685888_result%now\ <= \$14837_modulo6685888_result%next\;
        \$14677_modulo6685888_arg%now\ <= \$14677_modulo6685888_arg%next\;
        \$v6667%now\ <= \$v6667%next\;
        \$v7413%now\ <= \$v7413%next\;
        \$v6508%now\ <= \$v6508%next\;
        \$v6591%now\ <= \$v6591%next\;
        \$16284_v%now\ <= \$16284_v%next\;
        \$12808_aux664_result%now\ <= \$12808_aux664_result%next\;
        \$13816%now\ <= \$13816%next\;
        \$v6211%now\ <= \$v6211%next\;
        \$15874%now\ <= \$15874%next\;
        \$14829_modulo6685895_id%now\ <= \$14829_modulo6685895_id%next\;
        \$v7027%now\ <= \$v7027%next\;
        \$v6596%now\ <= \$v6596%next\;
        \$17746%now\ <= \$17746%next\;
        \$13950%now\ <= \$13950%next\;
        \$v5963%now\ <= \$v5963%next\;
        \$v5944%now\ <= \$v5944%next\;
        \$14597_modulo6685888_result%now\ <= \$14597_modulo6685888_result%next\;
        \$14582_res%now\ <= \$14582_res%next\;
        \$17891%now\ <= \$17891%next\;
        \$15397_modulo6685888_arg%now\ <= \$15397_modulo6685888_arg%next\;
        \$13927_branch_if648_result%now\ <= \$13927_branch_if648_result%next\;
        \$v7306%now\ <= \$v7306%next\;
        \$v7074%now\ <= \$v7074%next\;
        \$15021_modulo6685888_result%now\ <= \$15021_modulo6685888_result%next\;
        \$12707%now\ <= \$12707%next\;
        \$16881_compare6445898_result%now\ <= \$16881_compare6445898_result%next\;
        \$13679_w%now\ <= \$13679_w%next\;
        \$13663%now\ <= \$13663%next\;
        \$18447%now\ <= \$18447%next\;
        \$v6732%now\ <= \$v6732%next\;
        \$v6298%now\ <= \$v6298%next\;
        \$v6518%now\ <= \$v6518%next\;
        \$18278%now\ <= \$18278%next\;
        \$12544%now\ <= \$12544%next\;
        \$13218_w%now\ <= \$13218_w%next\;
        \$15932%now\ <= \$15932%next\;
        \$v7402%now\ <= \$v7402%next\;
        \$v7085%now\ <= \$v7085%next\;
        \$18731%now\ <= \$18731%next\;
        \$13519_w%now\ <= \$13519_w%next\;
        \$13606%now\ <= \$13606%next\;
        \$17776%now\ <= \$17776%next\;
        \$18644%now\ <= \$18644%next\;
        \$16327%now\ <= \$16327%next\;
        \$16169_v%now\ <= \$16169_v%next\;
        \$16551_compbranch6505926_arg%now\ <= \$16551_compbranch6505926_arg%next\;
        \$15229_modulo6685895_arg%now\ <= \$15229_modulo6685895_arg%next\;
        \$17457_aux664_result%now\ <= \$17457_aux664_result%next\;
        \$v6633%now\ <= \$v6633%next\;
        \$17665_hd%now\ <= \$17665_hd%next\;
        \$18159%now\ <= \$18159%next\;
        \$v6058%now\ <= \$v6058%next\;
        \$14122%now\ <= \$14122%next\;
        \$18563%now\ <= \$18563%next\;
        \$13310%now\ <= \$13310%next\;
        \$14012%now\ <= \$14012%next\;
        \$14677_modulo6685888_id%now\ <= \$14677_modulo6685888_id%next\;
        \$14181_sp%now\ <= \$14181_sp%next\;
        \$v6235%now\ <= \$v6235%next\;
        \$15961%now\ <= \$15961%next\;
        \$15476_modulo6685895_result%now\ <= \$15476_modulo6685895_result%next\;
        \$15237_modulo6685888_id%now\ <= \$15237_modulo6685888_id%next\;
        \$17505_forever6705894_arg%now\ <= \$17505_forever6705894_arg%next\;
        \$13388%now\ <= \$13388%next\;
        \$v6480%now\ <= \$v6480%next\;
        \$17001%now\ <= \$17001%next\;
        \$17963%now\ <= \$17963%next\;
        \$17803%now\ <= \$17803%next\;
        \$19142%now\ <= \$19142%next\;
        \$18679_forever6705881_id%now\ <= \$18679_forever6705881_id%next\;
        \$v6291%now\ <= \$v6291%next\;
        \$v6532%now\ <= \$v6532%next\;
        \$v7293%now\ <= \$v7293%next\;
        \$18919%now\ <= \$18919%next\;
        \$12685%now\ <= \$12685%next\;
        \$v6501%now\ <= \$v6501%next\;
        \$17238_sp%now\ <= \$17238_sp%next\;
        \$18186%now\ <= \$18186%next\;
        \$v7279%now\ <= \$v7279%next\;
        \$v6460%now\ <= \$v6460%next\;
        \$14431%now\ <= \$14431%next\;
        \$13667%now\ <= \$13667%next\;
        \$17455_loop666_arg%now\ <= \$17455_loop666_arg%next\;
        \$12851%now\ <= \$12851%next\;
        \$18188%now\ <= \$18188%next\;
        \$v6172%now\ <= \$v6172%next\;
        \$v7403%now\ <= \$v7403%next\;
        \$v7216%now\ <= \$v7216%next\;
        \$v7035%now\ <= \$v7035%next\;
        \$v6397%now\ <= \$v6397%next\;
        \$18709%now\ <= \$18709%next\;
        \$15720_compare6445897_id%now\ <= \$15720_compare6445897_id%next\;
        \$13823%now\ <= \$13823%next\;
        \$14177_hd%now\ <= \$14177_hd%next\;
        \result6503%now\ <= \result6503%next\;
        \$13395%now\ <= \$13395%next\;
        \$16353%now\ <= \$16353%next\;
        \$v6239%now\ <= \$v6239%next\;
        \$17559%now\ <= \$17559%next\;
        \$14351_v%now\ <= \$14351_v%next\;
        \$12808_aux664_id%now\ <= \$12808_aux664_id%next\;
        \$19269%now\ <= \$19269%next\;
        \$17412%now\ <= \$17412%next\;
        \$v7007%now\ <= \$v7007%next\;
        \$v6941%now\ <= \$v6941%next\;
        \$v6746%now\ <= \$v6746%next\;
        \$18925%now\ <= \$18925%next\;
        \$v6838%now\ <= \$v6838%next\;
        \$18733%now\ <= \$18733%next\;
        \$v5957%now\ <= \$v5957%next\;
        \$v6953%now\ <= \$v6953%next\;
        \$15783_v%now\ <= \$15783_v%next\;
        \$18279%now\ <= \$18279%next\;
        \$14207_loop_push6495899_result%now\ <= \$14207_loop_push6495899_result%next\;
        \$v6108%now\ <= \$v6108%next\;
        \$v7025%now\ <= \$v7025%next\;
        \$18120%now\ <= \$18120%next\;
        \$18566%now\ <= \$18566%next\;
        \$13016%now\ <= \$13016%next\;
        \$v6304%now\ <= \$v6304%next\;
        \$12692%now\ <= \$12692%next\;
        \$16037_v%now\ <= \$16037_v%next\;
        \$12935%now\ <= \$12935%next\;
        \$13625%now\ <= \$13625%next\;
        \$v7434%now\ <= \$v7434%next\;
        \$v6739%now\ <= \$v6739%next\;
        \$17509_forever6705890_arg%now\ <= \$17509_forever6705890_arg%next\;
        \$v6274%now\ <= \$v6274%next\;
        \$19001%now\ <= \$19001%next\;
        \$v7290%now\ <= \$v7290%next\;
        \$17498%now\ <= \$17498%next\;
        \$16945_b%now\ <= \$16945_b%next\;
        \$15298_v%now\ <= \$15298_v%next\;
        \$18346%now\ <= \$18346%next\;
        \$16589_compbranch6505927_id%now\ <= \$16589_compbranch6505927_id%next\;
        \$v6708%now\ <= \$v6708%next\;
        \$13157%now\ <= \$13157%next\;
        \$18909_hd%now\ <= \$18909_hd%next\;
        \$17674%now\ <= \$17674%next\;
        \$12712%now\ <= \$12712%next\;
        \$12945%now\ <= \$12945%next\;
        \$17354%now\ <= \$17354%next\;
        \$16574_compare6445898_result%now\ <= \$16574_compare6445898_result%next\;
        \$16365%now\ <= \$16365%next\;
        \$12715%now\ <= \$12715%next\;
        \$16510_forever6705925_id%now\ <= \$16510_forever6705925_id%next\;
        \$15218_v%now\ <= \$15218_v%next\;
        \$18699%now\ <= \$18699%next\;
        \$17591%now\ <= \$17591%next\;
        \$v6627%now\ <= \$v6627%next\;
        \$12915%now\ <= \$12915%next\;
        \$v6136%now\ <= \$v6136%next\;
        \$18045%now\ <= \$18045%next\;
        \$17460_aux664_id%now\ <= \$17460_aux664_id%next\;
        \$12807_loop665_id%now\ <= \$12807_loop665_id%next\;
        \$15069_modulo6685895_id%now\ <= \$15069_modulo6685895_id%next\;
        \$v6492%now\ <= \$v6492%next\;
        \$17487%now\ <= \$17487%next\;
        \$v6892%now\ <= \$v6892%next\;
        \$17387%now\ <= \$17387%next\;
        \$15386_r%now\ <= \$15386_r%next\;
        \$v6729%now\ <= \$v6729%next\;
        \$v6914%now\ <= \$v6914%next\;
        \$18915%now\ <= \$18915%next\;
        \$17105_w06555936_id%now\ <= \$17105_w06555936_id%next\;
        \$16589_compbranch6505927_arg%now\ <= \$16589_compbranch6505927_arg%next\;
        \$13890%now\ <= \$13890%next\;
        \$19144%now\ <= \$19144%next\;
        \$16677%now\ <= \$16677%next\;
        \$v7034%now\ <= \$v7034%next\;
        \$17678%now\ <= \$17678%next\;
        \$16875_b%now\ <= \$16875_b%next\;
        \$13927_branch_if648_arg%now\ <= \$13927_branch_if648_arg%next\;
        \$v6883%now\ <= \$v6883%next\;
        \$16438_v%now\ <= \$16438_v%next\;
        \$15612%now\ <= \$15612%next\;
        \$14773_modulo6685896_arg%now\ <= \$14773_modulo6685896_arg%next\;
        \$19140%now\ <= \$19140%next\;
        \$19071%now\ <= \$19071%next\;
        \$12848%now\ <= \$12848%next\;
        \$18831_hd%now\ <= \$18831_hd%next\;
        \$v6710%now\ <= \$v6710%next\;
        \$13468%now\ <= \$13468%next\;
        \$v6856%now\ <= \$v6856%next\;
        \$15317_modulo6685888_result%now\ <= \$15317_modulo6685888_result%next\;
        \$18570%now\ <= \$18570%next\;
        \$13623%now\ <= \$13623%next\;
        \$18128_next%now\ <= \$18128_next%next\;
        \$v7248%now\ <= \$v7248%next\;
        \$14644_binop_int6435901_result%now\ <= \$14644_binop_int6435901_result%next\;
        \$12679_loop666_id%now\ <= \$12679_loop666_id%next\;
        \$16399%now\ <= \$16399%next\;
        \$19263%now\ <= \$19263%next\;
        \$14749_modulo6685895_id%now\ <= \$14749_modulo6685895_id%next\;
        \$17794_w%now\ <= \$17794_w%next\;
        \result6468%now\ <= \result6468%next\;
        \$v7045%now\ <= \$v7045%next\;
        \$18816%now\ <= \$18816%next\;
        \$17885%now\ <= \$17885%next\;
        \$v7164%now\ <= \$v7164%next\;
        \$15101_modulo6685888_result%now\ <= \$15101_modulo6685888_result%next\;
        \$v7042%now\ <= \$v7042%next\;
        \$15500_modulo6685896_arg%now\ <= \$15500_modulo6685896_arg%next\;
        \$15333_modulo6685896_result%now\ <= \$15333_modulo6685896_result%next\;
        \$17761_copy_root_in_ram6635891_result%now\ <= \$17761_copy_root_in_ram6635891_result%next\;
        \$15720_compare6445897_arg%now\ <= \$15720_compare6445897_arg%next\;
        \$16713_v%now\ <= \$16713_v%next\;
        \$15697_binop_compare6455918_arg%now\ <= \$15697_binop_compare6455918_arg%next\;
        \$17250_v%now\ <= \$17250_v%next\;
        \$12887%now\ <= \$12887%next\;
        \$v6826%now\ <= \$v6826%next\;
        \$17394%now\ <= \$17394%next\;
        \$v6695%now\ <= \$v6695%next\;
        \$17333_sp%now\ <= \$17333_sp%next\;
        \$v7017%now\ <= \$v7017%next\;
        \$16158_forever6705923_arg%now\ <= \$16158_forever6705923_arg%next\;
        \$v6874%now\ <= \$v6874%next\;
        \$v6574%now\ <= \$v6574%next\;
        \$15853_v%now\ <= \$15853_v%next\;
        \$v7372%now\ <= \$v7372%next\;
        \$v6651%now\ <= \$v6651%next\;
        \$v7013%now\ <= \$v7013%next\;
        \$15181_modulo6685888_result%now\ <= \$15181_modulo6685888_result%next\;
        \$12691%now\ <= \$12691%next\;
        \$17962%now\ <= \$17962%next\;
        \$v6367%now\ <= \$v6367%next\;
        \$v6200%now\ <= \$v6200%next\;
        \$16612_compare6445898_result%now\ <= \$16612_compare6445898_result%next\;
        \$v6688%now\ <= \$v6688%next\;
        \$14330_v%now\ <= \$14330_v%next\;
        \$v7361%now\ <= \$v7361%next\;
        \$17319%now\ <= \$17319%next\;
        \$13941%now\ <= \$13941%next\;
        \$16078%now\ <= \$16078%next\;
        \$16165%now\ <= \$16165%next\;
        \$v7299%now\ <= \$v7299%next\;
        \$17012_sp%now\ <= \$17012_sp%next\;
        \$15261_modulo6685888_arg%now\ <= \$15261_modulo6685888_arg%next\;
        \$v6342%now\ <= \$v6342%next\;
        \$v5954%now\ <= \$v5954%next\;
        \$16606_b%now\ <= \$16606_b%next\;
        \$14986_r%now\ <= \$14986_r%next\;
        \$13301_hd%now\ <= \$13301_hd%next\;
        \$15847%now\ <= \$15847%next\;
        \$v7179%now\ <= \$v7179%next\;
        \$15021_modulo6685888_arg%now\ <= \$15021_modulo6685888_arg%next\;
        \$13127%now\ <= \$13127%next\;
        \$v7004%now\ <= \$v7004%next\;
        \$v7090%now\ <= \$v7090%next\;
        \$v6709%now\ <= \$v6709%next\;
        \$17321%now\ <= \$17321%next\;
        \$13530%now\ <= \$13530%next\;
        \$14222%now\ <= \$14222%next\;
        \$v6868%now\ <= \$v6868%next\;
        \$v6203%now\ <= \$v6203%next\;
        \$v5866%now\ <= \$v5866%next\;
        \$v5951%now\ <= \$v5951%next\;
        \$18450%now\ <= \$18450%next\;
        \$13296_w%now\ <= \$13296_w%next\;
        \$14724_binop_int6435902_id%now\ <= \$14724_binop_int6435902_id%next\;
        \$v7400%now\ <= \$v7400%next\;
        \$13013%now\ <= \$13013%next\;
        \$17349%now\ <= \$17349%next\;
        \$16192%now\ <= \$16192%next\;
        \$12834%now\ <= \$12834%next\;
        \$16441%now\ <= \$16441%next\;
        \$17167%now\ <= \$17167%next\;
        \$16042_v%now\ <= \$16042_v%next\;
        \$15697_binop_compare6455918_result%now\ <= \$15697_binop_compare6455918_result%next\;
        \$12679_loop666_result%now\ <= \$12679_loop666_result%next\;
        \$16234%now\ <= \$16234%next\;
        \$15625_binop_compare6455916_result%now\ <= \$15625_binop_compare6455916_result%next\;
        \$v7140%now\ <= \$v7140%next\;
        \$18163%now\ <= \$18163%next\;
        \$v6007%now\ <= \$v6007%next\;
        \$14933_modulo6685896_result%now\ <= \$14933_modulo6685896_result%next\;
        \$v7066%now\ <= \$v7066%next\;
        \$14818_v%now\ <= \$14818_v%next\;
        \$v6750%now\ <= \$v6750%next\;
        \$15976_v%now\ <= \$15976_v%next\;
        \$v6935%now\ <= \$v6935%next\;
        \$14338_v%now\ <= \$14338_v%next\;
        \$v6986%now\ <= \$v6986%next\;
        \$16805_b%now\ <= \$16805_b%next\;
        \$17961%now\ <= \$17961%next\;
        \$16439_v%now\ <= \$16439_v%next\;
        \$14933_modulo6685896_id%now\ <= \$14933_modulo6685896_id%next\;
        \$17681%now\ <= \$17681%next\;
        \$12910%now\ <= \$12910%next\;
        \$v6445%now\ <= \$v6445%next\;
        \$12741%now\ <= \$12741%next\;
        \$v7455%now\ <= \$v7455%next\;
        \$v6277%now\ <= \$v6277%next\;
        \$v6962%now\ <= \$v6962%next\;
        \$v7441%now\ <= \$v7441%next\;
        \$13962%now\ <= \$13962%next\;
        \$15010_r%now\ <= \$15010_r%next\;
        \$14829_modulo6685895_result%now\ <= \$14829_modulo6685895_result%next\;
        \$12521_loop665_arg%now\ <= \$12521_loop665_arg%next\;
        \$14161%now\ <= \$14161%next\;
        \$15805_binop_compare6455921_arg%now\ <= \$15805_binop_compare6455921_arg%next\;
        \$12843%now\ <= \$12843%next\;
        \$15413_modulo6685896_result%now\ <= \$15413_modulo6685896_result%next\;
        \$v7064%now\ <= \$v7064%next\;
        \$15484_modulo6685888_arg%now\ <= \$15484_modulo6685888_arg%next\;
        \$v7368%now\ <= \$v7368%next\;
        \$v6117%now\ <= \$v6117%next\;
        \$18634_aux664_result%now\ <= \$18634_aux664_result%next\;
        \$12943%now\ <= \$12943%next\;
        \$v6995%now\ <= \$v6995%next\;
        \$v6657%now\ <= \$v6657%next\;
        \$17600%now\ <= \$17600%next\;
        \$v6214%now\ <= \$v6214%next\;
        \$13957%now\ <= \$13957%next\;
        \$v7016%now\ <= \$v7016%next\;
        \$v6307%now\ <= \$v6307%next\;
        \$v6268%now\ <= \$v6268%next\;
        \$18982_w%now\ <= \$18982_w%next\;
        \$13103%now\ <= \$13103%next\;
        \$14517_v%now\ <= \$14517_v%next\;
        \$v7023%now\ <= \$v7023%next\;
        \$13692%now\ <= \$13692%next\;
        \$18479%now\ <= \$18479%next\;
        \$v7358%now\ <= \$v7358%next\;
        \$v6271%now\ <= \$v6271%next\;
        \$v6681%now\ <= \$v6681%next\;
        \$12806_loop666_result%now\ <= \$12806_loop666_result%next\;
        \$12680_loop665_result%now\ <= \$12680_loop665_result%next\;
        \$18734%now\ <= \$18734%next\;
        \$15484_modulo6685888_id%now\ <= \$15484_modulo6685888_id%next\;
        \$v6055%now\ <= \$v6055%next\;
        \$14746_r%now\ <= \$14746_r%next\;
        \$17327%now\ <= \$17327%next\;
        \$13153%now\ <= \$13153%next\;
        \$v6701%now\ <= \$v6701%next\;
        \$v7453%now\ <= \$v7453%next\;
        \$v6950%now\ <= \$v6950%next\;
        \$15733_binop_compare6455919_arg%now\ <= \$15733_binop_compare6455919_arg%next\;
        \$16436_v%now\ <= \$16436_v%next\;
        \$v7335%now\ <= \$v7335%next\;
        \$14837_modulo6685888_arg%now\ <= \$14837_modulo6685888_arg%next\;
        \$14558%now\ <= \$14558%next\;
        \$v6609%now\ <= \$v6609%next\;
        \$v6102%now\ <= \$v6102%next\;
        \$v6865%now\ <= \$v6865%next\;
        \$v7121%now\ <= \$v7121%next\;
        \$v6175%now\ <= \$v6175%next\;
        \$17520_copy_root_in_ram6635893_id%now\ <= \$17520_copy_root_in_ram6635893_id%next\;
        \$18818%now\ <= \$18818%next\;
        \$17018_w36575938_id%now\ <= \$17018_w36575938_id%next\;
        \$13946%now\ <= \$13946%next\;
        \$v7354%now\ <= \$v7354%next\;
        \$17315%now\ <= \$17315%next\;
        \$15204_binop_int6435908_id%now\ <= \$15204_binop_int6435908_id%next\;
        \$14658_v%now\ <= \$14658_v%next\;
        \$13307%now\ <= \$13307%next\;
        \$14042%now\ <= \$14042%next\;
        \$12939%now\ <= \$12939%next\;
        \$12891_copy_root_in_ram6635884_arg%now\ <= \$12891_copy_root_in_ram6635884_arg%next\;
        \$v7416%now\ <= \$v7416%next\;
        \$18166%now\ <= \$18166%next\;
        \$15556_modulo6685895_result%now\ <= \$15556_modulo6685895_result%next\;
        \$16035%now\ <= \$16035%next\;
        \$14853_modulo6685896_arg%now\ <= \$14853_modulo6685896_arg%next\;
        \$15124_binop_int6435907_arg%now\ <= \$15124_binop_int6435907_arg%next\;
        \$13928_w652_result%now\ <= \$13928_w652_result%next\;
        \$15317_modulo6685888_arg%now\ <= \$15317_modulo6685888_arg%next\;
        \$17377%now\ <= \$17377%next\;
        \$16126%now\ <= \$16126%next\;
        \$v7133%now\ <= \$v7133%next\;
        \$16127_v%now\ <= \$16127_v%next\;
        \$12878%now\ <= \$12878%next\;
        \$16031%now\ <= \$16031%next\;
        \$18836%now\ <= \$18836%next\;
        \$12857_forever6705883_arg%now\ <= \$12857_forever6705883_arg%next\;
        \$v7219%now\ <= \$v7219%next\;
        \$v6773%now\ <= \$v6773%next\;
        \$14114%now\ <= \$14114%next\;
        \$v7086%now\ <= \$v7086%next\;
        \$18999%now\ <= \$18999%next\;
        \$18637%now\ <= \$18637%next\;
        \$v6301%now\ <= \$v6301%next\;
        \$17734_copy_root_in_ram6635892_arg%now\ <= \$17734_copy_root_in_ram6635892_arg%next\;
        \$v5874%now\ <= \$v5874%next\;
        \$v7185%now\ <= \$v7185%next\;
        \$13693%now\ <= \$13693%next\;
        \$v6229%now\ <= \$v6229%next\;
        \$14285_v%now\ <= \$14285_v%next\;
        \$12734%now\ <= \$12734%next\;
        \$15341_modulo6685888_arg%now\ <= \$15341_modulo6685888_arg%next\;
        \$12904%now\ <= \$12904%next\;
        \$v7077%now\ <= \$v7077%next\;
        \$17513_forever6705889_id%now\ <= \$17513_forever6705889_id%next\;
        \$v6853%now\ <= \$v6853%next\;
        \$13466%now\ <= \$13466%next\;
        \$v7322%now\ <= \$v7322%next\;
        \$14804_binop_int6435903_arg%now\ <= \$14804_binop_int6435903_arg%next\;
        \$17463%now\ <= \$17463%next\;
        \$19115%now\ <= \$19115%next\;
        \$18904_w%now\ <= \$18904_w%next\;
        \$12818%now\ <= \$12818%next\;
        \$v6751%now\ <= \$v6751%next\;
        \$16292%now\ <= \$16292%next\;
        \$12844_next%now\ <= \$12844_next%next\;
        \$16395_v%now\ <= \$16395_v%next\;
        \$14964_binop_int6435905_id%now\ <= \$14964_binop_int6435905_id%next\;
        \$16767%now\ <= \$16767%next\;
        \$15093_modulo6685896_arg%now\ <= \$15093_modulo6685896_arg%next\;
        \$v6103%now\ <= \$v6103%next\;
        \$15648_compare6445897_id%now\ <= \$15648_compare6445897_id%next\;
        \$v6165%now\ <= \$v6165%next\;
        \$18104%now\ <= \$18104%next\;
        \$v7030%now\ <= \$v7030%next\;
        \$14613_modulo6685896_id%now\ <= \$14613_modulo6685896_id%next\;
        \$v6738%now\ <= \$v6738%next\;
        \$v6678%now\ <= \$v6678%next\;
        \$17491%now\ <= \$17491%next\;
        \$13078_copy_root_in_ram6635885_id%now\ <= \$13078_copy_root_in_ram6635885_id%next\;
        \$15981_v%now\ <= \$15981_v%next\;
        \$12560%now\ <= \$12560%next\;
        \$v7057%now\ <= \$v7057%next\;
        \$v6364%now\ <= \$v6364%next\;
        \$12702%now\ <= \$12702%next\;
        \$13312%now\ <= \$13312%next\;
        \$12520_loop666_arg%now\ <= \$12520_loop666_arg%next\;
        \$15792_compare6445897_result%now\ <= \$15792_compare6445897_result%next\;
        \$15341_modulo6685888_result%now\ <= \$15341_modulo6685888_result%next\;
        \$v7076%now\ <= \$v7076%next\;
        \$14669_modulo6685895_id%now\ <= \$14669_modulo6685895_id%next\;
        \$v5878%now\ <= \$v5878%next\;
        \$18711%now\ <= \$18711%next\;
        \$15828_compare6445897_id%now\ <= \$15828_compare6445897_id%next\;
        \$15237_modulo6685888_arg%now\ <= \$15237_modulo6685888_arg%next\;
        \$v6183%now\ <= \$v6183%next\;
        \$v5992%now\ <= \$v5992%next\;
        \$v6314%now\ <= \$v6314%next\;
        \$12522_wait662_result%now\ <= \$12522_wait662_result%next\;
        \$v6947%now\ <= \$v6947%next\;
        \$v6595%now\ <= \$v6595%next\;
        \$17455_loop666_result%now\ <= \$17455_loop666_result%next\;
        \$v7458%now\ <= \$v7458%next\;
        \$v6162%now\ <= \$v6162%next\;
        \$12838_next%now\ <= \$12838_next%next\;
        \$v6012%now\ <= \$v6012%next\;
        \$18472%now\ <= \$18472%next\;
        \$16036_sp%now\ <= \$16036_sp%next\;
        \$18185%now\ <= \$18185%next\;
        \$14424_v%now\ <= \$14424_v%next\;
        \$14254%now\ <= \$14254%next\;
        \$13389%now\ <= \$13389%next\;
        \$18677%now\ <= \$18677%next\;
        \$17348%now\ <= \$17348%next\;
        \$13393%now\ <= \$13393%next\;
        \$15769_binop_compare6455920_id%now\ <= \$15769_binop_compare6455920_id%next\;
        \$13387%now\ <= \$13387%next\;
        \$17590%now\ <= \$17590%next\;
        \$v7398%now\ <= \$v7398%next\;
        \$16823_compbranch6505931_id%now\ <= \$16823_compbranch6505931_id%next\;
        \$17495%now\ <= \$17495%next\;
        \$16379_v%now\ <= \$16379_v%next\;
        \$16881_compare6445898_arg%now\ <= \$16881_compare6445898_arg%next\;
        \$18679_forever6705881_arg%now\ <= \$18679_forever6705881_arg%next\;
        \$v6048%now\ <= \$v6048%next\;
        \$14677_modulo6685888_result%now\ <= \$14677_modulo6685888_result%next\;
        \$18288_next%now\ <= \$18288_next%next\;
        \$12538_cy%now\ <= \$12538_cy%next\;
        \$15378_v%now\ <= \$15378_v%next\;
        \$12941%now\ <= \$12941%next\;
        \$17783%now\ <= \$17783%next\;
        \$13794%now\ <= \$13794%next\;
        \$14693_modulo6685896_arg%now\ <= \$14693_modulo6685896_arg%next\;
        \$12914%now\ <= \$12914%next\;
        \$19262%now\ <= \$19262%next\;
        \$v6847%now\ <= \$v6847%next\;
        \$15382_res%now\ <= \$15382_res%next\;
        \$12521_loop665_result%now\ <= \$12521_loop665_result%next\;
        \$13238%now\ <= \$13238%next\;
        \$v6286%now\ <= \$v6286%next\;
        \$19070%now\ <= \$19070%next\;
        \$17254%now\ <= \$17254%next\;
        \$13694%now\ <= \$13694%next\;
        \$14941_modulo6685888_arg%now\ <= \$14941_modulo6685888_arg%next\;
        \$v7328%now\ <= \$v7328%next\;
        \$18356%now\ <= \$18356%next\;
        \$v7054%now\ <= \$v7054%next\;
        \$17761_copy_root_in_ram6635891_id%now\ <= \$17761_copy_root_in_ram6635891_id%next\;
        \$12695%now\ <= \$12695%next\;
        \$v6089%now\ <= \$v6089%next\;
        \$17774%now\ <= \$17774%next\;
        \$16231%now\ <= \$16231%next\;
        \$v7015%now\ <= \$v7015%next\;
        \$16202_ofs%now\ <= \$16202_ofs%next\;
        \$v7091%now\ <= \$v7091%next\;
        \$16217_hd%now\ <= \$16217_hd%next\;
        \$v6400%now\ <= \$v6400%next\;
        \$v6388%now\ <= \$v6388%next\;
        \$16024%now\ <= \$16024%next\;
        \$12913%now\ <= \$12913%next\;
        \$17048_w16565937_arg%now\ <= \$17048_w16565937_arg%next\;
        \$15476_modulo6685895_id%now\ <= \$15476_modulo6685895_id%next\;
        \$16823_compbranch6505931_result%now\ <= \$16823_compbranch6505931_result%next\;
        \$16928_compbranch6505934_result%now\ <= \$16928_compbranch6505934_result%next\;
        \$18475%now\ <= \$18475%next\;
        \$17890%now\ <= \$17890%next\;
        \$15580_modulo6685896_id%now\ <= \$15580_modulo6685896_id%next\;
        \$15828_compare6445897_result%now\ <= \$15828_compare6445897_result%next\;
        \$12936%now\ <= \$12936%next\;
        \$17165%now\ <= \$17165%next\;
        \$12660%now\ <= \$12660%next\;
        \$v7232%now\ <= \$v7232%next\;
        \$12736%now\ <= \$12736%next\;
        \$v6724%now\ <= \$v6724%next\;
        \$18724_hd%now\ <= \$18724_hd%next\;
        \$17775%now\ <= \$17775%next\;
        \$16630%now\ <= \$16630%next\;
        \$15341_modulo6685888_id%now\ <= \$15341_modulo6685888_id%next\;
        \$18187%now\ <= \$18187%next\;
        \$v6998%now\ <= \$v6998%next\;
        \$17580_w%now\ <= \$17580_w%next\;
        \$17785%now\ <= \$17785%next\;
        \$12716%now\ <= \$12716%next\;
        \$15253_modulo6685896_id%now\ <= \$15253_modulo6685896_id%next\;
        \$14135%now\ <= \$14135%next\;
        \$15828_compare6445897_arg%now\ <= \$15828_compare6445897_arg%next\;
        \$13129%now\ <= \$13129%next\;
        \$18194%now\ <= \$18194%next\;
        \$18193%now\ <= \$18193%next\;
        \$16916_compare6445898_arg%now\ <= \$16916_compare6445898_arg%next\;
        \$17812%now\ <= \$17812%next\;
        \$12806_loop666_id%now\ <= \$12806_loop666_id%next\;
        \$15204_binop_int6435908_result%now\ <= \$15204_binop_int6435908_result%next\;
        \$v7210%now\ <= \$v7210%next\;
        \$17457_aux664_arg%now\ <= \$17457_aux664_arg%next\;
        \$14453_next_acc%now\ <= \$14453_next_acc%next\;
        \$18571%now\ <= \$18571%next\;
        \$15309_modulo6685895_result%now\ <= \$15309_modulo6685895_result%next\;
        \$17879_hd%now\ <= \$17879_hd%next\;
        \$13138_w%now\ <= \$13138_w%next\;
        \$v6624%now\ <= \$v6624%next\;
        \$v6992%now\ <= \$v6992%next\;
        \$14644_binop_int6435901_arg%now\ <= \$14644_binop_int6435901_arg%next\;
        \$v6515%now\ <= \$v6515%next\;
        \$13507%now\ <= \$13507%next\;
        \$19235%now\ <= \$19235%next\;
        \$17593%now\ <= \$17593%next\;
        \$17460_aux664_result%now\ <= \$17460_aux664_result%next\;
        \$v7283%now\ <= \$v7283%next\;
        \$16986_compare6445898_result%now\ <= \$16986_compare6445898_result%next\;
        \$14930_r%now\ <= \$14930_r%next\;
        \$v6898%now\ <= \$v6898%next\;
        \$v6003%now\ <= \$v6003%next\;
        \$17466%now\ <= \$17466%next\;
        \$v6579%now\ <= \$v6579%next\;
        \$v6121%now\ <= \$v6121%next\;
        \$14621_modulo6685888_result%now\ <= \$14621_modulo6685888_result%next\;
        \$13689%now\ <= \$13689%next\;
        \$14804_binop_int6435903_result%now\ <= \$14804_binop_int6435903_result%next\;
        \$12782%now\ <= \$12782%next\;
        \$18995%now\ <= \$18995%next\;
        \$v6110%now\ <= \$v6110%next\;
        \$v6179%now\ <= \$v6179%next\;
        \$18043%now\ <= \$18043%next\;
        \$19251_w%now\ <= \$19251_w%next\;
        \$14381%now\ <= \$14381%next\;
        \$v6066%now\ <= \$v6066%next\;
        \$12546_dur%now\ <= \$12546_dur%next\;
        \$v6911%now\ <= \$v6911%next\;
        \$v6207%now\ <= \$v6207%next\;
        \$15253_modulo6685896_result%now\ <= \$15253_modulo6685896_result%next\;
        \$17889%now\ <= \$17889%next\;
        \$14311%now\ <= \$14311%next\;
        \$v6971%now\ <= \$v6971%next\;
        \$v5999%now\ <= \$v5999%next\;
        \$12906%now\ <= \$12906%next\;
        \$v7206%now\ <= \$v7206%next\;
        \$14917_modulo6685888_id%now\ <= \$14917_modulo6685888_id%next\;
        \$18661%now\ <= \$18661%next\;
        \$17957_hd%now\ <= \$17957_hd%next\;
        \$12924_w%now\ <= \$12924_w%next\;
        \$v6546%now\ <= \$v6546%next\;
        \$18280%now\ <= \$18280%next\;
        \$13148%now\ <= \$13148%next\;
        \$v6232%now\ <= \$v6232%next\;
        \$18633_loop665_arg%now\ <= \$18633_loop665_arg%next\;
        \$14757_modulo6685888_result%now\ <= \$14757_modulo6685888_result%next\;
        \$13922_wait662_result%now\ <= \$13922_wait662_result%next\;
        \$v7364%now\ <= \$v7364%next\;
        \$15580_modulo6685896_result%now\ <= \$15580_modulo6685896_result%next\;
        \$15421_modulo6685888_id%now\ <= \$15421_modulo6685888_id%next\;
        \$14610_r%now\ <= \$14610_r%next\;
        \$16916_compare6445898_id%now\ <= \$16916_compare6445898_id%next\;
        \$12886%now\ <= \$12886%next\;
        \$16195_forever6705924_id%now\ <= \$16195_forever6705924_id%next\;
        \$v6670%now\ <= \$v6670%next\;
        \$13817%now\ <= \$13817%next\;
        \$v6817%now\ <= \$v6817%next\;
        \$14221%now\ <= \$14221%next\;
        \$v6062%now\ <= \$v6062%next\;
        \$17389%now\ <= \$17389%next\;
        \$v6563%now\ <= \$v6563%next\;
        \$v6080%now\ <= \$v6080%next\;
        \$v6799%now\ <= \$v6799%next\;
        \$v7092%now\ <= \$v7092%next\;
        \$14296%now\ <= \$14296%next\;
        \$17815%now\ <= \$17815%next\;
        \$v6463%now\ <= \$v6463%next\;
        \$13100%now\ <= \$13100%next\;
        \$v6097%now\ <= \$v6097%next\;
        \$v7203%now\ <= \$v7203%next\;
        \$13808_hd%now\ <= \$13808_hd%next\;
        \$13822%now\ <= \$13822%next\;
        \$16121_v%now\ <= \$16121_v%next\;
        \$v6403%now\ <= \$v6403%next\;
        \$17000_sp%now\ <= \$17000_sp%next\;
        \$12735%now\ <= \$12735%next\;
        \$v6424%now\ <= \$v6424%next\;
        \$15261_modulo6685888_result%now\ <= \$15261_modulo6685888_result%next\;
        \$17500%now\ <= \$17500%next\;
        \$17805%now\ <= \$17805%next\;
        \$v6421%now\ <= \$v6421%next\;
        \$13510%now\ <= \$13510%next\;
        \$13940%now\ <= \$13940%next\;
        \$v7433%now\ <= \$v7433%next\;
        \$15309_modulo6685895_arg%now\ <= \$15309_modulo6685895_arg%next\;
        \$18657%now\ <= \$18657%next\;
        \$16574_compare6445898_arg%now\ <= \$16574_compare6445898_arg%next\;
        \$13317%now\ <= \$13317%next\;
        \$v6287%now\ <= \$v6287%next\;
        \$12903%now\ <= \$12903%next\;
        \$16382%now\ <= \$16382%next\;
        \$15897%now\ <= \$15897%next\;
        \$14941_modulo6685888_result%now\ <= \$14941_modulo6685888_result%next\;
        \$14909_modulo6685895_result%now\ <= \$14909_modulo6685895_result%next\;
        \$v7135%now\ <= \$v7135%next\;
        \$18806%now\ <= \$18806%next\;
        \$17458_loop666_arg%now\ <= \$17458_loop666_arg%next\;
        \$12938%now\ <= \$12938%next\;
        \$15531_binop_int6435913_id%now\ <= \$15531_binop_int6435913_id%next\;
        \$15284_binop_int6435909_id%now\ <= \$15284_binop_int6435909_id%next\;
        \$13700%now\ <= \$13700%next\;
        \$18843%now\ <= \$18843%next\;
        \$15364_binop_int6435910_id%now\ <= \$15364_binop_int6435910_id%next\;
        \$12523_make_block579_arg%now\ <= \$12523_make_block579_arg%next\;
        \$v7245%now\ <= \$v7245%next\;
        \$16317%now\ <= \$16317%next\;
        \$18348%now\ <= \$18348%next\;
        \$13101%now\ <= \$13101%next\;
        \$v6069%now\ <= \$v6069%next\;
        \$16063_w6515922_result%now\ <= \$16063_w6515922_result%next\;
        \$v6096%now\ <= \$v6096%next\;
        \$12864_copy_root_in_ram6635886_arg%now\ <= \$12864_copy_root_in_ram6635886_arg%next\;
        \$14669_modulo6685895_arg%now\ <= \$14669_modulo6685895_arg%next\;
        \$17561%now\ <= \$17561%next\;
        \$19118%now\ <= \$19118%next\;
        \$14837_modulo6685888_id%now\ <= \$14837_modulo6685888_id%next\;
        \$12694%now\ <= \$12694%next\;
        \$15284_binop_int6435909_arg%now\ <= \$15284_binop_int6435909_arg%next\;
        \$12701%now\ <= \$12701%next\;
        \$v7450%now\ <= \$v7450%next\;
        \$16158_forever6705923_id%now\ <= \$16158_forever6705923_id%next\;
        \$15101_modulo6685888_id%now\ <= \$15101_modulo6685888_id%next\;
        \$v7145%now\ <= \$v7145%next\;
        \$v6654%now\ <= \$v6654%next\;
        \$v6042%now\ <= \$v6042%next\;
        \$13234%now\ <= \$13234%next\;
        \$v6717%now\ <= \$v6717%next\;
        \$15580_modulo6685896_arg%now\ <= \$15580_modulo6685896_arg%next\;
        \$15500_modulo6685896_result%now\ <= \$15500_modulo6685896_result%next\;
        \$15447_forever6705911_arg%now\ <= \$15447_forever6705911_arg%next\;
        \$18189%now\ <= \$18189%next\;
        \rdy6469%now\ <= \rdy6469%next\;
        \$17964%now\ <= \$17964%next\;
        \$18319%now\ <= \$18319%next\;
        \$v6920%now\ <= \$v6920%next\;
        \$v6989%now\ <= \$v6989%next\;
        \$14315_v%now\ <= \$14315_v%next\;
        \$18124%now\ <= \$18124%next\;
        \$16321%now\ <= \$16321%next\;
        \$v5986%now\ <= \$v5986%next\;
        \$13384%now\ <= \$13384%next\;
        \$13379_hd%now\ <= \$13379_hd%next\;
        \$15421_modulo6685888_arg%now\ <= \$15421_modulo6685888_arg%next\;
        \$v7365%now\ <= \$v7365%next\;
        \$13922_wait662_id%now\ <= \$13922_wait662_id%next\;
        \$12549%now\ <= \$12549%next\;
        \$v6832%now\ <= \$v6832%next\;
        \$v6765%now\ <= \$v6765%next\;
        \$v6104%now\ <= \$v6104%next\;
        \$18730%now\ <= \$18730%next\;
        \$18184%now\ <= \$18184%next\;
        \$17892%now\ <= \$17892%next\;
        \$v6543%now\ <= \$v6543%next\;
        \$v6585%now\ <= \$v6585%next\;
        \$17671%now\ <= \$17671%next\;
        \$v6106%now\ <= \$v6106%next\;
        \$12704%now\ <= \$12704%next\;
        \$v7399%now\ <= \$v7399%next\;
        \$v7110%now\ <= \$v7110%next\;
        \$18118%now\ <= \$18118%next\;
        \$13540%now\ <= \$13540%next\;
        \$v6862%now\ <= \$v6862%next\;
        \$15508_modulo6685888_result%now\ <= \$15508_modulo6685888_result%next\;
        \$v7100%now\ <= \$v7100%next\;
        \$17513_forever6705889_arg%now\ <= \$17513_forever6705889_arg%next\;
        \$v6835%now\ <= \$v6835%next\;
        \$16203%now\ <= \$16203%next\;
        \$15229_modulo6685895_result%now\ <= \$15229_modulo6685895_result%next\;
        \$15910%now\ <= \$15910%next\;
        \$17456_loop665_result%now\ <= \$17456_loop665_result%next\;
        \$v5995%now\ <= \$v5995%next\;
        \$13765%now\ <= \$13765%next\;
        \$12807_loop665_result%now\ <= \$12807_loop665_result%next\;
        \$v6373%now\ <= \$v6373%next\;
        \$v6171%now\ <= \$v6171%next\;
        \$18473%now\ <= \$18473%next\;
        \$v6758%now\ <= \$v6758%next\;
        \$v7332%now\ <= \$v7332%next\;
        \$v6646%now\ <= \$v6646%next\;
        \$v6692%now\ <= \$v6692%next\;
        \$v7188%now\ <= \$v7188%next\;
        \$16063_w6515922_id%now\ <= \$16063_w6515922_id%next\;
        \$v6562%now\ <= \$v6562%next\;
        \$v6743%now\ <= \$v6743%next\;
        \$v7426%now\ <= \$v7426%next\;
        \$13463%now\ <= \$13463%next\;
        \$18686_copy_root_in_ram6635880_id%now\ <= \$18686_copy_root_in_ram6635880_id%next\;
        \$v7378%now\ <= \$v7378%next\;
        \$v6742%now\ <= \$v6742%next\;
        \$14989_modulo6685895_result%now\ <= \$14989_modulo6685895_result%next\;
        \$v7375%now\ <= \$v7375%next\;
        \$15204_binop_int6435908_arg%now\ <= \$15204_binop_int6435908_arg%next\;
        \$18845%now\ <= \$18845%next\;
        \$14008%now\ <= \$14008%next\;
        \$v6328%now\ <= \$v6328%next\;
        \$v7355%now\ <= \$v7355%next\;
        \$v7044%now\ <= \$v7044%next\;
        \$v6319%now\ <= \$v6319%next\;
        \$15364_binop_int6435910_arg%now\ <= \$15364_binop_int6435910_arg%next\;
        \$v6965%now\ <= \$v6965%next\;
        \$12879%now\ <= \$12879%next\;
        \$15284_binop_int6435909_result%now\ <= \$15284_binop_int6435909_result%next\;
        \$12804_loop665_result%now\ <= \$12804_loop665_result%next\;
        \$18546%now\ <= \$18546%next\;
        \$v7020%now\ <= \$v7020%next\;
        \$15564_modulo6685888_result%now\ <= \$15564_modulo6685888_result%next\;
        \$v7081%now\ <= \$v7081%next\;
        \$v5872%now\ <= \$v5872%next\;
        \$v7393%now\ <= \$v7393%next\;
        \$14152%now\ <= \$14152%next\;
        \$v6766%now\ <= \$v6766%next\;
        \$18841%now\ <= \$18841%next\;
        \$15661_binop_compare6455917_result%now\ <= \$15661_binop_compare6455917_result%next\;
        \$13316%now\ <= \$13316%next\;
        \$13009_hd%now\ <= \$13009_hd%next\;
        \$14909_modulo6685895_arg%now\ <= \$14909_modulo6685895_arg%next\;
        \$12682_make_block579_result%now\ <= \$12682_make_block579_result%next\;
        \$18738%now\ <= \$18738%next\;
        \$16509%now\ <= \$16509%next\;
        \$12688%now\ <= \$12688%next\;
        \$15577_r%now\ <= \$15577_r%next\;
        \$v6093%now\ <= \$v6093%next\;
        \$v6109%now\ <= \$v6109%next\;
        \$15564_modulo6685888_arg%now\ <= \$15564_modulo6685888_arg%next\;
        \$16928_compbranch6505934_id%now\ <= \$16928_compbranch6505934_id%next\;
        \$14884_binop_int6435904_arg%now\ <= \$14884_binop_int6435904_arg%next\;
        \$v6553%now\ <= \$v6553%next\;
        \$14092%now\ <= \$14092%next\;
        \$v6535%now\ <= \$v6535%next\;
        \$18732%now\ <= \$18732%next\;
        \$17066%now\ <= \$17066%next\;
        \$15389_modulo6685895_id%now\ <= \$15389_modulo6685895_id%next\;
        \$v6660%now\ <= \$v6660%next\;
        \$17337%now\ <= \$17337%next\;
        \$18826_w%now\ <= \$18826_w%next\;
        \$v6036%now\ <= \$v6036%next\;
        \$17374_v%now\ <= \$17374_v%next\;
        \$17502%now\ <= \$17502%next\;
        \$12942%now\ <= \$12942%next\;
        \$14773_modulo6685896_id%now\ <= \$14773_modulo6685896_id%next\;
        \$14757_modulo6685888_id%now\ <= \$14757_modulo6685888_id%next\;
        \$18041%now\ <= \$18041%next\;
        \$v6547%now\ <= \$v6547%next\;
        \$v6184%now\ <= \$v6184%next\;
        \$12864_copy_root_in_ram6635886_id%now\ <= \$12864_copy_root_in_ram6635886_id%next\;
        \$18470%now\ <= \$18470%next\;
        \$12835%now\ <= \$12835%next\;
        \$15909%now\ <= \$15909%next\;
        \$v6902%now\ <= \$v6902%next\;
        \$17009_sp%now\ <= \$17009_sp%next\;
        \$18476%now\ <= \$18476%next\;
        \$16626%now\ <= \$16626%next\;
        \$17804%now\ <= \$17804%next\;
        \$18443%now\ <= \$18443%next\;
        \$14701_modulo6685888_result%now\ <= \$14701_modulo6685888_result%next\;
        \$v7167%now\ <= \$v7167%next\;
        \$14902_res%now\ <= \$14902_res%next\;
        \$12717%now\ <= \$12717%next\;
        \$v6908%now\ <= \$v6908%next\;
        \$13917%now\ <= \$13917%next\;
        \$16749_sp%now\ <= \$16749_sp%next\;
        \$v6155%now\ <= \$v6155%next\;
        \$17243%now\ <= \$17243%next\;
        \$v6442%now\ <= \$v6442%next\;
        \$13923_make_block579_result%now\ <= \$13923_make_block579_result%next\;
        \$v7445%now\ <= \$v7445%next\;
        \$v6354%now\ <= \$v6354%next\;
        \$14508_v%now\ <= \$14508_v%next\;
        \$15157_modulo6685888_arg%now\ <= \$15157_modulo6685888_arg%next\;
        \$19267%now\ <= \$19267%next\;
        \$16846_compare6445898_id%now\ <= \$16846_compare6445898_id%next\;
        \$15170_r%now\ <= \$15170_r%next\;
        \$v6616%now\ <= \$v6616%next\;
        \$13926_make_block_n646_id%now\ <= \$13926_make_block_n646_id%next\;
        \$18478%now\ <= \$18478%next\;
        \$16440%now\ <= \$16440%next\;
        \$15451_binop_int6435912_arg%now\ <= \$15451_binop_int6435912_arg%next\;
        \$15980_v%now\ <= \$15980_v%next\;
        \$v6623%now\ <= \$v6623%next\;
        \$14909_modulo6685895_id%now\ <= \$14909_modulo6685895_id%next\;
        \$12830%now\ <= \$12830%next\;
        \$13149%now\ <= \$13149%next\;
        \$17164%now\ <= \$17164%next\;
        \$14463_v%now\ <= \$14463_v%next\;
        \$13019%now\ <= \$13019%next\;
        \$15613%now\ <= \$15613%next\;
        \$17535%now\ <= \$17535%next\;
        \$13818%now\ <= \$13818%next\;
        \$v6521%now\ <= \$v6521%next\;
        \$16763_v%now\ <= \$16763_v%next\;
        \$18669%now\ <= \$18669%next\;
        \$18660%now\ <= \$18660%next\;
        \$v6137%now\ <= \$v6137%next\;
        \$v6790%now\ <= \$v6790%next\;
        \$v7117%now\ <= \$v7117%next\;
        \$v6223%now\ <= \$v6223%next\;
        \$13105_copy_root_in_ram6635884_arg%now\ <= \$13105_copy_root_in_ram6635884_arg%next\;
        \$v7387%now\ <= \$v7387%next\;
        \$17547_copy_root_in_ram6635891_id%now\ <= \$17547_copy_root_in_ram6635891_id%next\;
        \$15157_modulo6685888_id%now\ <= \$15157_modulo6685888_id%next\;
        \$18632_loop666_arg%now\ <= \$18632_loop666_arg%next\;
        \$17173%now\ <= \$17173%next\;
        \$15447_forever6705911_id%now\ <= \$15447_forever6705911_id%next\;
        \$15861_v%now\ <= \$15861_v%next\;
        \$13223_hd%now\ <= \$13223_hd%next\;
        \$13524_hd%now\ <= \$13524_hd%next\;
        \$16336%now\ <= \$16336%next\;
        \$v6899%now\ <= \$v6899%next\;
        \$v7156%now\ <= \$v7156%next\;
        \$15302_res%now\ <= \$15302_res%next\;
        \$19268%now\ <= \$19268%next\;
        \$18572%now\ <= \$18572%next\;
        \$v7459%now\ <= \$v7459%next\;
        \$v7229%now\ <= \$v7229%next\;
        \$17883%now\ <= \$17883%next\;
        \$18048%now\ <= \$18048%next\;
        \$13385%now\ <= \$13385%next\;
        \$17239_v%now\ <= \$17239_v%next\;
        \$14773_modulo6685896_result%now\ <= \$14773_modulo6685896_result%next\;
        \$17592%now\ <= \$17592%next\;
        \$13926_make_block_n646_result%now\ <= \$13926_make_block_n646_result%next\;
        \$17749%now\ <= \$17749%next\;
        \$18668%now\ <= \$18668%next\;
        \$v7093%now\ <= \$v7093%next\;
        \$v6176%now\ <= \$v6176%next\;
        \$12710%now\ <= \$12710%next\;
        \$18913%now\ <= \$18913%next\;
        \$v7107%now\ <= \$v7107%next\;
        \$v6075%now\ <= \$v6075%next\;
        \$v6031%now\ <= \$v6031%next\;
        \$14861_modulo6685888_arg%now\ <= \$14861_modulo6685888_arg%next\;
        \$v6352%now\ <= \$v6352%next\;
        \$13924_apply638_result%now\ <= \$13924_apply638_result%next\;
        \$15883%now\ <= \$15883%next\;
        \$v6684%now\ <= \$v6684%next\;
        \$13309%now\ <= \$13309%next\;
        \$12829%now\ <= \$12829%next\;
        \$14273%now\ <= \$14273%next\;
        \rdy6504%now\ <= \rdy6504%next\;
        \$v6938%now\ <= \$v6938%next\;
        \$17371_v%now\ <= \$17371_v%next\;
        \$v6880%now\ <= \$v6880%next\;
        \$v7011%now\ <= \$v7011%next\;
        \$17232%now\ <= \$17232%next\;
        \$12864_copy_root_in_ram6635886_result%now\ <= \$12864_copy_root_in_ram6635886_result%next\;
        \$v6829%now\ <= \$v6829%next\;
        \$v7056%now\ <= \$v7056%next\;
        \$14139%now\ <= \$14139%next\;
        \$v6379%now\ <= \$v6379%next\;
        \$17332_sp%now\ <= \$17332_sp%next\;
        \$17048_w16565937_result%now\ <= \$17048_w16565937_result%next\;
        \$19266%now\ <= \$19266%next\;
        \$15588_modulo6685888_result%now\ <= \$15588_modulo6685888_result%next\;
        \$v7260%now\ <= \$v7260%next\;
        \$14621_modulo6685888_arg%now\ <= \$14621_modulo6685888_arg%next\;
        \$13924_apply638_arg%now\ <= \$13924_apply638_arg%next\;
        \$v6643%now\ <= \$v6643%next\;
        \$v6152%now\ <= \$v6152%next\;
        \$18994%now\ <= \$18994%next\;
        \$15250_r%now\ <= \$15250_r%next\;
        \$15044_binop_int6435906_result%now\ <= \$15044_binop_int6435906_result%next\;
        \$16650_sp%now\ <= \$16650_sp%next\;
        \$v7350%now\ <= \$v7350%next\;
        \$18633_loop665_result%now\ <= \$18633_loop665_result%next\;
        \$12553%now\ <= \$12553%next\;
        \$18044%now\ <= \$18044%next\;
        \$12720%now\ <= \$12720%next\;
        \$17594%now\ <= \$17594%next\;
        \$v6190%now\ <= \$v6190%next\;
        \$v5964%now\ <= \$v5964%next\;
        \$13926_make_block_n646_arg%now\ <= \$13926_make_block_n646_arg%next\;
        \$15077_modulo6685888_id%now\ <= \$15077_modulo6685888_id%next\;
        \$v7021%now\ <= \$v7021%next\;
        \$17018_w36575938_result%now\ <= \$17018_w36575938_result%next\;
        \$v6180%now\ <= \$v6180%next\;
        \$v6889%now\ <= \$v6889%next\;
        \$15715_res%now\ <= \$15715_res%next\;
        \$16349_v%now\ <= \$16349_v%next\;
        \$14964_binop_int6435905_arg%now\ <= \$14964_binop_int6435905_arg%next\;
        \$18998%now\ <= \$18998%next\;
        \$13158%now\ <= \$13158%next\;
        \$v6283%now\ <= \$v6283%next\;
        \$17393%now\ <= \$17393%next\;
        \$v5948%now\ <= \$v5948%next\;
        \$13092%now\ <= \$13092%next\;
        \$v6714%now\ <= \$v6714%next\;
        \$v6325%now\ <= \$v6325%next\;
        \$14997_modulo6685888_result%now\ <= \$14997_modulo6685888_result%next\;
        \$v6550%now\ <= \$v6550%next\;
        \$v6236%now\ <= \$v6236%next\;
        \$12934%now\ <= \$12934%next\;
        \$v6588%now\ <= \$v6588%next\;
        \$v6256%now\ <= \$v6256%next\;
        \$17458_loop666_id%now\ <= \$17458_loop666_id%next\;
        \$17032%now\ <= \$17032%next\;
        \$12706%now\ <= \$12706%next\;
        \$16673_v%now\ <= \$16673_v%next\;
        \$13688%now\ <= \$13688%next\;
        \$v7427%now\ <= \$v7427%next\;
        \$17458_loop666_result%now\ <= \$17458_loop666_result%next\;
        \$12681_wait662_arg%now\ <= \$12681_wait662_arg%next\;
        \$18673%now\ <= \$18673%next\;
        \$17324%now\ <= \$17324%next\;
        \$14070_v%now\ <= \$14070_v%next\;
        \$12737%now\ <= \$12737%next\;
        \$19214%now\ <= \$19214%next\;
        \$15787_res%now\ <= \$15787_res%next\;
        \$14589_modulo6685895_arg%now\ <= \$14589_modulo6685895_arg%next\;
        \$v5967%now\ <= \$v5967%next\;
        \$17968%now\ <= \$17968%next\;
        \$14738_v%now\ <= \$14738_v%next\;
        \$v5998%now\ <= \$v5998%next\;
        \$18639%now\ <= \$18639%next\;
        \$13766%now\ <= \$13766%next\;
        \$15413_modulo6685896_arg%now\ <= \$15413_modulo6685896_arg%next\;
        \$15860%now\ <= \$15860%next\;
        \$v7010%now\ <= \$v7010%next\;
        \$18564%now\ <= \$18564%next\;
        \$v7449%now\ <= \$v7449%next\;
        \$v7046%now\ <= \$v7046%next\;
        \$17532%now\ <= \$17532%next\;
        \$v6243%now\ <= \$v6243%next\;
        \$19213%now\ <= \$19213%next\;
        \$13529%now\ <= \$13529%next\;
        \$v6493%now\ <= \$v6493%next\;
        \$15421_modulo6685888_result%now\ <= \$15421_modulo6685888_result%next\;
        \$18191%now\ <= \$18191%next\;
        \$14564_binop_int6435900_id%now\ <= \$14564_binop_int6435900_id%next\;
        \$12679_loop666_arg%now\ <= \$12679_loop666_arg%next\;
        \$14406_v%now\ <= \$14406_v%next\;
        \$15619%now\ <= \$15619%next\;
        \$v6917%now\ <= \$v6917%next\;
        \$16507%now\ <= \$16507%next\;
        \$v7116%now\ <= \$v7116%next\;
        \$v7273%now\ <= \$v7273%next\;
        \$14165%now\ <= \$14165%next\;
        \$13920_loop666_id%now\ <= \$13920_loop666_id%next\;
        \$15618%now\ <= \$15618%next\;
        \$16403%now\ <= \$16403%next\;
        \$17476%now\ <= \$17476%next\;
        \$13626%now\ <= \$13626%next\;
        \$17967%now\ <= \$17967%next\;
        \$12709%now\ <= \$12709%next\;
        \$v7213%now\ <= \$v7213%next\;
        \$14861_modulo6685888_id%now\ <= \$14861_modulo6685888_id%next\;
        \$v6844%now\ <= \$v6844%next\;
        \$12804_loop665_arg%now\ <= \$12804_loop665_arg%next\;
        \$14281%now\ <= \$14281%next\;
        \$16272%now\ <= \$16272%next\;
        \$17572%now\ <= \$17572%next\;
        \$12705%now\ <= \$12705%next\;
        \$12696%now\ <= \$12696%next\;
        \$13117%now\ <= \$13117%next\;
        \$13605%now\ <= \$13605%next\;
        \$16288%now\ <= \$16288%next\;
        \$12853_forever6705887_id%now\ <= \$12853_forever6705887_id%next\;
        \$17734_copy_root_in_ram6635892_result%now\ <= \$17734_copy_root_in_ram6635892_result%next\;
        \$17759%now\ <= \$17759%next\;
        \$v6247%now\ <= \$v6247%next\;
        \$16986_compare6445898_id%now\ <= \$16986_compare6445898_id%next\;
        \$17314%now\ <= \$17314%next\;
        \$v7197%now\ <= \$v7197%next\;
        \$12680_loop665_arg%now\ <= \$12680_loop665_arg%next\;
        \$18119%now\ <= \$18119%next\;
        \$v6072%now\ <= \$v6072%next\;
        \$12760%now\ <= \$12760%next\;
        \$12548_dis%now\ <= \$12548_dis%next\;
        \$15077_modulo6685888_arg%now\ <= \$15077_modulo6685888_arg%next\;
        \$14853_modulo6685896_result%now\ <= \$14853_modulo6685896_result%next\;
        \$18737%now\ <= \$18737%next\;
        \$18918%now\ <= \$18918%next\;
        \$17237_sp%now\ <= \$17237_sp%next\;
        \$15173_modulo6685896_arg%now\ <= \$15173_modulo6685896_arg%next\;
        \$17595%now\ <= \$17595%next\;
        \$17008%now\ <= \$17008%next\;
        \$17761_copy_root_in_ram6635891_arg%now\ <= \$17761_copy_root_in_ram6635891_arg%next\;
        \$v7101%now\ <= \$v7101%next\;
        \$12847%now\ <= \$12847%next\;
        \$v6859%now\ <= \$v6859%next\;
        \$12889%now\ <= \$12889%next\;
        \$18051%now\ <= \$18051%next\;
        \$v6219%now\ <= \$v6219%next\;
        \$14826_r%now\ <= \$14826_r%next\;
        \$14033%now\ <= \$14033%next\;
        \$v6606%now\ <= \$v6606%next\;
        \$18326%now\ <= \$18326%next\;
        \$18921%now\ <= \$18921%next\;
        \$13691%now\ <= \$13691%next\;
        \$v7083%now\ <= \$v7083%next\;
        \$v6956%now\ <= \$v6956%next\;
        \$15679_res%now\ <= \$15679_res%next\;
        \$v6666%now\ <= \$v6666%next\;
        \$19239%now\ <= \$19239%next\;
        \$14024%now\ <= \$14024%next\;
        \$v7442%now\ <= \$v7442%next\;
        \$16811_compare6445898_result%now\ <= \$16811_compare6445898_result%next\;
        \$14781_modulo6685888_arg%now\ <= \$14781_modulo6685888_arg%next\;
        \$v6335%now\ <= \$v6335%next\;
        \$19260%now\ <= \$19260%next\;
        \$17347%now\ <= \$17347%next\;
        \$15333_modulo6685896_id%now\ <= \$15333_modulo6685896_id%next\;
        \$18196%now\ <= \$18196%next\;
        \$v6752%now\ <= \$v6752%next\;
        \$16300%now\ <= \$16300%next\;
        \$17673%now\ <= \$17673%next\;
        \$13227%now\ <= \$13227%next\;
        \$16612_compare6445898_arg%now\ <= \$16612_compare6445898_arg%next\;
        \$13925_offsetclosure_n639_result%now\ <= \$13925_offsetclosure_n639_result%next\;
        \$v6409%now\ <= \$v6409%next\;
        \$17814%now\ <= \$17814%next\;
        \$17585_hd%now\ <= \$17585_hd%next\;
        \$17509_forever6705890_id%now\ <= \$17509_forever6705890_id%next\;
        \$17566%now\ <= \$17566%next\;
        \$12814%now\ <= \$12814%next\;
        \$19242%now\ <= \$19242%next\;
        \$17497%now\ <= \$17497%next\;
        \$13695%now\ <= \$13695%next\;
        \$v6394%now\ <= \$v6394%next\;
        \$v7397%now\ <= \$v7397%next\;
        \$v7289%now\ <= \$v7289%next\;
        \$v7194%now\ <= \$v7194%next\;
        \$17874_w%now\ <= \$17874_w%next\;
        \$18844%now\ <= \$18844%next\;
        \$15181_modulo6685888_arg%now\ <= \$15181_modulo6685888_arg%next\;
        \$18175_w%now\ <= \$18175_w%next\;
        \$v5876%now\ <= \$v5876%next\;
        \$18676%now\ <= \$18676%next\;
        \$17539%now\ <= \$17539%next\;
        \$v7115%now\ <= \$v7115%next\;
        \$v6263%now\ <= \$v6263%next\;
        \$v6353%now\ <= \$v6353%next\;
        \$18335_w%now\ <= \$18335_w%next\;
        \$18993%now\ <= \$18993%next\;
        \$13928_w652_id%now\ <= \$13928_w652_id%next\;
        \$17504%now\ <= \$17504%next\;
        \$18046%now\ <= \$18046%next\;
        \$12670%now\ <= \$12670%next\;
        \$v5972%now\ <= \$v5972%next\;
        \$v6133%now\ <= \$v6133%next\;
        \$12743%now\ <= \$12743%next\;
        \$13539%now\ <= \$13539%next\;
        \$v5947%now\ <= \$v5947%next\;
        \$17117_v%now\ <= \$17117_v%next\;
        \$15173_modulo6685896_result%now\ <= \$15173_modulo6685896_result%next\;
        \$15819_v%now\ <= \$15819_v%next\;
        \$17547_copy_root_in_ram6635891_arg%now\ <= \$17547_copy_root_in_ram6635891_arg%next\;
        \$12681_wait662_id%now\ <= \$12681_wait662_id%next\;
        \$14043_v%now\ <= \$14043_v%next\;
        \$13814%now\ <= \$13814%next\;
        \$12803_loop666_arg%now\ <= \$12803_loop666_arg%next\;
        \$v6436%now\ <= \$v6436%next\;
        \$19136%now\ <= \$19136%next\;
        \$18674%now\ <= \$18674%next\;
        \$v6784%now\ <= \$v6784%next\;
        \$v7296%now\ <= \$v7296%next\;
        \$17395%now\ <= \$17395%next\;
        \$13236%now\ <= \$13236%next\;
        \$13464%now\ <= \$13464%next\;
        \$14051%now\ <= \$14051%next\;
        \$v7014%now\ <= \$v7014%next\;
        \$17320%now\ <= \$17320%next\;
        \$v7095%now\ <= \$v7095%next\;
        \$v6433%now\ <= \$v6433%next\;
        \$12681_wait662_result%now\ <= \$12681_wait662_result%next\;
        \$13383%now\ <= \$13383%next\;
        \$14578_v%now\ <= \$14578_v%next\;
        \$v7112%now\ <= \$v7112%next\;
        \$17675%now\ <= \$17675%next\;
        \$19127_w%now\ <= \$19127_w%next\;
        \$18808%now\ <= \$18808%next\;
        \$14148%now\ <= \$14148%next\;
        \$18705%now\ <= \$18705%next\;
        \$14804_binop_int6435903_id%now\ <= \$14804_binop_int6435903_id%next\;
        \$v6650%now\ <= \$v6650%next\;
        \$v7267%now\ <= \$v7267%next\;
        \$13624%now\ <= \$13624%next\;
        \$15588_modulo6685888_arg%now\ <= \$15588_modulo6685888_arg%next\;
        \$v7051%now\ <= \$v7051%next\;
        \$v5867%now\ <= \$v5867%next\;
        \$17388%now\ <= \$17388%next\;
        \$15173_modulo6685896_id%now\ <= \$15173_modulo6685896_id%next\;
        \$16589_compbranch6505927_result%now\ <= \$16589_compbranch6505927_result%next\;
        \$14069%now\ <= \$14069%next\;
        \$v6531%now\ <= \$v6531%next\;
        \$12713%now\ <= \$12713%next\;
        \$13021%now\ <= \$13021%next\;
        \$18666_next%now\ <= \$18666_next%next\;
        \$14446_v%now\ <= \$14446_v%next\;
        \$17677%now\ <= \$17677%next\;
        \$18740%now\ <= \$18740%next\;
        \$18842%now\ <= \$18842%next\;
        \$17972%now\ <= \$17972%next\;
        \$14989_modulo6685895_id%now\ <= \$14989_modulo6685895_id%next\;
        \$17598%now\ <= \$17598%next\;
        \$12522_wait662_id%now\ <= \$12522_wait662_id%next\;
        \$18701%now\ <= \$18701%next\;
        \$16662_fill6535928_arg%now\ <= \$16662_fill6535928_arg%next\;
        \$17490_next%now\ <= \$17490_next%next\;
        \$v6759%now\ <= \$v6759%next\;
        \$16928_compbranch6505934_arg%now\ <= \$16928_compbranch6505934_arg%next\;
        \$18922%now\ <= \$18922%next\;
        \$18464_hd%now\ <= \$18464_hd%next\;
        \$16963_compbranch6505935_result%now\ <= \$16963_compbranch6505935_result%next\;
        \$13992_v%now\ <= \$13992_v%next\;
        \$15508_modulo6685888_arg%now\ <= \$15508_modulo6685888_arg%next\;
        \$12929_hd%now\ <= \$12929_hd%next\;
        \$v7457%now\ <= \$v7457%next\;
        \$13538%now\ <= \$13538%next\;
        \$16457%now\ <= \$16457%next\;
        \$15306_r%now\ <= \$15306_r%next\;
        \$v6705%now\ <= \$v6705%next\;
        \$18122%now\ <= \$18122%next\;
        \$v7102%now\ <= \$v7102%next\;
        \$19143%now\ <= \$19143%next\;
        \$18670_next%now\ <= \$18670_next%next\;
        \$18634_aux664_arg%now\ <= \$18634_aux664_arg%next\;
        \$18793_copy_root_in_ram6635879_id%now\ <= \$18793_copy_root_in_ram6635879_id%next\;
        \$15149_modulo6685895_id%now\ <= \$15149_modulo6685895_id%next\;
        \$16788_compbranch6505930_result%now\ <= \$16788_compbranch6505930_result%next\;
        \$13535%now\ <= \$13535%next\;
        \$15545_v%now\ <= \$15545_v%next\;
        \$17482%now\ <= \$17482%next\;
        \$v7061%now\ <= \$v7061%next\;
        \$v6253%now\ <= \$v6253%next\;
        \$13897%now\ <= \$13897%next\;
        \$18735%now\ <= \$18735%next\;
        \$v7126%now\ <= \$v7126%next\;
        \$18281%now\ <= \$18281%next\;
        \$16473%now\ <= \$16473%next\;
        \$14917_modulo6685888_result%now\ <= \$14917_modulo6685888_result%next\;
        \$16741%now\ <= \$16741%next\;
        \$16510_forever6705925_arg%now\ <= \$16510_forever6705925_arg%next\;
        \$v6536%now\ <= \$v6536%next\;
        \$12811%now\ <= \$12811%next\;
        \$v6796%now\ <= \$v6796%next\;
        \$18459_w%now\ <= \$18459_w%next\;
        \$14413_v%now\ <= \$14413_v%next\;
        \$12520_loop666_result%now\ <= \$12520_loop666_result%next\;
        \$16612_compare6445898_id%now\ <= \$16612_compare6445898_id%next\;
        \$17747%now\ <= \$17747%next\;
        \$v7104%now\ <= \$v7104%next\;
        \$13939%now\ <= \$13939%next\;
        \$15661_binop_compare6455917_id%now\ <= \$15661_binop_compare6455917_id%next\;
        \$17973%now\ <= \$17973%next\;
        \$12804_loop665_id%now\ <= \$12804_loop665_id%next\;
        \$17758%now\ <= \$17758%next\;
        \$12719%now\ <= \$12719%next\;
        \$15397_modulo6685888_id%now\ <= \$15397_modulo6685888_id%next\;
        \$17105_w06555936_arg%now\ <= \$17105_w06555936_arg%next\;
        \$12792%now\ <= \$12792%next\;
        \$16194%now\ <= \$16194%next\;
        \$v7176%now\ <= \$v7176%next\;
        \$14829_modulo6685895_arg%now\ <= \$14829_modulo6685895_arg%next\;
        \$18049%now\ <= \$18049%next\;
        \$13536%now\ <= \$13536%next\;
        \$12842%now\ <= \$12842%next\;
        \$v7182%now\ <= \$v7182%next\;
        \$v6511%now\ <= \$v6511%next\;
        \$14693_modulo6685896_id%now\ <= \$14693_modulo6685896_id%next\;
        \$13023%now\ <= \$13023%next\;
        \$v6098%now\ <= \$v6098%next\;
        \$15792_compare6445897_arg%now\ <= \$15792_compare6445897_arg%next\;
        \$v6905%now\ <= \$v6905%next\;
        \$13313%now\ <= \$13313%next\;
        \$14552%now\ <= \$14552%next\;
        \$16840_b%now\ <= \$16840_b%next\;
        \$16568_b%now\ <= \$16568_b%next\;
        \$14423_v%now\ <= \$14423_v%next\;
        \$v6527%now\ <= \$v6527%next\;
        \$18262%now\ <= \$18262%next\;
        \$13078_copy_root_in_ram6635885_result%now\ <= \$13078_copy_root_in_ram6635885_result%next\;
        \$18351%now\ <= \$18351%next\;
        \$16232%now\ <= \$16232%next\;
        \$16133%now\ <= \$16133%next\;
        \$15711_v%now\ <= \$15711_v%next\;
        \$15614_forever6705914_id%now\ <= \$15614_forever6705914_id%next\;
        \$13004_w%now\ <= \$13004_w%next\;
        \$12803_loop666_id%now\ <= \$12803_loop666_id%next\;
        \$12744%now\ <= \$12744%next\;
        \$13311%now\ <= \$13311%next\;
        \$18664_next%now\ <= \$18664_next%next\;
        \$19264%now\ <= \$19264%next\;
        \$13472_next%now\ <= \$13472_next%next\;
        \$16858_compbranch6505932_id%now\ <= \$16858_compbranch6505932_id%next\;
        \$v7096%now\ <= \$v7096%next\;
        \$17966%now\ <= \$17966%next\;
        \$v6787%now\ <= \$v6787%next\;
        \$17459_loop665_result%now\ <= \$17459_loop665_result%next\;
        \$v7120%now\ <= \$v7120%next\;
        \$17310%now\ <= \$17310%next\;
        \$17492_next%now\ <= \$17492_next%next\;
        \$v6045%now\ <= \$v6045%next\;
        \$17748%now\ <= \$17748%next\;
        \$18638%now\ <= \$18638%next\;
        \$15792_compare6445897_id%now\ <= \$15792_compare6445897_id%next\;
        \$13963%now\ <= \$13963%next\;
        \$v6140%now\ <= \$v6140%next\;
        \$12933%now\ <= \$12933%next\;
        \$18640%now\ <= \$18640%next\;
        \$13528%now\ <= \$13528%next\;
        \$v7254%now\ <= \$v7254%next\;
        \$16881_compare6445898_id%now\ <= \$16881_compare6445898_id%next\;
        \$17460_aux664_arg%now\ <= \$17460_aux664_arg%next\;
        \$12523_make_block579_result%now\ <= \$12523_make_block579_result%next\;
        \$13922_wait662_arg%now\ <= \$13922_wait662_arg%next\;
        \$v6156%now\ <= \$v6156%next\;
        \$v6814%now\ <= \$v6814%next\;
        \$v7419%now\ <= \$v7419%next\;
        \$15451_binop_int6435912_result%now\ <= \$15451_binop_int6435912_result%next\;
        \$v6322%now\ <= \$v6322%next\;
        \$17331_sp%now\ <= \$17331_sp%next\;
        \$17894%now\ <= \$17894%next\;
        \$v6002%now\ <= \$v6002%next\;
        \$v6476%now\ <= \$v6476%next\;
        \$13239%now\ <= \$13239%next\;
        \$12708%now\ <= \$12708%next\;
        \$18812%now\ <= \$18812%next\;
        \$v6187%now\ <= \$v6187%next\;
        \$v7072%now\ <= \$v7072%next\;
        \rdy6148%now\ <= \rdy6148%next\;
        \$18047%now\ <= \$18047%next\;
        \$14644_binop_int6435901_id%now\ <= \$14644_binop_int6435901_id%next\;
        \$14597_modulo6685888_id%now\ <= \$14597_modulo6685888_id%next\;
        \$v7103%now\ <= \$v7103%next\;
        \$19261%now\ <= \$19261%next\;
        \$16893_compbranch6505933_arg%now\ <= \$16893_compbranch6505933_arg%next\;
        \$13390%now\ <= \$13390%next\;
        \$16534%now\ <= \$16534%next\;
        \$v7191%now\ <= \$v7191%next\;
        \$19002%now\ <= \$19002%next\;
        \$v7041%now\ <= \$v7041%next\;
        \$v6968%now\ <= \$v6968%next\;
        \$v7127%now\ <= \$v7127%next\;
        \$17520_copy_root_in_ram6635893_result%now\ <= \$17520_copy_root_in_ram6635893_result%next\;
        \$v6332%now\ <= \$v6332%next\;
        \$13229%now\ <= \$13229%next\;
        \$v6159%now\ <= \$v6159%next\;
        \$15684_compare6445897_id%now\ <= \$15684_compare6445897_id%next\;
        \$v7114%now\ <= \$v7114%next\;
        \$17544%now\ <= \$17544%next\;
        \$v6704%now\ <= \$v6704%next\;
        \$18040%now\ <= \$18040%next\;
        \$17786%now\ <= \$17786%next\;
        \$v7233%now\ <= \$v7233%next\;
        \$14207_loop_push6495899_arg%now\ <= \$14207_loop_push6495899_arg%next\;
        \$16709%now\ <= \$16709%next\;
        \$v7113%now\ <= \$v7113%next\;
        \$14724_binop_int6435902_arg%now\ <= \$14724_binop_int6435902_arg%next\;
        \$13232%now\ <= \$13232%next\;
        \$16986_compare6445898_arg%now\ <= \$16986_compare6445898_arg%next\;
        \$v6054%now\ <= \$v6054%next\;
        \$16074_v%now\ <= \$16074_v%next\;
        \$v6781%now\ <= \$v6781%next\;
        \$v7047%now\ <= \$v7047%next\;
        \$17503%now\ <= \$17503%next\;
        \$13147%now\ <= \$13147%next\;
        \$v6259%now\ <= \$v6259%next\;
        \$v6144%now\ <= \$v6144%next\;
        \$13018%now\ <= \$13018%next\;
        \$v6603%now\ <= \$v6603%next\;
        \$14016_v%now\ <= \$14016_v%next\;
        \$16752_fill6545929_id%now\ <= \$16752_fill6545929_id%next\;
        \$v5973%now\ <= \$v5973%next\;
        \$13815%now\ <= \$13815%next\;
        \$v7033%now\ <= \$v7033%next\;
        \$v5983%now\ <= \$v5983%next\;
        \$19271%now\ <= \$19271%next\;
        \$v6735%now\ <= \$v6735%next\;
        \$v6769%now\ <= \$v6769%next\;
        \$v7242%now\ <= \$v7242%next\;
        \$16508%now\ <= \$16508%next\;
        \$12808_aux664_arg%now\ <= \$12808_aux664_arg%next\;
        \$18708%now\ <= \$18708%next\;
        \$18991%now\ <= \$18991%next\;
        \$14471%now\ <= \$14471%next\;
        \$v7070%now\ <= \$v7070%next\;
        \$12547%now\ <= \$12547%next\;
        \$v7031%now\ <= \$v7031%next\;
        \$v6315%now\ <= \$v6315%next\;
        \$12674%now\ <= \$12674%next\;
        \$12846%now\ <= \$12846%next\;
        \$17010%now\ <= \$17010%next\;
        \$17560%now\ <= \$17560%next\;
        \$16156%now\ <= \$16156%next\;
        \$15021_modulo6685888_id%now\ <= \$15021_modulo6685888_id%next\;
        \$13925_offsetclosure_n639_arg%now\ <= \$13925_offsetclosure_n639_arg%next\;
        \$14898_v%now\ <= \$14898_v%next\;
        \$14693_modulo6685896_result%now\ <= \$14693_modulo6685896_result%next\;
        \$15497_r%now\ <= \$15497_r%next\;
        \$13105_copy_root_in_ram6635884_id%now\ <= \$13105_copy_root_in_ram6635884_id%next\;
        \$17434%now\ <= \$17434%next\;
        \$16515%now\ <= \$16515%next\;
        \$14512_v%now\ <= \$14512_v%next\;
        \$14300_v%now\ <= \$14300_v%next\;
        \$18261%now\ <= \$18261%next\;
        \$17207_arg%now\ <= \$17207_arg%next\;
        \$13315%now\ <= \$13315%next\;
        \$18992%now\ <= \$18992%next\;
        \$18344%now\ <= \$18344%next\;
        \$17183%now\ <= \$17183%next\;
        \$v7032%now\ <= \$v7032%next\;
        \result6112%now\ <= \result6112%next\;
        \$v5960%now\ <= \$v5960%next\;
        \$v7084%now\ <= \$v7084%next\;
        \$v6639%now\ <= \$v6639%next\;
        \$v7060%now\ <= \$v7060%next\;
        \$18030_w%now\ <= \$18030_w%next\;
        \$18190%now\ <= \$18190%next\;
        \$16380_v%now\ <= \$16380_v%next\;
        \$v6295%now\ <= \$v6295%next\;
        \$18924%now\ <= \$18924%next\;
        \$12659%now\ <= \$12659%next\;
        \$v6111%now\ <= \$v6111%next\;
        \$v6011%now\ <= \$v6011%next\;
        \$12891_copy_root_in_ram6635884_result%now\ <= \$12891_copy_root_in_ram6635884_result%next\;
        \$18621%now\ <= \$18621%next\;
        \$14185_next_env%now\ <= \$14185_next_env%next\;
        \$17166%now\ <= \$17166%next\;
        \$v6059%now\ <= \$v6059%next\;
        \$12703%now\ <= \$12703%next\;
        \$v6358%now\ <= \$v6358%next\;
        \$12832%now\ <= \$12832%next\;
        \$15684_compare6445897_result%now\ <= \$15684_compare6445897_result%next\;
        \$v7111%now\ <= \$v7111%next\;
        \$17895%now\ <= \$17895%next\;
        \$13812%now\ <= \$13812%next\;
        \$18632_loop666_id%now\ <= \$18632_loop666_id%next\;
        \$17952_w%now\ <= \$17952_w%next\;
        \$13820%now\ <= \$13820%next\;
        \$13533%now\ <= \$13533%next\;
        \$15805_binop_compare6455921_result%now\ <= \$15805_binop_compare6455921_result%next\;
        \$15413_modulo6685896_id%now\ <= \$15413_modulo6685896_id%next\;
        \$13977_v%now\ <= \$13977_v%next\;
        \$v6294%now\ <= \$v6294%next\;
        \$12857_forever6705883_id%now\ <= \$12857_forever6705883_id%next\;
        \$v7438%now\ <= \$v7438%next\;
        \$v7082%now\ <= \$v7082%next\;
        \$v6415%now\ <= \$v6415%next\;
        \$v5982%now\ <= \$v5982%next\;
        \$19265%now\ <= \$19265%next\;
        \$17011%now\ <= \$17011%next\;
        \$v7012%now\ <= \$v7012%next\;
        \$17505_forever6705894_id%now\ <= \$17505_forever6705894_id%next\;
        \$v7282%now\ <= \$v7282%next\;
        \$12813%now\ <= \$12813%next\;
        \$17499%now\ <= \$17499%next\;
        \$v6457%now\ <= \$v6457%next\;
        \$13150%now\ <= \$13150%next\;
        \$17808%now\ <= \$17808%next\;
        \$v6820%now\ <= \$v6820%next\;
        \$17970%now\ <= \$17970%next\;
        \$12803_loop666_result%now\ <= \$12803_loop666_result%next\;
        \$v7276%now\ <= \$v7276%next\;
        \$14964_binop_int6435905_result%now\ <= \$14964_binop_int6435905_result%next\;
        \$v7134%now\ <= \$v7134%next\;
        \$17809%now\ <= \$17809%next\;
        \$16404%now\ <= \$16404%next\;
        \$v7157%now\ <= \$v7157%next\;
        \$17969%now\ <= \$17969%next\;
        \$v6280%now\ <= \$v6280%next\;
        \$12845%now\ <= \$12845%next\;
        \$v6361%now\ <= \$v6361%next\;
        \$12561%now\ <= \$12561%next\;
        \$17545%now\ <= \$17545%next\;
        \$18634_aux664_id%now\ <= \$18634_aux664_id%next\;
        \$15410_r%now\ <= \$15410_r%next\;
        \$v6582%now\ <= \$v6582%next\;
        \$v6600%now\ <= \$v6600%next\;
        \$15062_res%now\ <= \$15062_res%next\;
        \$v6264%now\ <= \$v6264%next\;
        \$14342%now\ <= \$14342%next\;
        \$v6691%now\ <= \$v6691%next\;
        \$12562%now\ <= \$12562%next\;
        \result5939%now\ <= \result5939%next\;
        \$12657%now\ <= \$12657%next\;
        \$v7130%now\ <= \$v7130%next\;
        \$16193%now\ <= \$16193%next\;
        \$16916_compare6445898_result%now\ <= \$16916_compare6445898_result%next\;
        \$18839%now\ <= \$18839%next\;
        \$13787%now\ <= \$13787%next\;
        \$v7303%now\ <= \$v7303%next\;
        \$19146%now\ <= \$19146%next\;
        \$15684_compare6445897_arg%now\ <= \$15684_compare6445897_arg%next\;
        \$15142_res%now\ <= \$15142_res%next\;
        \$12905%now\ <= \$12905%next\;
        \$v6267%now\ <= \$v6267%next\;
        \$18658%now\ <= \$18658%next\;
        \$13386%now\ <= \$13386%next\;
        \$17465%now\ <= \$17465%next\;
        \$v6477%now\ <= \$v6477%next\;
        \$13025%now\ <= \$13025%next\;
        \$18678%now\ <= \$18678%next\;
        \$16461%now\ <= \$16461%next\;
        \$v6774%now\ <= \$v6774%next\;
        \$18180_hd%now\ <= \$18180_hd%next\;
        \$v6811%now\ <= \$v6811%next\;
        \$13791%now\ <= \$13791%next\;
        \$14464_v%now\ <= \$14464_v%next\;
        \$15851_argument1%now\ <= \$15851_argument1%next\;
        \$13022%now\ <= \$13022%next\;
        \$15101_modulo6685888_arg%now\ <= \$15101_modulo6685888_arg%next\;
        \$13124%now\ <= \$13124%next\;
        \$v6762%now\ <= \$v6762%next\;
        \$v6720%now\ <= \$v6720%next\;
        \$v6528%now\ <= \$v6528%next\;
        \$v6083%now\ <= \$v6083%next\;
        \$16724%now\ <= \$16724%next\;
        \$v6524%now\ <= \$v6524%next\;
        \$v6448%now\ <= \$v6448%next\;
        \$17184%now\ <= \$17184%next\;
        \$13228%now\ <= \$13228%next\;
        \$19139%now\ <= \$19139%next\;
        \$v7036%now\ <= \$v7036%next\;
        \$v6755%now\ <= \$v6755%next\;
        \$17533%now\ <= \$17533%next\;
        \result5974%now\ <= \result5974%next\;
        \$v7037%now\ <= \$v7037%next\;
        \$18589%now\ <= \$18589%next\;
        \$14669_modulo6685895_result%now\ <= \$14669_modulo6685895_result%next\;
        \$13813%now\ <= \$13813%next\;
        \$17105_w06555936_result%now\ <= \$17105_w06555936_result%next\;
        \$13921_loop665_arg%now\ <= \$13921_loop665_arg%next\;
        \$17599%now\ <= \$17599%next\;
        \$13921_loop665_result%now\ <= \$13921_loop665_result%next\;
        \$v7401%now\ <= \$v7401%next\;
        \$v6980%now\ <= \$v6980%next\;
        \$16337%now\ <= \$16337%next\;
        \$17534%now\ <= \$17534%next\;
        \$12558%now\ <= \$12558%next\;
        \$v6926%now\ <= \$v6926%next\;
        \$16811_compare6445898_id%now\ <= \$16811_compare6445898_id%next\;
        \$v5989%now\ <= \$v5989%next\;
        \$14103%now\ <= \$14103%next\;
        \$15556_modulo6685895_arg%now\ <= \$15556_modulo6685895_arg%next\;
        \$19147%now\ <= \$19147%next\;
        \$16383%now\ <= \$16383%next\;
        \$v7149%now\ <= \$v7149%next\;
        \$13314%now\ <= \$13314%next\;
        \$15639_v%now\ <= \$15639_v%next\;
        \$16624_argument2%now\ <= \$16624_argument2%next\;
        \$15069_modulo6685895_result%now\ <= \$15069_modulo6685895_result%next\;
        \$16662_fill6535928_id%now\ <= \$16662_fill6535928_id%next\;
        \rdy6113%now\ <= \rdy6113%next\;
        \$17542%now\ <= \$17542%next\;
        \$v6345%now\ <= \$v6345%next\;
        \$v6194%now\ <= \$v6194%next\;
        \$v6571%now\ <= \$v6571%next\;
        \$15531_binop_int6435913_result%now\ <= \$15531_binop_int6435913_result%next\;
        \$v6439%now\ <= \$v6439%next\;
        \$v6079%now\ <= \$v6079%next\;
        \$15621_forever6705915_arg%now\ <= \$15621_forever6705915_arg%next\;
        \$17884%now\ <= \$17884%next\;
        \$v7097%now\ <= \$v7097%next\;
        \$13927_branch_if648_id%now\ <= \$13927_branch_if648_id%next\;
        \$14982_res%now\ <= \$14982_res%next\;
        \$18353%now\ <= \$18353%next\;
        \$v7347%now\ <= \$v7347%next\;
        \$16846_compare6445898_arg%now\ <= \$16846_compare6445898_arg%next\;
        \$v6895%now\ <= \$v6895%next\;
        \$16195_forever6705924_arg%now\ <= \$16195_forever6705924_arg%next\;
        \$17589%now\ <= \$17589%next\;
        \$13017%now\ <= \$13017%next\;
        \$15747_v%now\ <= \$15747_v%next\;
        \$16662_fill6535928_result%now\ <= \$16662_fill6535928_result%next\;
        \$18345%now\ <= \$18345%next\;
        \$v7122%now\ <= \$v7122%next\;
        \$17048_w16565937_id%now\ <= \$17048_w16565937_id%next\;
        \$18686_copy_root_in_ram6635880_result%now\ <= \$18686_copy_root_in_ram6635880_result%next\;
        \$15093_modulo6685896_id%now\ <= \$15093_modulo6685896_id%next\;
        \$18736%now\ <= \$18736%next\;
        \$18671%now\ <= \$18671%next\;
        \$15500_modulo6685896_id%now\ <= \$15500_modulo6685896_id%next\;
        \$v7226%now\ <= \$v7226%next\;
        \$17459_loop665_id%now\ <= \$17459_loop665_id%next\;
        \$15333_modulo6685896_arg%now\ <= \$15333_modulo6685896_arg%next\;
        \$17807%now\ <= \$17807%next\;
        \$v6220%now\ <= \$v6220%next\;
        \$13821%now\ <= \$13821%next\;
        \$18035_hd%now\ <= \$18035_hd%next\;
        \$v6290%now\ <= \$v6290%next\;
        \$17172%now\ <= \$17172%next\;
        \$13394%now\ <= \$13394%next\;
        \$19338%now\ <= \$19338%next\;
        \$17368_v%now\ <= \$17368_v%next\;
        \$v5871%now\ <= \$v5871%next\;
        \$13958%now\ <= \$13958%next\;
        \$12824%now\ <= \$12824%next\;
        \$17562%now\ <= \$17562%next\;
        \$16322%now\ <= \$16322%next\;
        \$v7105%now\ <= \$v7105%next\;
        \$13698%now\ <= \$13698%next\;
        \$17520_copy_root_in_ram6635893_arg%now\ <= \$17520_copy_root_in_ram6635893_arg%next\;
        \$15556_modulo6685895_id%now\ <= \$15556_modulo6685895_id%next\;
        \$13105_copy_root_in_ram6635884_result%now\ <= \$13105_copy_root_in_ram6635884_result%next\;
        \$12891_copy_root_in_ram6635884_id%now\ <= \$12891_copy_root_in_ram6635884_id%next\;
        \$12806_loop666_arg%now\ <= \$12806_loop666_arg%next\;
        \$v6566%now\ <= \$v6566%next\;
        \$15181_modulo6685888_id%now\ <= \$15181_modulo6685888_id%next\;
        \$v7080%now\ <= \$v7080%next\;
        \$v6675%now\ <= \$v6675%next\;
        \$v6576%now\ <= \$v6576%next\;
        \$16998_argument3%now\ <= \$16998_argument3%next\;
        \$v7423%now\ <= \$v7423%next\;
        \$18728%now\ <= \$18728%next\;
        \$16157%now\ <= \$16157%next\;
        \$13684_hd%now\ <= \$13684_hd%next\;
        \$19111%now\ <= \$19111%next\;
        \$v6647%now\ <= \$v6647%next\;
        \$13091%now\ <= \$13091%next\;
        \$13143_hd%now\ <= \$13143_hd%next\;
        \$18793_copy_root_in_ram6635879_result%now\ <= \$18793_copy_root_in_ram6635879_result%next\;
        \$15769_binop_compare6455920_result%now\ <= \$15769_binop_compare6455920_result%next\;
        \$16462%now\ <= \$16462%next\;
        \$14265%now\ <= \$14265%next\;
        \$12916%now\ <= \$12916%next\;
        \$v6244%now\ <= \$v6244%next\;
        \$12742%now\ <= \$12742%next\;
        \$13119%now\ <= \$13119%next\;
        \$13972_v%now\ <= \$13972_v%next\;
        \$14884_binop_int6435904_result%now\ <= \$14884_binop_int6435904_result%next\;
        \$13951%now\ <= \$13951%next\;
        \$v7024%now\ <= \$v7024%next\;
        \$13923_make_block579_arg%now\ <= \$13923_make_block579_arg%next\;
        \$15648_compare6445897_result%now\ <= \$15648_compare6445897_result%next\;
        \$17330_sp%now\ <= \$17330_sp%next\;
        \$v6620%now\ <= \$v6620%next\;
        \$17353%now\ <= \$17353%next\;
        \$v6983%now\ <= \$v6983%next\;
        \$v7257%now\ <= \$v7257%next\;
        \$v6663%now\ <= \$v6663%next\;
        \$13118%now\ <= \$13118%next\;
        \$v6032%now\ <= \$v6032%next\;
        \$18672%now\ <= \$18672%next\;
        \$19074%now\ <= \$19074%next\;
        \$15309_modulo6685895_id%now\ <= \$15309_modulo6685895_id%next\;
        \$v6260%now\ <= \$v6260%next\;
        \$19076%now\ <= \$19076%next\;
        \rdy5975%now\ <= \rdy5975%next\;
        \$15124_binop_int6435907_result%now\ <= \$15124_binop_int6435907_result%next\;
        \$16334_v%now\ <= \$16334_v%next\;
        \$v7270%now\ <= \$v7270%next\;
        \$18042%now\ <= \$18042%next\;
        \$18611%now\ <= \$18611%next\;
        \$14377_v%now\ <= \$14377_v%next\;
        \$16381_v%now\ <= \$16381_v%next\;
        \$v6076%now\ <= \$v6076%next\;
        \$15908%now\ <= \$15908%next\;
        \$12563%now\ <= \$12563%next\;
        \$v7026%now\ <= \$v7026%next\;
        \$v6698%now\ <= \$v6698%next\;
        \$15013_modulo6685896_result%now\ <= \$15013_modulo6685896_result%next\;
        \$12805_aux664_arg%now\ <= \$12805_aux664_arg%next\;
        \$v7075%now\ <= \$v7075%next\;
        \$13024%now\ <= \$13024%next\;
        \$13965%now\ <= \$13965%next\;
        \$18573%now\ <= \$18573%next\;
        \$v6124%now\ <= \$v6124%next\;
        \$17481%now\ <= \$17481%next\;
        \$v6215%now\ <= \$v6215%next\;
        \$15720_compare6445897_result%now\ <= \$15720_compare6445897_result%next\;
        \$v7160%now\ <= \$v7160%next\;
        \$v6497%now\ <= \$v6497%next\;
        \$15044_binop_int6435906_arg%now\ <= \$15044_binop_int6435906_arg%next\;
        \$13097%now\ <= \$13097%next\;
        \$17456_loop665_arg%now\ <= \$17456_loop665_arg%next\;
        \$13952%now\ <= \$13952%next\;
        \$15093_modulo6685896_result%now\ <= \$15093_modulo6685896_result%next\;
        \$13924_apply638_id%now\ <= \$13924_apply638_id%next\;
        \$v6556%now\ <= \$v6556%next\;
        \$14701_modulo6685888_id%now\ <= \$14701_modulo6685888_id%next\;
        \$12687%now\ <= \$12687%next\;
        \$15473_r%now\ <= \$15473_r%next\;
        \$17061%now\ <= \$17061%next\;
        \$16725%now\ <= \$16725%next\;
        \$v6412%now\ <= \$v6412%next\;
        \$v7407%now\ <= \$v7407%next\;
        \$v6747%now\ <= \$v6747%next\;
        \$12831%now\ <= \$12831%next\;
        \$16651%now\ <= \$16651%next\;
        \$14781_modulo6685888_id%now\ <= \$14781_modulo6685888_id%next\;
        \$16658%now\ <= \$16658%next\;
        \$v7136%now\ <= \$v7136%next\;
        \$14589_modulo6685895_id%now\ <= \$14589_modulo6685895_id%next\;
        \$v5968%now\ <= \$v5968%next\;
        \$v6339%now\ <= \$v6339%next\;
        \$16788_compbranch6505930_id%now\ <= \$16788_compbranch6505930_id%next\;
        \$17486%now\ <= \$17486%next\;
        \$v6331%now\ <= \$v6331%next\;
        \$18553%now\ <= \$18553%next\;
        \$14034_v%now\ <= \$14034_v%next\;
        \$v7410%now\ <= \$v7410%next\;
        \$v7131%now\ <= \$v7131%next\;
        \$18284%now\ <= \$18284%next\;
        \$v7390%now\ <= \$v7390%next\;
        \$13306%now\ <= \$13306%next\;
        \$v6539%now\ <= \$v6539%next\;
        \$v7341%now\ <= \$v7341%next\;
        \$15090_r%now\ <= \$15090_r%next\;
        \$14906_r%now\ <= \$14906_r%next\;
        \$13462%now\ <= \$13462%next\;
        \$19270%now\ <= \$19270%next\;
        \$v6850%now\ <= \$v6850%next\;
        \$v7430%now\ <= \$v7430%next\;
        \$v6671%now\ <= \$v6671%next\;
        \$15149_modulo6685895_result%now\ <= \$15149_modulo6685895_result%next\;
        \$15756_compare6445897_id%now\ <= \$15756_compare6445897_id%next\;
        \$v6418%now\ <= \$v6418%next\;
        \$v6250%now\ <= \$v6250%next\;
        \$v6051%now\ <= \$v6051%next\;
        \$15621_forever6705915_id%now\ <= \$15621_forever6705915_id%next\;
        \$v6886%now\ <= \$v6886%next\;
        \$16858_compbranch6505932_result%now\ <= \$16858_compbranch6505932_result%next\;
        \$15222_res%now\ <= \$15222_res%next\;
        \$v6770%now\ <= \$v6770%next\;
        \$v7040%now\ <= \$v7040%next\;
        \$16301%now\ <= \$16301%next\;
        \$13911%now\ <= \$13911%next\;
        \$17680%now\ <= \$17680%next\;
        \$v6191%now\ <= \$v6191%next\;
        \$15138_v%now\ <= \$15138_v%next\;
        \$v6486%now\ <= \$v6486%next\;
        \$13152%now\ <= \$13152%next\;
        \$16155%now\ <= \$16155%next\;
        \$14933_modulo6685896_arg%now\ <= \$14933_modulo6685896_arg%next\;
        \$12693%now\ <= \$12693%next\;
        \$v7106%now\ <= \$v7106%next\;
        \$v7067%now\ <= \$v7067%next\;
        \$13920_loop666_result%now\ <= \$13920_loop666_result%next\;
        \$16293%now\ <= \$16293%next\;
        \$13159%now\ <= \$13159%next\;
        \$13953%now\ <= \$13953%next\;
        \$15625_binop_compare6455916_arg%now\ <= \$15625_binop_compare6455916_arg%next\;
        \$13015%now\ <= \$13015%next\;
        \$17799_hd%now\ <= \$17799_hd%next\;
        \$v6039%now\ <= \$v6039%next\;
        \$15611%now\ <= \$15611%next\;
        \$v6808%now\ <= \$v6808%next\;
        \$17444%now\ <= \$17444%next\;
        \$14853_modulo6685896_id%now\ <= \$14853_modulo6685896_id%next\;
        \$18665%now\ <= \$18665%next\;
        \$19132_hd%now\ <= \$19132_hd%next\;
        \$16313_v%now\ <= \$16313_v%next\;
        \$14757_modulo6685888_arg%now\ <= \$14757_modulo6685888_arg%next\;
        \$18710%now\ <= \$18710%next\;
        \$v5979%now\ <= \$v5979%next\;
        \$v6006%now\ <= \$v6006%next\;
        \$14621_modulo6685888_id%now\ <= \$14621_modulo6685888_id%next\;
        \$14941_modulo6685888_id%now\ <= \$14941_modulo6685888_id%next\;
        \$19073%now\ <= \$19073%next\;
        \$15733_binop_compare6455919_id%now\ <= \$15733_binop_compare6455919_id%next\;
        \$15620%now\ <= \$15620%next\;
        \$17596%now\ <= \$17596%next\;
        \$16413%now\ <= \$16413%next\;
        \$19141%now\ <= \$19141%next\;
        \$17753%now\ <= \$17753%next\;
        \$16706%now\ <= \$16706%next\;
        \$16296%now\ <= \$16296%next\;
        \$v7001%now\ <= \$v7001%next\;
        \$18468%now\ <= \$18468%next\;
        \$19000%now\ <= \$19000%next\;
        \$v5877%now\ <= \$v5877%next\;
        \$16951_compare6445898_id%now\ <= \$16951_compare6445898_id%next\;
        \$13231%now\ <= \$13231%next\;
        \$v6024%now\ <= \$v6024%next\;
        \$13130%now\ <= \$13130%next\;
        \$15469_res%now\ <= \$15469_res%next\;
        \$18471%now\ <= \$18471%next\;
        \$v6793%now\ <= \$v6793%next\;
        \$v7266%now\ <= \$v7266%next\;
        \$18350%now\ <= \$18350%next\;
        \$16357%now\ <= \$16357%next\;
        \$15149_modulo6685895_arg%now\ <= \$15149_modulo6685895_arg%next\;
        \$13987_v%now\ <= \$13987_v%next\;
        \$v7055%now\ <= \$v7055%next\;
        \$17483%now\ <= \$17483%next\;
        \$14260%now\ <= \$14260%next\;
        \$15588_modulo6685888_id%now\ <= \$15588_modulo6685888_id%next\;
        \$v7309%now\ <= \$v7309%next\;
        \$15643_res%now\ <= \$15643_res%next\;
        \$13078_copy_root_in_ram6635885_arg%now\ <= \$13078_copy_root_in_ram6635885_arg%next\;
        \$18914%now\ <= \$18914%next\;
        \$17660_w%now\ <= \$17660_w%next\;
        \$16846_compare6445898_result%now\ <= \$16846_compare6445898_result%next\;
        \$18817%now\ <= \$18817%next\;
        \$v6871%now\ <= \$v6871%next\;
        \$17672%now\ <= \$17672%next\;
        \$19148%now\ <= \$19148%next\;
        \$v7329%now\ <= \$v7329%next\;
        \$19072%now\ <= \$19072%next\;
        \$15733_binop_compare6455919_result%now\ <= \$15733_binop_compare6455919_result%next\;
        \$14081%now\ <= \$14081%next\;
        \$18545%now\ <= \$18545%next\;
        \$13889%now\ <= \$13889%next\;
        \$14015%now\ <= \$14015%next\;
        \$12840_next%now\ <= \$12840_next%next\;
        \$18686_copy_root_in_ram6635880_arg%now\ <= \$18686_copy_root_in_ram6635880_arg%next\;
        \$14742_res%now\ <= \$14742_res%next\;
        \$14586_r%now\ <= \$14586_r%next\;
        \$18195%now\ <= \$18195%next\;
        \$v6540%now\ <= \$v6540%next\;
        \$18793_copy_root_in_ram6635879_arg%now\ <= \$18793_copy_root_in_ram6635879_arg%next\;
        \$15317_modulo6685888_id%now\ <= \$15317_modulo6685888_id%next\;
        \$16551_compbranch6505926_result%now\ <= \$16551_compbranch6505926_result%next\;
        \$17811%now\ <= \$17811%next\;
        \$16980_b%now\ <= \$16980_b%next\;
        \$18349%now\ <= \$18349%next\;
        \$15451_binop_int6435912_id%now\ <= \$15451_binop_int6435912_id%next\;
        \$14002_v%now\ <= \$14002_v%next\;
        \$14997_modulo6685888_arg%now\ <= \$14997_modulo6685888_arg%next\;
        \$16335_v%now\ <= \$16335_v%next\;
        \$13014%now\ <= \$13014%next\;
        \$v6977%now\ <= \$v6977%next\;
        \$18039%now\ <= \$18039%next\;
        \$13448%now\ <= \$13448%next\;
        \$17571%now\ <= \$17571%next\;
        \$17757%now\ <= \$17757%next\;
        \$v6018%now\ <= \$v6018%next\;
        \$16358%now\ <= \$16358%next\;
        \$v7052%now\ <= \$v7052%next\;
        \$17352%now\ <= \$17352%next\;
        \$17756%now\ <= \$17756%next\;
        \$v6141%now\ <= \$v6141%next\;
        \$13391%now\ <= \$13391%next\;
        \$v6086%now\ <= \$v6086%next\;
        \$v6145%now\ <= \$v6145%next\;
        \$15066_r%now\ <= \$15066_r%next\;
        \result6147%now\ <= \result6147%next\;
        \$15446%now\ <= \$15446%next\;
        \$v6877%now\ <= \$v6877%next\;
        \$16041_v%now\ <= \$16041_v%next\;
        \$16063_w6515922_arg%now\ <= \$16063_w6515922_arg%next\;
        \$12700%now\ <= \$12700%next\;
        \$16951_compare6445898_result%now\ <= \$16951_compare6445898_result%next\;
        \$v6210%now\ <= \$v6210%next\;
        \$15564_modulo6685888_id%now\ <= \$15564_modulo6685888_id%next\;
        \$12721%now\ <= \$12721%next\;
        \$18920%now\ <= \$18920%next\;
        \$14393_hd%now\ <= \$14393_hd%next\;
        \$18282%now\ <= \$18282%next\;
        \$v7141%now\ <= \$v7141%next\;
        \$15157_modulo6685888_result%now\ <= \$15157_modulo6685888_result%next\;
        \$14850_r%now\ <= \$14850_r%next\;
        \$17601%now\ <= \$17601%next\;
        \$v6310%now\ <= \$v6310%next\;
        \$14493_v%now\ <= \$14493_v%next\;
        \$12711%now\ <= \$12711%next\;
        \$v5864%now\ <= \$v5864%next\;
        \$v6483%now\ <= \$v6483%next\;
        \$13819%now\ <= \$13819%next\;
        \$v7325%now\ <= \$v7325%next\;
        \$13120%now\ <= \$13120%next\;
        \$v7087%now\ <= \$v7087%next\;
        \$v6615%now\ <= \$v6615%next\;
        \$15146_r%now\ <= \$15146_r%next\;
        \$v7394%now\ <= \$v7394%next\;
        \$18347%now\ <= \$18347%next\;
        \$18700%now\ <= \$18700%next\;
        \$v6777%now\ <= \$v6777%next\;
        \$12940%now\ <= \$12940%next\;
        \$v7173%now\ <= \$v7173%next\;
        \$17062%now\ <= \$17062%next\;
        \$v7073%now\ <= \$v7073%next\;
        \$14025_v%now\ <= \$14025_v%next\;
        \$14561%now\ <= \$14561%next\;
        \$16437_v%now\ <= \$16437_v%next\;
        \$15549_res%now\ <= \$15549_res%next\;
        \$15253_modulo6685896_arg%now\ <= \$15253_modulo6685896_arg%next\;
        \$15013_modulo6685896_arg%now\ <= \$15013_modulo6685896_arg%next\;
        \$14822_res%now\ <= \$14822_res%next\;
        \$18847%now\ <= \$18847%next\;
        \$18840%now\ <= \$18840%next\;
        \$18340_hd%now\ <= \$18340_hd%next\;
        \$v7148%now\ <= \$v7148%next\;
        \$14884_binop_int6435904_id%now\ <= \$14884_binop_int6435904_id%next\;
        \$18632_loop666_result%now\ <= \$18632_loop666_result%next\;
        \$15226_r%now\ <= \$15226_r%next\;
        \$18422%now\ <= \$18422%next\;
        \$15444%now\ <= \$15444%next\;
        \$19137%now\ <= \$19137%next\;
        \$18923%now\ <= \$18923%next\;
        \$17161%now\ <= \$17161%next\;
        \$12662%now\ <= \$12662%next\;
        \$v7065%now\ <= \$v7065%next\;
        \$14662_res%now\ <= \$14662_res%next\;
        \$v6226%now\ <= \$v6226%next\;
        \$v7319%now\ <= \$v7319%next\;
        \$17396%now\ <= \$17396%next\;
        \$17806%now\ <= \$17806%next\;
        \$v6612%now\ <= \$v6612%next\;
        \$15805_binop_compare6455921_id%now\ <= \$15805_binop_compare6455921_id%next\;
        \$13305%now\ <= \$13305%next\;
        \$13230%now\ <= \$13230%next\;
        \$19056%now\ <= \$19056%next\;
        \$18469%now\ <= \$18469%next\;
        \$v7286%now\ <= \$v7286%next\;
        \$13534%now\ <= \$13534%next\;
        \$v7152%now\ <= \$v7152%next\;
        \$v6929%now\ <= \$v6929%next\;
        \$16910_b%now\ <= \$16910_b%next\;
        \$v7043%now\ <= \$v7043%next\;
        \$12850%now\ <= \$12850%next\;
        \$17456_loop665_id%now\ <= \$17456_loop665_id%next\;
        \$18477%now\ <= \$18477%next\;
        \$v7225%now\ <= \$v7225%next\;
        \$v6923%now\ <= \$v6923%next\;
        \$v6674%now\ <= \$v6674%next\;
        \$13699%now\ <= \$13699%next\;
        \$v6944%now\ <= \$v6944%next\;
        \$13923_make_block579_id%now\ <= \$13923_make_block579_id%next\;
        \$14207_loop_push6495899_id%now\ <= \$14207_loop_push6495899_id%next\;
        \$15648_compare6445897_arg%now\ <= \$15648_compare6445897_arg%next\;
        \$13803_w%now\ <= \$13803_w%next\;
        \$17780%now\ <= \$17780%next\;
        \$12876%now\ <= \$12876%next\;
        \$18656%now\ <= \$18656%next\;
        \$v6687%now\ <= \$v6687%next\;
        \$v6107%now\ <= \$v6107%next\;
        \$12661%now\ <= \$12661%next\;
        \$v6630%now\ <= \$v6630%next\;
        \$15697_binop_compare6455918_id%now\ <= \$15697_binop_compare6455918_id%next\;
        \$v7124%now\ <= \$v7124%next\;
        \$v7384%now\ <= \$v7384%next\;
        \$v7063%now\ <= \$v7063%next\;
        \$13928_w652_arg%now\ <= \$13928_w652_arg%next\;
        \$15465_v%now\ <= \$15465_v%next\;
        \$13622%now\ <= \$13622%next\;
        \$14355%now\ <= \$14355%next\;
        \$v7312%now\ <= \$v7312%next\;
        \$v6636%now\ <= \$v6636%next\;
        \$14770_r%now\ <= \$14770_r%next\;
        \$v6063%now\ <= \$v6063%next\;
        \$15013_modulo6685896_id%now\ <= \$15013_modulo6685896_id%next\;
        \$14690_r%now\ <= \$14690_r%next\;
        \$12807_loop665_arg%now\ <= \$12807_loop665_arg%next\;
        \$v6120%now\ <= \$v6120%next\;
        \$17810%now\ <= \$17810%next\;
        \$v6168%now\ <= \$v6168%next\;
        \$v7053%now\ <= \$v7053%next\;
        \$v7239%now\ <= \$v7239%next\;
        \$17236%now\ <= \$17236%next\;
        \$v7209%now\ <= \$v7209%next\;
        \$13128%now\ <= \$13128%next\;
        \$15229_modulo6685895_id%now\ <= \$15229_modulo6685895_id%next\;
        \$v7316%now\ <= \$v7316%next\;
        \$12690%now\ <= \$12690%next\;
        \$13925_offsetclosure_n639_id%now\ <= \$13925_offsetclosure_n639_id%next\;
        \$13020%now\ <= \$13020%next\;
        \$v6932%now\ <= \$v6932%next\;
        \$12539%now\ <= \$12539%next\;
        \$v6592%now\ <= \$v6592%next\;
        \$v6010%now\ <= \$v6010%next\;
        \$13093%now\ <= \$13093%next\;
        \$18323%now\ <= \$18323%next\;
        \$17965%now\ <= \$17965%next\;
        \$v5971%now\ <= \$v5971%next\;
        \$16659_sp%now\ <= \$16659_sp%next\;
        \$17547_copy_root_in_ram6635891_result%now\ <= \$17547_copy_root_in_ram6635891_result%next\;
        \$13690%now\ <= \$13690%next\;
        \$13628%now\ <= \$13628%next\;
        \$v6349%now\ <= \$v6349%next\;
        \$13465%now\ <= \$13465%next\;
        \$12812%now\ <= \$12812%next\;
        \$v6028%now\ <= \$v6028%next\;
        \$13374_w%now\ <= \$13374_w%next\;
        \$14368%now\ <= \$14368%next\;
        \$12718%now\ <= \$12718%next\;
        \$17784%now\ <= \$17784%next\;
        \$15508_modulo6685888_id%now\ <= \$15508_modulo6685888_id%next\;
        \$15364_binop_int6435910_result%now\ <= \$15364_binop_int6435910_result%next\;
        \$14613_modulo6685896_arg%now\ <= \$14613_modulo6685896_arg%next\;
        \$15751_res%now\ <= \$15751_res%next\;
        \$13537%now\ <= \$13537%next\;
        \$12654%now\ <= \$12654%next\;
        \$v7071%now\ <= \$v7071%next\;
        \$v6311%now\ <= \$v6311%next\;
        \$ram_lock%now\ <= \$ram_lock%next\;
        \$global_end_lock%now\ <= \$global_end_lock%next\;
        \$code_lock%now\ <= \$code_lock%next\;
        \state_var7464%now\ <= \state_var7464%next\;
        \state_var7463%now\ <= \state_var7463%next\;
        \state_var7462%now\ <= \state_var7462%next\;
        \state_var7461%now\ <= \state_var7461%next\;
        \state_var7460%now\ <= \state_var7460%next\;
        \state%now\ <= \state%next\;
      end if;
    end process;
      
      process(argument,\state%now\, clk,\state_var7464%now\,\state_var7463%now\,\state_var7462%now\,\state_var7461%now\,\state_var7460%now\, \$ram_value\, \$global_end_value\, \$code_value\, \$12559%now\, \$14060%now\, \$v6454%now\, \$14516_v%now\, \$15069_modulo6685895_arg%now\, \$18421%now\, \$v6570%now\, \$14564_binop_int6435900_arg%now\, \$17813%now\, \$v6841%now\, \$14666_r%now\, \$v7022%now\, \$14589_modulo6685895_result%now\, \$13392%now\, \$18996%now\, \$12673_rdy%now\, \$v6130%now\, \$v7263%now\, \$14917_modulo6685888_arg%now\, \$v6197%now\, \$19272%now\, \$v7123%now\, \$v6642%now\, \$18729%now\, \$18192%now\, \$13670%now\, \$v6127%now\, \$15675_v%now\, \$15077_modulo6685888_result%now\, \$v6725%now\, \$16182%now\, \$14052_v%now\, \$18354%now\, \$14749_modulo6685895_result%now\, \$v6451%now\, \$12545_x%now\, \$v7062%now\, \$17496_next%now\, \$12852%now\, \$13503%now\, \$v6473%now\, \$15531_binop_int6435913_arg%now\, \$17887%now\, \$18997%now\, \$18835%now\, \$v6567%now\, \$v7313%now\, \$14724_binop_int6435902_result%now\, \$12699%now\, \$v7125%now\, \$14989_modulo6685895_arg%now\, \$13090%now\, \$19003%now\, \$12522_wait662_arg%now\, \$16811_compare6445898_arg%now\, \$17893%now\, \$15661_binop_compare6455917_arg%now\, \$14126%now\, \$v7437%now\, \$17570%now\, \$16453_v%now\, \$17676%now\, \$18121%now\, \$v7222%now\, \$v6512%now\, \$13308%now\, \$17018_w36575938_arg%now\, \$v6206%now\, \$15484_modulo6685888_result%now\, \$v7170%now\, \$15614_forever6705914_arg%now\, \$16858_compbranch6505932_arg%now\, \$v7236%now\, \$v7153%now\, \$16893_compbranch6505933_id%now\, \$14597_modulo6685888_arg%now\, \$16141%now\, \$v6105%now\, \$v7446%now\, \$13156%now\, \$v6575%now\, \$19138%now\, \$16178_v%now\, \$13945%now\, \$v7094%now\, \$v6391%now\, \$18838%now\, \$13824%now\, \$v6959%now\, \$13531%now\, \$16788_compbranch6505930_arg%now\, \$17971%now\, \$v6348%now\, \$17121%now\, \$16752_fill6545929_arg%now\, \$v6382%now\, \$12853_forever6705887_arg%now\, \$v7251%now\, \$15769_binop_compare6455920_arg%now\, \$17494%now\, \$v6385%now\, \$14326%now\, \$v6240%now\, \$19080_next%now\, \$17386%now\, \$13982_v%now\, \$17459_loop665_arg%now\, \$18719_w%now\, \$15445%now\, \$v7353%now\, \$16752_fill6545929_result%now\, \$14997_modulo6685888_id%now\, \$18050%now\, \$12883%now\, \$16823_compbranch6505931_arg%now\, \$16233%now\, \$16271%now\, \$12682_make_block579_arg%now\, \$18655%now\, \$v7371%now\, \$18987_hd%now\, \$v6619%now\, \$v6427%now\, \$16748%now\, \$v6974%now\, \$18474%now\, \$17886%now\, \$15756_compare6445897_arg%now\, \$13151%now\, \$v6805%now\, \$17569%now\, \$12698%now\, \$15389_modulo6685895_arg%now\, \$v6035%now\, \$15553_r%now\, \$15237_modulo6685888_result%now\, \$12944%now\, \$14613_modulo6685896_result%now\, \$v7381%now\, \$18846%now\, \$18917%now\, \$v6092%now\, \$18916%now\, \$15261_modulo6685888_id%now\, \$17679%now\, \$13154%now\, \$v6336%now\, \$16527_f0%now\, \$18352%now\, \$13964%now\, \$v7420%now\, \$13632_next%now\, \$v6502%now\, \$v6370%now\, \$18739%now\, \$12714%now\, \$17484%now\, \$17597%now\, \$15756_compare6445897_result%now\, \$v7137%now\, \$13532%now\, \$v6823%now\, \$14781_modulo6685888_result%now\, \$v6721%now\, \$17734_copy_root_in_ram6635892_id%now\, \$v7338%now\, \$14749_modulo6685895_arg%now\, \$v7050%now\, \$16299_v%now\, \$12689%now\, \$18807%now\, \$13920_loop666_arg%now\, \$17455_loop666_id%now\, \$v6027%now\, \$18650%now\, \$18837%now\, \$16951_compare6445898_arg%now\, \$14861_modulo6685888_result%now\, \$18805%now\, \$17543%now\, \$13997_v%now\, \$16574_compare6445898_id%now\, \$v6728%now\, \$v6500%now\, \$v5869%now\, \$v6496%now\, \$14978_v%now\, \$v7454%now\, \$13237%now\, \$v6146%now\, \$15330_r%now\, \$12839%now\, \$14061_v%now\, \$14701_modulo6685888_arg%now\, \$12697%now\, \$17773%now\, \$v7344%now\, \$12888%now\, \$13155%now\, \$12937%now\, \$16115%now\, \$12805_aux664_result%now\, \$v6021%now\, \$13697%now\, \$v6466%now\, \$18355%now\, \rdy5940%now\, \$13102%now\, \$13235%now\, \$15044_binop_int6435906_id%now\, \$16729_v%now\, \$v6376%now\, \$13233%now\, \$17670%now\, \$14555%now\, \$14564_binop_int6435900_result%now\, \$v6802%now\, \$15058_v%now\, \$17464%now\, \$v6599%now\, \$v6430%now\, \$v6318%now\, \$v7161%now\, \$17669%now\, \$16963_compbranch6505935_id%now\, \$13967_v%now\, \$13696%now\, \$v6015%now\, \$15476_modulo6685895_arg%now\, \$17470%now\, \$12520_loop666_id%now\, \$18815%now\, \$v6559%now\, \$18565%now\, \$16551_compbranch6505926_id%now\, \$15397_modulo6685888_result%now\, \$12877%now\, \$18698%now\, \$18480%now\, \$v7300%now\, \$15389_modulo6685895_result%now\, \$v7144%now\, \$v6780%now\, \$19256_hd%now\, \$15823_res%now\, \$15124_binop_int6435907_id%now\, \$v6218%now\, \$v7406%now\, \$16963_compbranch6505935_arg%now\, \$v7132%now\, \$v7200%now\, \$18633_loop665_id%now\, \$17888%now\, \$19145%now\, \$15625_binop_compare6455916_id%now\, \$19337%now\, \$15893%now\, \$14364_v%now\, \$16893_compbranch6505933_result%now\, \$v6406%now\, \$v6489%now\, \$14837_modulo6685888_result%now\, \$14677_modulo6685888_arg%now\, \$v6667%now\, \$v7413%now\, \$v6508%now\, \$v6591%now\, \$16284_v%now\, \$12808_aux664_result%now\, \$13816%now\, \$v6211%now\, \$15874%now\, \$14829_modulo6685895_id%now\, \$v7027%now\, \$v6596%now\, \$17746%now\, \$13950%now\, \$v5963%now\, \$v5944%now\, \$14597_modulo6685888_result%now\, \$14582_res%now\, \$17891%now\, \$15397_modulo6685888_arg%now\, \$13927_branch_if648_result%now\, \$v7306%now\, \$v7074%now\, \$15021_modulo6685888_result%now\, \$12707%now\, \$16881_compare6445898_result%now\, \$13679_w%now\, \$13663%now\, \$18447%now\, \$v6732%now\, \$v6298%now\, \$v6518%now\, \$18278%now\, \$12544%now\, \$13218_w%now\, \$15932%now\, \$v7402%now\, \$v7085%now\, \$18731%now\, \$13519_w%now\, \$13606%now\, \$17776%now\, \$18644%now\, \$16327%now\, \$16169_v%now\, \$16551_compbranch6505926_arg%now\, \$15229_modulo6685895_arg%now\, \$17457_aux664_result%now\, \$v6633%now\, \$17665_hd%now\, \$18159%now\, \$v6058%now\, \$14122%now\, \$18563%now\, \$13310%now\, \$14012%now\, \$14677_modulo6685888_id%now\, \$14181_sp%now\, \$v6235%now\, \$15961%now\, \$15476_modulo6685895_result%now\, \$15237_modulo6685888_id%now\, \$17505_forever6705894_arg%now\, \$13388%now\, \$v6480%now\, \$17001%now\, \$17963%now\, \$17803%now\, \$19142%now\, \$18679_forever6705881_id%now\, \$v6291%now\, \$v6532%now\, \$v7293%now\, \$18919%now\, \$12685%now\, \$v6501%now\, \$17238_sp%now\, \$18186%now\, \$v7279%now\, \$v6460%now\, \$14431%now\, \$13667%now\, \$17455_loop666_arg%now\, \$12851%now\, \$18188%now\, \$v6172%now\, \$v7403%now\, \$v7216%now\, \$v7035%now\, \$v6397%now\, \$18709%now\, \$15720_compare6445897_id%now\, \$13823%now\, \$14177_hd%now\, \result6503%now\, \$13395%now\, \$16353%now\, \$v6239%now\, \$17559%now\, \$14351_v%now\, \$12808_aux664_id%now\, \$19269%now\, \$17412%now\, \$v7007%now\, \$v6941%now\, \$v6746%now\, \$18925%now\, \$v6838%now\, \$18733%now\, \$v5957%now\, \$v6953%now\, \$15783_v%now\, \$18279%now\, \$14207_loop_push6495899_result%now\, \$v6108%now\, \$v7025%now\, \$18120%now\, \$18566%now\, \$13016%now\, \$v6304%now\, \$12692%now\, \$16037_v%now\, \$12935%now\, \$13625%now\, \$v7434%now\, \$v6739%now\, \$17509_forever6705890_arg%now\, \$v6274%now\, \$19001%now\, \$v7290%now\, \$17498%now\, \$16945_b%now\, \$15298_v%now\, \$18346%now\, \$16589_compbranch6505927_id%now\, \$v6708%now\, \$13157%now\, \$18909_hd%now\, \$17674%now\, \$12712%now\, \$12945%now\, \$17354%now\, \$16574_compare6445898_result%now\, \$16365%now\, \$12715%now\, \$16510_forever6705925_id%now\, \$15218_v%now\, \$18699%now\, \$17591%now\, \$v6627%now\, \$12915%now\, \$v6136%now\, \$18045%now\, \$17460_aux664_id%now\, \$12807_loop665_id%now\, \$15069_modulo6685895_id%now\, \$v6492%now\, \$17487%now\, \$v6892%now\, \$17387%now\, \$15386_r%now\, \$v6729%now\, \$v6914%now\, \$18915%now\, \$17105_w06555936_id%now\, \$16589_compbranch6505927_arg%now\, \$13890%now\, \$19144%now\, \$16677%now\, \$v7034%now\, \$17678%now\, \$16875_b%now\, \$13927_branch_if648_arg%now\, \$v6883%now\, \$16438_v%now\, \$15612%now\, \$14773_modulo6685896_arg%now\, \$19140%now\, \$19071%now\, \$12848%now\, \$18831_hd%now\, \$v6710%now\, \$13468%now\, \$v6856%now\, \$15317_modulo6685888_result%now\, \$18570%now\, \$13623%now\, \$18128_next%now\, \$v7248%now\, \$14644_binop_int6435901_result%now\, \$12679_loop666_id%now\, \$16399%now\, \$19263%now\, \$14749_modulo6685895_id%now\, \$17794_w%now\, \result6468%now\, \$v7045%now\, \$18816%now\, \$17885%now\, \$v7164%now\, \$15101_modulo6685888_result%now\, \$v7042%now\, \$15500_modulo6685896_arg%now\, \$15333_modulo6685896_result%now\, \$17761_copy_root_in_ram6635891_result%now\, \$15720_compare6445897_arg%now\, \$16713_v%now\, \$15697_binop_compare6455918_arg%now\, \$17250_v%now\, \$12887%now\, \$v6826%now\, \$17394%now\, \$v6695%now\, \$17333_sp%now\, \$v7017%now\, \$16158_forever6705923_arg%now\, \$v6874%now\, \$v6574%now\, \$15853_v%now\, \$v7372%now\, \$v6651%now\, \$v7013%now\, \$15181_modulo6685888_result%now\, \$12691%now\, \$17962%now\, \$v6367%now\, \$v6200%now\, \$16612_compare6445898_result%now\, \$v6688%now\, \$14330_v%now\, \$v7361%now\, \$17319%now\, \$13941%now\, \$16078%now\, \$16165%now\, \$v7299%now\, \$17012_sp%now\, \$15261_modulo6685888_arg%now\, \$v6342%now\, \$v5954%now\, \$16606_b%now\, \$14986_r%now\, \$13301_hd%now\, \$15847%now\, \$v7179%now\, \$15021_modulo6685888_arg%now\, \$13127%now\, \$v7004%now\, \$v7090%now\, \$v6709%now\, \$17321%now\, \$13530%now\, \$14222%now\, \$v6868%now\, \$v6203%now\, \$v5866%now\, \$v5951%now\, \$18450%now\, \$13296_w%now\, \$14724_binop_int6435902_id%now\, \$v7400%now\, \$13013%now\, \$17349%now\, \$16192%now\, \$12834%now\, \$16441%now\, \$17167%now\, \$16042_v%now\, \$15697_binop_compare6455918_result%now\, \$12679_loop666_result%now\, \$16234%now\, \$15625_binop_compare6455916_result%now\, \$v7140%now\, \$18163%now\, \$v6007%now\, \$14933_modulo6685896_result%now\, \$v7066%now\, \$14818_v%now\, \$v6750%now\, \$15976_v%now\, \$v6935%now\, \$14338_v%now\, \$v6986%now\, \$16805_b%now\, \$17961%now\, \$16439_v%now\, \$14933_modulo6685896_id%now\, \$17681%now\, \$12910%now\, \$v6445%now\, \$12741%now\, \$v7455%now\, \$v6277%now\, \$v6962%now\, \$v7441%now\, \$13962%now\, \$15010_r%now\, \$14829_modulo6685895_result%now\, \$12521_loop665_arg%now\, \$14161%now\, \$15805_binop_compare6455921_arg%now\, \$12843%now\, \$15413_modulo6685896_result%now\, \$v7064%now\, \$15484_modulo6685888_arg%now\, \$v7368%now\, \$v6117%now\, \$18634_aux664_result%now\, \$12943%now\, \$v6995%now\, \$v6657%now\, \$17600%now\, \$v6214%now\, \$13957%now\, \$v7016%now\, \$v6307%now\, \$v6268%now\, \$18982_w%now\, \$13103%now\, \$14517_v%now\, \$v7023%now\, \$13692%now\, \$18479%now\, \$v7358%now\, \$v6271%now\, \$v6681%now\, \$12806_loop666_result%now\, \$12680_loop665_result%now\, \$18734%now\, \$15484_modulo6685888_id%now\, \$v6055%now\, \$14746_r%now\, \$17327%now\, \$13153%now\, \$v6701%now\, \$v7453%now\, \$v6950%now\, \$15733_binop_compare6455919_arg%now\, \$16436_v%now\, \$v7335%now\, \$14837_modulo6685888_arg%now\, \$14558%now\, \$v6609%now\, \$v6102%now\, \$v6865%now\, \$v7121%now\, \$v6175%now\, \$17520_copy_root_in_ram6635893_id%now\, \$18818%now\, \$17018_w36575938_id%now\, \$13946%now\, \$v7354%now\, \$17315%now\, \$15204_binop_int6435908_id%now\, \$14658_v%now\, \$13307%now\, \$14042%now\, \$12939%now\, \$12891_copy_root_in_ram6635884_arg%now\, \$v7416%now\, \$18166%now\, \$15556_modulo6685895_result%now\, \$16035%now\, \$14853_modulo6685896_arg%now\, \$15124_binop_int6435907_arg%now\, \$13928_w652_result%now\, \$15317_modulo6685888_arg%now\, \$17377%now\, \$16126%now\, \$v7133%now\, \$16127_v%now\, \$12878%now\, \$16031%now\, \$18836%now\, \$12857_forever6705883_arg%now\, \$v7219%now\, \$v6773%now\, \$14114%now\, \$v7086%now\, \$18999%now\, \$18637%now\, \$v6301%now\, \$17734_copy_root_in_ram6635892_arg%now\, \$v5874%now\, \$v7185%now\, \$13693%now\, \$v6229%now\, \$14285_v%now\, \$12734%now\, \$15341_modulo6685888_arg%now\, \$12904%now\, \$v7077%now\, \$17513_forever6705889_id%now\, \$v6853%now\, \$13466%now\, \$v7322%now\, \$14804_binop_int6435903_arg%now\, \$17463%now\, \$19115%now\, \$18904_w%now\, \$12818%now\, \$v6751%now\, \$16292%now\, \$12844_next%now\, \$16395_v%now\, \$14964_binop_int6435905_id%now\, \$16767%now\, \$15093_modulo6685896_arg%now\, \$v6103%now\, \$15648_compare6445897_id%now\, \$v6165%now\, \$18104%now\, \$v7030%now\, \$14613_modulo6685896_id%now\, \$v6738%now\, \$v6678%now\, \$17491%now\, \$13078_copy_root_in_ram6635885_id%now\, \$15981_v%now\, \$12560%now\, \$v7057%now\, \$v6364%now\, \$12702%now\, \$13312%now\, \$12520_loop666_arg%now\, \$15792_compare6445897_result%now\, \$15341_modulo6685888_result%now\, \$v7076%now\, \$14669_modulo6685895_id%now\, \$v5878%now\, \$18711%now\, \$15828_compare6445897_id%now\, \$15237_modulo6685888_arg%now\, \$v6183%now\, \$v5992%now\, \$v6314%now\, \$12522_wait662_result%now\, \$v6947%now\, \$v6595%now\, \$17455_loop666_result%now\, \$v7458%now\, \$v6162%now\, \$12838_next%now\, \$v6012%now\, \$18472%now\, \$16036_sp%now\, \$18185%now\, \$14424_v%now\, \$14254%now\, \$13389%now\, \$18677%now\, \$17348%now\, \$13393%now\, \$15769_binop_compare6455920_id%now\, \$13387%now\, \$17590%now\, \$v7398%now\, \$16823_compbranch6505931_id%now\, \$17495%now\, \$16379_v%now\, \$16881_compare6445898_arg%now\, \$18679_forever6705881_arg%now\, \$v6048%now\, \$14677_modulo6685888_result%now\, \$18288_next%now\, \$12538_cy%now\, \$15378_v%now\, \$12941%now\, \$17783%now\, \$13794%now\, \$14693_modulo6685896_arg%now\, \$12914%now\, \$19262%now\, \$v6847%now\, \$15382_res%now\, \$12521_loop665_result%now\, \$13238%now\, \$v6286%now\, \$19070%now\, \$17254%now\, \$13694%now\, \$14941_modulo6685888_arg%now\, \$v7328%now\, \$18356%now\, \$v7054%now\, \$17761_copy_root_in_ram6635891_id%now\, \$12695%now\, \$v6089%now\, \$17774%now\, \$16231%now\, \$v7015%now\, \$16202_ofs%now\, \$v7091%now\, \$16217_hd%now\, \$v6400%now\, \$v6388%now\, \$16024%now\, \$12913%now\, \$17048_w16565937_arg%now\, \$15476_modulo6685895_id%now\, \$16823_compbranch6505931_result%now\, \$16928_compbranch6505934_result%now\, \$18475%now\, \$17890%now\, \$15580_modulo6685896_id%now\, \$15828_compare6445897_result%now\, \$12936%now\, \$17165%now\, \$12660%now\, \$v7232%now\, \$12736%now\, \$v6724%now\, \$18724_hd%now\, \$17775%now\, \$16630%now\, \$15341_modulo6685888_id%now\, \$18187%now\, \$v6998%now\, \$17580_w%now\, \$17785%now\, \$12716%now\, \$15253_modulo6685896_id%now\, \$14135%now\, \$15828_compare6445897_arg%now\, \$13129%now\, \$18194%now\, \$18193%now\, \$16916_compare6445898_arg%now\, \$17812%now\, \$12806_loop666_id%now\, \$15204_binop_int6435908_result%now\, \$v7210%now\, \$17457_aux664_arg%now\, \$14453_next_acc%now\, \$18571%now\, \$15309_modulo6685895_result%now\, \$17879_hd%now\, \$13138_w%now\, \$v6624%now\, \$v6992%now\, \$14644_binop_int6435901_arg%now\, \$v6515%now\, \$13507%now\, \$19235%now\, \$17593%now\, \$17460_aux664_result%now\, \$v7283%now\, \$16986_compare6445898_result%now\, \$14930_r%now\, \$v6898%now\, \$v6003%now\, \$17466%now\, \$v6579%now\, \$v6121%now\, \$14621_modulo6685888_result%now\, \$13689%now\, \$14804_binop_int6435903_result%now\, \$12782%now\, \$18995%now\, \$v6110%now\, \$v6179%now\, \$18043%now\, \$19251_w%now\, \$14381%now\, \$v6066%now\, \$12546_dur%now\, \$v6911%now\, \$v6207%now\, \$15253_modulo6685896_result%now\, \$17889%now\, \$14311%now\, \$v6971%now\, \$v5999%now\, \$12906%now\, \$v7206%now\, \$14917_modulo6685888_id%now\, \$18661%now\, \$17957_hd%now\, \$12924_w%now\, \$v6546%now\, \$18280%now\, \$13148%now\, \$v6232%now\, \$18633_loop665_arg%now\, \$14757_modulo6685888_result%now\, \$13922_wait662_result%now\, \$v7364%now\, \$15580_modulo6685896_result%now\, \$15421_modulo6685888_id%now\, \$14610_r%now\, \$16916_compare6445898_id%now\, \$12886%now\, \$16195_forever6705924_id%now\, \$v6670%now\, \$13817%now\, \$v6817%now\, \$14221%now\, \$v6062%now\, \$17389%now\, \$v6563%now\, \$v6080%now\, \$v6799%now\, \$v7092%now\, \$14296%now\, \$17815%now\, \$v6463%now\, \$13100%now\, \$v6097%now\, \$v7203%now\, \$13808_hd%now\, \$13822%now\, \$16121_v%now\, \$v6403%now\, \$17000_sp%now\, \$12735%now\, \$v6424%now\, \$15261_modulo6685888_result%now\, \$17500%now\, \$17805%now\, \$v6421%now\, \$13510%now\, \$13940%now\, \$v7433%now\, \$15309_modulo6685895_arg%now\, \$18657%now\, \$16574_compare6445898_arg%now\, \$13317%now\, \$v6287%now\, \$12903%now\, \$16382%now\, \$15897%now\, \$14941_modulo6685888_result%now\, \$14909_modulo6685895_result%now\, \$v7135%now\, \$18806%now\, \$17458_loop666_arg%now\, \$12938%now\, \$15531_binop_int6435913_id%now\, \$15284_binop_int6435909_id%now\, \$13700%now\, \$18843%now\, \$15364_binop_int6435910_id%now\, \$12523_make_block579_arg%now\, \$v7245%now\, \$16317%now\, \$18348%now\, \$13101%now\, \$v6069%now\, \$16063_w6515922_result%now\, \$v6096%now\, \$12864_copy_root_in_ram6635886_arg%now\, \$14669_modulo6685895_arg%now\, \$17561%now\, \$19118%now\, \$14837_modulo6685888_id%now\, \$12694%now\, \$15284_binop_int6435909_arg%now\, \$12701%now\, \$v7450%now\, \$16158_forever6705923_id%now\, \$15101_modulo6685888_id%now\, \$v7145%now\, \$v6654%now\, \$v6042%now\, \$13234%now\, \$v6717%now\, \$15580_modulo6685896_arg%now\, \$15500_modulo6685896_result%now\, \$15447_forever6705911_arg%now\, \$18189%now\, \rdy6469%now\, \$17964%now\, \$18319%now\, \$v6920%now\, \$v6989%now\, \$14315_v%now\, \$18124%now\, \$16321%now\, \$v5986%now\, \$13384%now\, \$13379_hd%now\, \$15421_modulo6685888_arg%now\, \$v7365%now\, \$13922_wait662_id%now\, \$12549%now\, \$v6832%now\, \$v6765%now\, \$v6104%now\, \$18730%now\, \$18184%now\, \$17892%now\, \$v6543%now\, \$v6585%now\, \$17671%now\, \$v6106%now\, \$12704%now\, \$v7399%now\, \$v7110%now\, \$18118%now\, \$13540%now\, \$v6862%now\, \$15508_modulo6685888_result%now\, \$v7100%now\, \$17513_forever6705889_arg%now\, \$v6835%now\, \$16203%now\, \$15229_modulo6685895_result%now\, \$15910%now\, \$17456_loop665_result%now\, \$v5995%now\, \$13765%now\, \$12807_loop665_result%now\, \$v6373%now\, \$v6171%now\, \$18473%now\, \$v6758%now\, \$v7332%now\, \$v6646%now\, \$v6692%now\, \$v7188%now\, \$16063_w6515922_id%now\, \$v6562%now\, \$v6743%now\, \$v7426%now\, \$13463%now\, \$18686_copy_root_in_ram6635880_id%now\, \$v7378%now\, \$v6742%now\, \$14989_modulo6685895_result%now\, \$v7375%now\, \$15204_binop_int6435908_arg%now\, \$18845%now\, \$14008%now\, \$v6328%now\, \$v7355%now\, \$v7044%now\, \$v6319%now\, \$15364_binop_int6435910_arg%now\, \$v6965%now\, \$12879%now\, \$15284_binop_int6435909_result%now\, \$12804_loop665_result%now\, \$18546%now\, \$v7020%now\, \$15564_modulo6685888_result%now\, \$v7081%now\, \$v5872%now\, \$v7393%now\, \$14152%now\, \$v6766%now\, \$18841%now\, \$15661_binop_compare6455917_result%now\, \$13316%now\, \$13009_hd%now\, \$14909_modulo6685895_arg%now\, \$12682_make_block579_result%now\, \$18738%now\, \$16509%now\, \$12688%now\, \$15577_r%now\, \$v6093%now\, \$v6109%now\, \$15564_modulo6685888_arg%now\, \$16928_compbranch6505934_id%now\, \$14884_binop_int6435904_arg%now\, \$v6553%now\, \$14092%now\, \$v6535%now\, \$18732%now\, \$17066%now\, \$15389_modulo6685895_id%now\, \$v6660%now\, \$17337%now\, \$18826_w%now\, \$v6036%now\, \$17374_v%now\, \$17502%now\, \$12942%now\, \$14773_modulo6685896_id%now\, \$14757_modulo6685888_id%now\, \$18041%now\, \$v6547%now\, \$v6184%now\, \$12864_copy_root_in_ram6635886_id%now\, \$18470%now\, \$12835%now\, \$15909%now\, \$v6902%now\, \$17009_sp%now\, \$18476%now\, \$16626%now\, \$17804%now\, \$18443%now\, \$14701_modulo6685888_result%now\, \$v7167%now\, \$14902_res%now\, \$12717%now\, \$v6908%now\, \$13917%now\, \$16749_sp%now\, \$v6155%now\, \$17243%now\, \$v6442%now\, \$13923_make_block579_result%now\, \$v7445%now\, \$v6354%now\, \$14508_v%now\, \$15157_modulo6685888_arg%now\, \$19267%now\, \$16846_compare6445898_id%now\, \$15170_r%now\, \$v6616%now\, \$13926_make_block_n646_id%now\, \$18478%now\, \$16440%now\, \$15451_binop_int6435912_arg%now\, \$15980_v%now\, \$v6623%now\, \$14909_modulo6685895_id%now\, \$12830%now\, \$13149%now\, \$17164%now\, \$14463_v%now\, \$13019%now\, \$15613%now\, \$17535%now\, \$13818%now\, \$v6521%now\, \$16763_v%now\, \$18669%now\, \$18660%now\, \$v6137%now\, \$v6790%now\, \$v7117%now\, \$v6223%now\, \$13105_copy_root_in_ram6635884_arg%now\, \$v7387%now\, \$17547_copy_root_in_ram6635891_id%now\, \$15157_modulo6685888_id%now\, \$18632_loop666_arg%now\, \$17173%now\, \$15447_forever6705911_id%now\, \$15861_v%now\, \$13223_hd%now\, \$13524_hd%now\, \$16336%now\, \$v6899%now\, \$v7156%now\, \$15302_res%now\, \$19268%now\, \$18572%now\, \$v7459%now\, \$v7229%now\, \$17883%now\, \$18048%now\, \$13385%now\, \$17239_v%now\, \$14773_modulo6685896_result%now\, \$17592%now\, \$13926_make_block_n646_result%now\, \$17749%now\, \$18668%now\, \$v7093%now\, \$v6176%now\, \$12710%now\, \$18913%now\, \$v7107%now\, \$v6075%now\, \$v6031%now\, \$14861_modulo6685888_arg%now\, \$v6352%now\, \$13924_apply638_result%now\, \$15883%now\, \$v6684%now\, \$13309%now\, \$12829%now\, \$14273%now\, \rdy6504%now\, \$v6938%now\, \$17371_v%now\, \$v6880%now\, \$v7011%now\, \$17232%now\, \$12864_copy_root_in_ram6635886_result%now\, \$v6829%now\, \$v7056%now\, \$14139%now\, \$v6379%now\, \$17332_sp%now\, \$17048_w16565937_result%now\, \$19266%now\, \$15588_modulo6685888_result%now\, \$v7260%now\, \$14621_modulo6685888_arg%now\, \$13924_apply638_arg%now\, \$v6643%now\, \$v6152%now\, \$18994%now\, \$15250_r%now\, \$15044_binop_int6435906_result%now\, \$16650_sp%now\, \$v7350%now\, \$18633_loop665_result%now\, \$12553%now\, \$18044%now\, \$12720%now\, \$17594%now\, \$v6190%now\, \$v5964%now\, \$13926_make_block_n646_arg%now\, \$15077_modulo6685888_id%now\, \$v7021%now\, \$17018_w36575938_result%now\, \$v6180%now\, \$v6889%now\, \$15715_res%now\, \$16349_v%now\, \$14964_binop_int6435905_arg%now\, \$18998%now\, \$13158%now\, \$v6283%now\, \$17393%now\, \$v5948%now\, \$13092%now\, \$v6714%now\, \$v6325%now\, \$14997_modulo6685888_result%now\, \$v6550%now\, \$v6236%now\, \$12934%now\, \$v6588%now\, \$v6256%now\, \$17458_loop666_id%now\, \$17032%now\, \$12706%now\, \$16673_v%now\, \$13688%now\, \$v7427%now\, \$17458_loop666_result%now\, \$12681_wait662_arg%now\, \$18673%now\, \$17324%now\, \$14070_v%now\, \$12737%now\, \$19214%now\, \$15787_res%now\, \$14589_modulo6685895_arg%now\, \$v5967%now\, \$17968%now\, \$14738_v%now\, \$v5998%now\, \$18639%now\, \$13766%now\, \$15413_modulo6685896_arg%now\, \$15860%now\, \$v7010%now\, \$18564%now\, \$v7449%now\, \$v7046%now\, \$17532%now\, \$v6243%now\, \$19213%now\, \$13529%now\, \$v6493%now\, \$15421_modulo6685888_result%now\, \$18191%now\, \$14564_binop_int6435900_id%now\, \$12679_loop666_arg%now\, \$14406_v%now\, \$15619%now\, \$v6917%now\, \$16507%now\, \$v7116%now\, \$v7273%now\, \$14165%now\, \$13920_loop666_id%now\, \$15618%now\, \$16403%now\, \$17476%now\, \$13626%now\, \$17967%now\, \$12709%now\, \$v7213%now\, \$14861_modulo6685888_id%now\, \$v6844%now\, \$12804_loop665_arg%now\, \$14281%now\, \$16272%now\, \$17572%now\, \$12705%now\, \$12696%now\, \$13117%now\, \$13605%now\, \$16288%now\, \$12853_forever6705887_id%now\, \$17734_copy_root_in_ram6635892_result%now\, \$17759%now\, \$v6247%now\, \$16986_compare6445898_id%now\, \$17314%now\, \$v7197%now\, \$12680_loop665_arg%now\, \$18119%now\, \$v6072%now\, \$12760%now\, \$12548_dis%now\, \$15077_modulo6685888_arg%now\, \$14853_modulo6685896_result%now\, \$18737%now\, \$18918%now\, \$17237_sp%now\, \$15173_modulo6685896_arg%now\, \$17595%now\, \$17008%now\, \$17761_copy_root_in_ram6635891_arg%now\, \$v7101%now\, \$12847%now\, \$v6859%now\, \$12889%now\, \$18051%now\, \$v6219%now\, \$14826_r%now\, \$14033%now\, \$v6606%now\, \$18326%now\, \$18921%now\, \$13691%now\, \$v7083%now\, \$v6956%now\, \$15679_res%now\, \$v6666%now\, \$19239%now\, \$14024%now\, \$v7442%now\, \$16811_compare6445898_result%now\, \$14781_modulo6685888_arg%now\, \$v6335%now\, \$19260%now\, \$17347%now\, \$15333_modulo6685896_id%now\, \$18196%now\, \$v6752%now\, \$16300%now\, \$17673%now\, \$13227%now\, \$16612_compare6445898_arg%now\, \$13925_offsetclosure_n639_result%now\, \$v6409%now\, \$17814%now\, \$17585_hd%now\, \$17509_forever6705890_id%now\, \$17566%now\, \$12814%now\, \$19242%now\, \$17497%now\, \$13695%now\, \$v6394%now\, \$v7397%now\, \$v7289%now\, \$v7194%now\, \$17874_w%now\, \$18844%now\, \$15181_modulo6685888_arg%now\, \$18175_w%now\, \$v5876%now\, \$18676%now\, \$17539%now\, \$v7115%now\, \$v6263%now\, \$v6353%now\, \$18335_w%now\, \$18993%now\, \$13928_w652_id%now\, \$17504%now\, \$18046%now\, \$12670%now\, \$v5972%now\, \$v6133%now\, \$12743%now\, \$13539%now\, \$v5947%now\, \$17117_v%now\, \$15173_modulo6685896_result%now\, \$15819_v%now\, \$17547_copy_root_in_ram6635891_arg%now\, \$12681_wait662_id%now\, \$14043_v%now\, \$13814%now\, \$12803_loop666_arg%now\, \$v6436%now\, \$19136%now\, \$18674%now\, \$v6784%now\, \$v7296%now\, \$17395%now\, \$13236%now\, \$13464%now\, \$14051%now\, \$v7014%now\, \$17320%now\, \$v7095%now\, \$v6433%now\, \$12681_wait662_result%now\, \$13383%now\, \$14578_v%now\, \$v7112%now\, \$17675%now\, \$19127_w%now\, \$18808%now\, \$14148%now\, \$18705%now\, \$14804_binop_int6435903_id%now\, \$v6650%now\, \$v7267%now\, \$13624%now\, \$15588_modulo6685888_arg%now\, \$v7051%now\, \$v5867%now\, \$17388%now\, \$15173_modulo6685896_id%now\, \$16589_compbranch6505927_result%now\, \$14069%now\, \$v6531%now\, \$12713%now\, \$13021%now\, \$18666_next%now\, \$14446_v%now\, \$17677%now\, \$18740%now\, \$18842%now\, \$17972%now\, \$14989_modulo6685895_id%now\, \$17598%now\, \$12522_wait662_id%now\, \$18701%now\, \$16662_fill6535928_arg%now\, \$17490_next%now\, \$v6759%now\, \$16928_compbranch6505934_arg%now\, \$18922%now\, \$18464_hd%now\, \$16963_compbranch6505935_result%now\, \$13992_v%now\, \$15508_modulo6685888_arg%now\, \$12929_hd%now\, \$v7457%now\, \$13538%now\, \$16457%now\, \$15306_r%now\, \$v6705%now\, \$18122%now\, \$v7102%now\, \$19143%now\, \$18670_next%now\, \$18634_aux664_arg%now\, \$18793_copy_root_in_ram6635879_id%now\, \$15149_modulo6685895_id%now\, \$16788_compbranch6505930_result%now\, \$13535%now\, \$15545_v%now\, \$17482%now\, \$v7061%now\, \$v6253%now\, \$13897%now\, \$18735%now\, \$v7126%now\, \$18281%now\, \$16473%now\, \$14917_modulo6685888_result%now\, \$16741%now\, \$16510_forever6705925_arg%now\, \$v6536%now\, \$12811%now\, \$v6796%now\, \$18459_w%now\, \$14413_v%now\, \$12520_loop666_result%now\, \$16612_compare6445898_id%now\, \$17747%now\, \$v7104%now\, \$13939%now\, \$15661_binop_compare6455917_id%now\, \$17973%now\, \$12804_loop665_id%now\, \$17758%now\, \$12719%now\, \$15397_modulo6685888_id%now\, \$17105_w06555936_arg%now\, \$12792%now\, \$16194%now\, \$v7176%now\, \$14829_modulo6685895_arg%now\, \$18049%now\, \$13536%now\, \$12842%now\, \$v7182%now\, \$v6511%now\, \$14693_modulo6685896_id%now\, \$13023%now\, \$v6098%now\, \$15792_compare6445897_arg%now\, \$v6905%now\, \$13313%now\, \$14552%now\, \$16840_b%now\, \$16568_b%now\, \$14423_v%now\, \$v6527%now\, \$18262%now\, \$13078_copy_root_in_ram6635885_result%now\, \$18351%now\, \$16232%now\, \$16133%now\, \$15711_v%now\, \$15614_forever6705914_id%now\, \$13004_w%now\, \$12803_loop666_id%now\, \$12744%now\, \$13311%now\, \$18664_next%now\, \$19264%now\, \$13472_next%now\, \$16858_compbranch6505932_id%now\, \$v7096%now\, \$17966%now\, \$v6787%now\, \$17459_loop665_result%now\, \$v7120%now\, \$17310%now\, \$17492_next%now\, \$v6045%now\, \$17748%now\, \$18638%now\, \$15792_compare6445897_id%now\, \$13963%now\, \$v6140%now\, \$12933%now\, \$18640%now\, \$13528%now\, \$v7254%now\, \$16881_compare6445898_id%now\, \$17460_aux664_arg%now\, \$12523_make_block579_result%now\, \$13922_wait662_arg%now\, \$v6156%now\, \$v6814%now\, \$v7419%now\, \$15451_binop_int6435912_result%now\, \$v6322%now\, \$17331_sp%now\, \$17894%now\, \$v6002%now\, \$v6476%now\, \$13239%now\, \$12708%now\, \$18812%now\, \$v6187%now\, \$v7072%now\, \rdy6148%now\, \$18047%now\, \$14644_binop_int6435901_id%now\, \$14597_modulo6685888_id%now\, \$v7103%now\, \$19261%now\, \$16893_compbranch6505933_arg%now\, \$13390%now\, \$16534%now\, \$v7191%now\, \$19002%now\, \$v7041%now\, \$v6968%now\, \$v7127%now\, \$17520_copy_root_in_ram6635893_result%now\, \$v6332%now\, \$13229%now\, \$v6159%now\, \$15684_compare6445897_id%now\, \$v7114%now\, \$17544%now\, \$v6704%now\, \$18040%now\, \$17786%now\, \$v7233%now\, \$14207_loop_push6495899_arg%now\, \$16709%now\, \$v7113%now\, \$14724_binop_int6435902_arg%now\, \$13232%now\, \$16986_compare6445898_arg%now\, \$v6054%now\, \$16074_v%now\, \$v6781%now\, \$v7047%now\, \$17503%now\, \$13147%now\, \$v6259%now\, \$v6144%now\, \$13018%now\, \$v6603%now\, \$14016_v%now\, \$16752_fill6545929_id%now\, \$v5973%now\, \$13815%now\, \$v7033%now\, \$v5983%now\, \$19271%now\, \$v6735%now\, \$v6769%now\, \$v7242%now\, \$16508%now\, \$12808_aux664_arg%now\, \$18708%now\, \$18991%now\, \$14471%now\, \$v7070%now\, \$12547%now\, \$v7031%now\, \$v6315%now\, \$12674%now\, \$12846%now\, \$17010%now\, \$17560%now\, \$16156%now\, \$15021_modulo6685888_id%now\, \$13925_offsetclosure_n639_arg%now\, \$14898_v%now\, \$14693_modulo6685896_result%now\, \$15497_r%now\, \$13105_copy_root_in_ram6635884_id%now\, \$17434%now\, \$16515%now\, \$14512_v%now\, \$14300_v%now\, \$18261%now\, \$17207_arg%now\, \$13315%now\, \$18992%now\, \$18344%now\, \$17183%now\, \$v7032%now\, \result6112%now\, \$v5960%now\, \$v7084%now\, \$v6639%now\, \$v7060%now\, \$18030_w%now\, \$18190%now\, \$16380_v%now\, \$v6295%now\, \$18924%now\, \$12659%now\, \$v6111%now\, \$v6011%now\, \$12891_copy_root_in_ram6635884_result%now\, \$18621%now\, \$14185_next_env%now\, \$17166%now\, \$v6059%now\, \$12703%now\, \$v6358%now\, \$12832%now\, \$15684_compare6445897_result%now\, \$v7111%now\, \$17895%now\, \$13812%now\, \$18632_loop666_id%now\, \$17952_w%now\, \$13820%now\, \$13533%now\, \$15805_binop_compare6455921_result%now\, \$15413_modulo6685896_id%now\, \$13977_v%now\, \$v6294%now\, \$12857_forever6705883_id%now\, \$v7438%now\, \$v7082%now\, \$v6415%now\, \$v5982%now\, \$19265%now\, \$17011%now\, \$v7012%now\, \$17505_forever6705894_id%now\, \$v7282%now\, \$12813%now\, \$17499%now\, \$v6457%now\, \$13150%now\, \$17808%now\, \$v6820%now\, \$17970%now\, \$12803_loop666_result%now\, \$v7276%now\, \$14964_binop_int6435905_result%now\, \$v7134%now\, \$17809%now\, \$16404%now\, \$v7157%now\, \$17969%now\, \$v6280%now\, \$12845%now\, \$v6361%now\, \$12561%now\, \$17545%now\, \$18634_aux664_id%now\, \$15410_r%now\, \$v6582%now\, \$v6600%now\, \$15062_res%now\, \$v6264%now\, \$14342%now\, \$v6691%now\, \$12562%now\, \result5939%now\, \$12657%now\, \$v7130%now\, \$16193%now\, \$16916_compare6445898_result%now\, \$18839%now\, \$13787%now\, \$v7303%now\, \$19146%now\, \$15684_compare6445897_arg%now\, \$15142_res%now\, \$12905%now\, \$v6267%now\, \$18658%now\, \$13386%now\, \$17465%now\, \$v6477%now\, \$13025%now\, \$18678%now\, \$16461%now\, \$v6774%now\, \$18180_hd%now\, \$v6811%now\, \$13791%now\, \$14464_v%now\, \$15851_argument1%now\, \$13022%now\, \$15101_modulo6685888_arg%now\, \$13124%now\, \$v6762%now\, \$v6720%now\, \$v6528%now\, \$v6083%now\, \$16724%now\, \$v6524%now\, \$v6448%now\, \$17184%now\, \$13228%now\, \$19139%now\, \$v7036%now\, \$v6755%now\, \$17533%now\, \result5974%now\, \$v7037%now\, \$18589%now\, \$14669_modulo6685895_result%now\, \$13813%now\, \$17105_w06555936_result%now\, \$13921_loop665_arg%now\, \$17599%now\, \$13921_loop665_result%now\, \$v7401%now\, \$v6980%now\, \$16337%now\, \$17534%now\, \$12558%now\, \$v6926%now\, \$16811_compare6445898_id%now\, \$v5989%now\, \$14103%now\, \$15556_modulo6685895_arg%now\, \$19147%now\, \$16383%now\, \$v7149%now\, \$13314%now\, \$15639_v%now\, \$16624_argument2%now\, \$15069_modulo6685895_result%now\, \$16662_fill6535928_id%now\, \rdy6113%now\, \$17542%now\, \$v6345%now\, \$v6194%now\, \$v6571%now\, \$15531_binop_int6435913_result%now\, \$v6439%now\, \$v6079%now\, \$15621_forever6705915_arg%now\, \$17884%now\, \$v7097%now\, \$13927_branch_if648_id%now\, \$14982_res%now\, \$18353%now\, \$v7347%now\, \$16846_compare6445898_arg%now\, \$v6895%now\, \$16195_forever6705924_arg%now\, \$17589%now\, \$13017%now\, \$15747_v%now\, \$16662_fill6535928_result%now\, \$18345%now\, \$v7122%now\, \$17048_w16565937_id%now\, \$18686_copy_root_in_ram6635880_result%now\, \$15093_modulo6685896_id%now\, \$18736%now\, \$18671%now\, \$15500_modulo6685896_id%now\, \$v7226%now\, \$17459_loop665_id%now\, \$15333_modulo6685896_arg%now\, \$17807%now\, \$v6220%now\, \$13821%now\, \$18035_hd%now\, \$v6290%now\, \$17172%now\, \$13394%now\, \$19338%now\, \$17368_v%now\, \$v5871%now\, \$13958%now\, \$12824%now\, \$17562%now\, \$16322%now\, \$v7105%now\, \$13698%now\, \$17520_copy_root_in_ram6635893_arg%now\, \$15556_modulo6685895_id%now\, \$13105_copy_root_in_ram6635884_result%now\, \$12891_copy_root_in_ram6635884_id%now\, \$12806_loop666_arg%now\, \$v6566%now\, \$15181_modulo6685888_id%now\, \$v7080%now\, \$v6675%now\, \$v6576%now\, \$16998_argument3%now\, \$v7423%now\, \$18728%now\, \$16157%now\, \$13684_hd%now\, \$19111%now\, \$v6647%now\, \$13091%now\, \$13143_hd%now\, \$18793_copy_root_in_ram6635879_result%now\, \$15769_binop_compare6455920_result%now\, \$16462%now\, \$14265%now\, \$12916%now\, \$v6244%now\, \$12742%now\, \$13119%now\, \$13972_v%now\, \$14884_binop_int6435904_result%now\, \$13951%now\, \$v7024%now\, \$13923_make_block579_arg%now\, \$15648_compare6445897_result%now\, \$17330_sp%now\, \$v6620%now\, \$17353%now\, \$v6983%now\, \$v7257%now\, \$v6663%now\, \$13118%now\, \$v6032%now\, \$18672%now\, \$19074%now\, \$15309_modulo6685895_id%now\, \$v6260%now\, \$19076%now\, \rdy5975%now\, \$15124_binop_int6435907_result%now\, \$16334_v%now\, \$v7270%now\, \$18042%now\, \$18611%now\, \$14377_v%now\, \$16381_v%now\, \$v6076%now\, \$15908%now\, \$12563%now\, \$v7026%now\, \$v6698%now\, \$15013_modulo6685896_result%now\, \$12805_aux664_arg%now\, \$v7075%now\, \$13024%now\, \$13965%now\, \$18573%now\, \$v6124%now\, \$17481%now\, \$v6215%now\, \$15720_compare6445897_result%now\, \$v7160%now\, \$v6497%now\, \$15044_binop_int6435906_arg%now\, \$13097%now\, \$17456_loop665_arg%now\, \$13952%now\, \$15093_modulo6685896_result%now\, \$13924_apply638_id%now\, \$v6556%now\, \$14701_modulo6685888_id%now\, \$12687%now\, \$15473_r%now\, \$17061%now\, \$16725%now\, \$v6412%now\, \$v7407%now\, \$v6747%now\, \$12831%now\, \$16651%now\, \$14781_modulo6685888_id%now\, \$16658%now\, \$v7136%now\, \$14589_modulo6685895_id%now\, \$v5968%now\, \$v6339%now\, \$16788_compbranch6505930_id%now\, \$17486%now\, \$v6331%now\, \$18553%now\, \$14034_v%now\, \$v7410%now\, \$v7131%now\, \$18284%now\, \$v7390%now\, \$13306%now\, \$v6539%now\, \$v7341%now\, \$15090_r%now\, \$14906_r%now\, \$13462%now\, \$19270%now\, \$v6850%now\, \$v7430%now\, \$v6671%now\, \$15149_modulo6685895_result%now\, \$15756_compare6445897_id%now\, \$v6418%now\, \$v6250%now\, \$v6051%now\, \$15621_forever6705915_id%now\, \$v6886%now\, \$16858_compbranch6505932_result%now\, \$15222_res%now\, \$v6770%now\, \$v7040%now\, \$16301%now\, \$13911%now\, \$17680%now\, \$v6191%now\, \$15138_v%now\, \$v6486%now\, \$13152%now\, \$16155%now\, \$14933_modulo6685896_arg%now\, \$12693%now\, \$v7106%now\, \$v7067%now\, \$13920_loop666_result%now\, \$16293%now\, \$13159%now\, \$13953%now\, \$15625_binop_compare6455916_arg%now\, \$13015%now\, \$17799_hd%now\, \$v6039%now\, \$15611%now\, \$v6808%now\, \$17444%now\, \$14853_modulo6685896_id%now\, \$18665%now\, \$19132_hd%now\, \$16313_v%now\, \$14757_modulo6685888_arg%now\, \$18710%now\, \$v5979%now\, \$v6006%now\, \$14621_modulo6685888_id%now\, \$14941_modulo6685888_id%now\, \$19073%now\, \$15733_binop_compare6455919_id%now\, \$15620%now\, \$17596%now\, \$16413%now\, \$19141%now\, \$17753%now\, \$16706%now\, \$16296%now\, \$v7001%now\, \$18468%now\, \$19000%now\, \$v5877%now\, \$16951_compare6445898_id%now\, \$13231%now\, \$v6024%now\, \$13130%now\, \$15469_res%now\, \$18471%now\, \$v6793%now\, \$v7266%now\, \$18350%now\, \$16357%now\, \$15149_modulo6685895_arg%now\, \$13987_v%now\, \$v7055%now\, \$17483%now\, \$14260%now\, \$15588_modulo6685888_id%now\, \$v7309%now\, \$15643_res%now\, \$13078_copy_root_in_ram6635885_arg%now\, \$18914%now\, \$17660_w%now\, \$16846_compare6445898_result%now\, \$18817%now\, \$v6871%now\, \$17672%now\, \$19148%now\, \$v7329%now\, \$19072%now\, \$15733_binop_compare6455919_result%now\, \$14081%now\, \$18545%now\, \$13889%now\, \$14015%now\, \$12840_next%now\, \$18686_copy_root_in_ram6635880_arg%now\, \$14742_res%now\, \$14586_r%now\, \$18195%now\, \$v6540%now\, \$18793_copy_root_in_ram6635879_arg%now\, \$15317_modulo6685888_id%now\, \$16551_compbranch6505926_result%now\, \$17811%now\, \$16980_b%now\, \$18349%now\, \$15451_binop_int6435912_id%now\, \$14002_v%now\, \$14997_modulo6685888_arg%now\, \$16335_v%now\, \$13014%now\, \$v6977%now\, \$18039%now\, \$13448%now\, \$17571%now\, \$17757%now\, \$v6018%now\, \$16358%now\, \$v7052%now\, \$17352%now\, \$17756%now\, \$v6141%now\, \$13391%now\, \$v6086%now\, \$v6145%now\, \$15066_r%now\, \result6147%now\, \$15446%now\, \$v6877%now\, \$16041_v%now\, \$16063_w6515922_arg%now\, \$12700%now\, \$16951_compare6445898_result%now\, \$v6210%now\, \$15564_modulo6685888_id%now\, \$12721%now\, \$18920%now\, \$14393_hd%now\, \$18282%now\, \$v7141%now\, \$15157_modulo6685888_result%now\, \$14850_r%now\, \$17601%now\, \$v6310%now\, \$14493_v%now\, \$12711%now\, \$v5864%now\, \$v6483%now\, \$13819%now\, \$v7325%now\, \$13120%now\, \$v7087%now\, \$v6615%now\, \$15146_r%now\, \$v7394%now\, \$18347%now\, \$18700%now\, \$v6777%now\, \$12940%now\, \$v7173%now\, \$17062%now\, \$v7073%now\, \$14025_v%now\, \$14561%now\, \$16437_v%now\, \$15549_res%now\, \$15253_modulo6685896_arg%now\, \$15013_modulo6685896_arg%now\, \$14822_res%now\, \$18847%now\, \$18840%now\, \$18340_hd%now\, \$v7148%now\, \$14884_binop_int6435904_id%now\, \$18632_loop666_result%now\, \$15226_r%now\, \$18422%now\, \$15444%now\, \$19137%now\, \$18923%now\, \$17161%now\, \$12662%now\, \$v7065%now\, \$14662_res%now\, \$v6226%now\, \$v7319%now\, \$17396%now\, \$17806%now\, \$v6612%now\, \$15805_binop_compare6455921_id%now\, \$13305%now\, \$13230%now\, \$19056%now\, \$18469%now\, \$v7286%now\, \$13534%now\, \$v7152%now\, \$v6929%now\, \$16910_b%now\, \$v7043%now\, \$12850%now\, \$17456_loop665_id%now\, \$18477%now\, \$v7225%now\, \$v6923%now\, \$v6674%now\, \$13699%now\, \$v6944%now\, \$13923_make_block579_id%now\, \$14207_loop_push6495899_id%now\, \$15648_compare6445897_arg%now\, \$13803_w%now\, \$17780%now\, \$12876%now\, \$18656%now\, \$v6687%now\, \$v6107%now\, \$12661%now\, \$v6630%now\, \$15697_binop_compare6455918_id%now\, \$v7124%now\, \$v7384%now\, \$v7063%now\, \$13928_w652_arg%now\, \$15465_v%now\, \$13622%now\, \$14355%now\, \$v7312%now\, \$v6636%now\, \$14770_r%now\, \$v6063%now\, \$15013_modulo6685896_id%now\, \$14690_r%now\, \$12807_loop665_arg%now\, \$v6120%now\, \$17810%now\, \$v6168%now\, \$v7053%now\, \$v7239%now\, \$17236%now\, \$v7209%now\, \$13128%now\, \$15229_modulo6685895_id%now\, \$v7316%now\, \$12690%now\, \$13925_offsetclosure_n639_id%now\, \$13020%now\, \$v6932%now\, \$12539%now\, \$v6592%now\, \$v6010%now\, \$13093%now\, \$18323%now\, \$17965%now\, \$v5971%now\, \$16659_sp%now\, \$17547_copy_root_in_ram6635891_result%now\, \$13690%now\, \$13628%now\, \$v6349%now\, \$13465%now\, \$12812%now\, \$v6028%now\, \$13374_w%now\, \$14368%now\, \$12718%now\, \$17784%now\, \$15508_modulo6685888_id%now\, \$15364_binop_int6435910_result%now\, \$14613_modulo6685896_arg%now\, \$15751_res%now\, \$13537%now\, \$12654%now\, \$v7071%now\, \$v6311%now\, \$ram_lock%now\, \$global_end_lock%now\, \$code_lock%now\)
        variable \$12670\ : value(0 to 1) := (others => '0');
        variable \$12807_loop665_arg\, \$16651\, \$17456_loop665_arg\, 
                 \$13921_loop665_arg\, \$12523_make_block579_result\, 
                 \$17105_w06555936_arg\, \$16741\, \$12680_loop665_arg\, 
                 \$12804_loop665_arg\, \$17232\, 
                 \$13923_make_block579_result\, 
                 \$12682_make_block579_result\, \$18633_loop665_arg\, 
                 \$16024\, \$12521_loop665_arg\, \$17001\, 
                 \$17459_loop665_arg\ : value(0 to 95) := (others => '0');
        variable \$13928_w652_arg\, \$16063_w6515922_arg\, 
                 \$12805_aux664_arg\, \$12806_loop666_arg\, 
                 \$12808_aux664_arg\, \$14207_loop_push6495899_arg\, 
                 \$17460_aux664_arg\, \$18634_aux664_arg\, 
                 \$12803_loop666_arg\, \$12679_loop666_arg\, 
                 \$18632_loop666_arg\, \$17458_loop666_arg\, 
                 \$17457_aux664_arg\, \$12520_loop666_arg\, 
                 \$17455_loop666_arg\, \$13920_loop666_arg\ : value(0 to 63) := (others => '0');
        variable \$18323\, \$17780\, \$17753\, \$13097\, \$13124\, \$13791\, 
                 \$18812\, \$18705\, \$17539\, \$17566\, \$19239\, 
                 \$12548_dis\, \$17324\, \$12835\, \$18661\, \$13507\, 
                 \$12818\, \$19115\, \$17327\, \$12910\, \$18163\, \$17321\, 
                 \$17487\, \$13667\, \$18644\, \$18447\, \$17470\, \$12883\ : value(0 to 47) := (others => '0');
        variable \$15648_compare6445897_arg\, \$16846_compare6445898_arg\, 
                 \$15684_compare6445897_arg\, \$16986_compare6445898_arg\, 
                 \$15792_compare6445897_arg\, \$16612_compare6445898_arg\, 
                 \$16574_compare6445898_arg\, \$16916_compare6445898_arg\, 
                 \$15828_compare6445897_arg\, \$16881_compare6445898_arg\, 
                 \$15720_compare6445897_arg\, \$16951_compare6445898_arg\, 
                 \$15756_compare6445897_arg\, \$16811_compare6445898_arg\ : value(0 to 93) := (others => '0');
        variable \$13911\, \$13897\, \$13917\, \$13927_branch_if648_arg\ : value(0 to 122) := (others => '0');
        variable \$17547_copy_root_in_ram6635891_result\, \$16659_sp\, 
                 \$12840_next\, \$18665\, \$17330_sp\, 
                 \$18793_copy_root_in_ram6635879_result\, 
                 \$13105_copy_root_in_ram6635884_result\, 
                 \$18686_copy_root_in_ram6635880_result\, 
                 \$16662_fill6535928_result\, \$13921_loop665_result\, 
                 \$17105_w06555936_result\, 
                 \$12891_copy_root_in_ram6635884_result\, 
                 \$17520_copy_root_in_ram6635893_result\, \$17331_sp\, 
                 \$17492_next\, \$17459_loop665_result\, \$13472_next\, 
                 \$18664_next\, \$13078_copy_root_in_ram6635885_result\, 
                 \$18670_next\, \$17490_next\, \$18666_next\, \$17237_sp\, 
                 \$17734_copy_root_in_ram6635892_result\, 
                 \$17018_w36575938_result\, \$18633_loop665_result\, 
                 \$16650_sp\, \$17332_sp\, 
                 \$12864_copy_root_in_ram6635886_result\, \$16749_sp\, 
                 \$17009_sp\, \$12804_loop665_result\, 
                 \$12807_loop665_result\, \$17456_loop665_result\, 
                 \$16063_w6515922_result\, \$17000_sp\, 
                 \$17460_aux664_result\, \$16202_ofs\, 
                 \$12521_loop665_result\, \$18288_next\, \$16036_sp\, 
                 \$12838_next\, \$17491\, \$12844_next\, 
                 \$12680_loop665_result\, \$18634_aux664_result\, 
                 \$17012_sp\, \$17333_sp\, 
                 \$17761_copy_root_in_ram6635891_result\, \$18128_next\, 
                 \$14207_loop_push6495899_result\, \$17238_sp\, \$14181_sp\, 
                 \$17457_aux664_result\, \$12808_aux664_result\, 
                 \$12805_aux664_result\, \$12839\, \$13632_next\, 
                 \$16752_fill6545929_result\, \$19080_next\, \$17496_next\ : value(0 to 15) := (others => '0');
        variable \$12563\, \$12558\, \$12562\, \$12561\, \$v7438\, \$v7442\, 
                 \$v7450\, \$12560\, \$v7446\, \$12559\ : value(0 to 7) := (others => '0');
        variable \$14613_modulo6685896_arg\, \$15013_modulo6685896_arg\, 
                 \$15253_modulo6685896_arg\, \$14997_modulo6685888_arg\, 
                 \$15149_modulo6685895_arg\, \$14757_modulo6685888_arg\, 
                 \$14933_modulo6685896_arg\, \$15333_modulo6685896_arg\, 
                 \$15556_modulo6685895_arg\, \$15101_modulo6685888_arg\, 
                 \$14829_modulo6685895_arg\, \$15508_modulo6685888_arg\, 
                 \$15588_modulo6685888_arg\, \$15181_modulo6685888_arg\, 
                 \$14781_modulo6685888_arg\, \$15173_modulo6685896_arg\, 
                 \$15077_modulo6685888_arg\, \$15413_modulo6685896_arg\, 
                 \$14589_modulo6685895_arg\, \$14621_modulo6685888_arg\, 
                 \$14861_modulo6685888_arg\, \$15157_modulo6685888_arg\, 
                 \$15564_modulo6685888_arg\, \$14909_modulo6685895_arg\, 
                 \$15421_modulo6685888_arg\, \$15580_modulo6685896_arg\, 
                 \$14669_modulo6685895_arg\, \$15309_modulo6685895_arg\, 
                 \$14941_modulo6685888_arg\, \$14693_modulo6685896_arg\, 
                 \$15237_modulo6685888_arg\, \$15093_modulo6685896_arg\, 
                 \$15341_modulo6685888_arg\, \$15317_modulo6685888_arg\, 
                 \$14853_modulo6685896_arg\, \$14837_modulo6685888_arg\, 
                 \$15484_modulo6685888_arg\, \$15021_modulo6685888_arg\, 
                 \$15261_modulo6685888_arg\, \$15500_modulo6685896_arg\, 
                 \$14773_modulo6685896_arg\, \$15229_modulo6685895_arg\, 
                 \$15397_modulo6685888_arg\, \$14677_modulo6685888_arg\, 
                 \$15476_modulo6685895_arg\, \$14701_modulo6685888_arg\, 
                 \$14749_modulo6685895_arg\, \$15389_modulo6685895_arg\, 
                 \$14597_modulo6685888_arg\, \$14989_modulo6685895_arg\, 
                 \$14917_modulo6685888_arg\, \$15069_modulo6685895_arg\ : value(0 to 61) := (others => '0');
        variable \$13922_wait662_arg\, \$12681_wait662_arg\, 
                 \$12522_wait662_arg\ : value(0 to 96) := (others => '0');
        variable result5939 : value(0 to 57) := (others => '0');
        variable \$12539\, \$v6107\, \$12662\, \$v6106\, \$v6104\, \$v6103\, 
                 \$v6108\, \$v6105\ : value(0 to 3) := (others => '0');
        variable \$15508_modulo6685888_id\, \$13925_offsetclosure_n639_id\, 
                 \$15229_modulo6685895_id\, \$15013_modulo6685896_id\, 
                 \$15697_binop_compare6455918_id\, 
                 \$14207_loop_push6495899_id\, \$13923_make_block579_id\, 
                 \$17456_loop665_id\, \$15805_binop_compare6455921_id\, 
                 \$14884_binop_int6435904_id\, \$15564_modulo6685888_id\, 
                 \$15451_binop_int6435912_id\, \$15317_modulo6685888_id\, 
                 \$15588_modulo6685888_id\, \$16951_compare6445898_id\, 
                 \$15733_binop_compare6455919_id\, \$14941_modulo6685888_id\, 
                 \$14621_modulo6685888_id\, \$14853_modulo6685896_id\, 
                 \$15621_forever6705915_id\, \$15756_compare6445897_id\, 
                 \$16788_compbranch6505930_id\, \$14589_modulo6685895_id\, 
                 \$14781_modulo6685888_id\, \$14701_modulo6685888_id\, 
                 \$13924_apply638_id\, \$15309_modulo6685895_id\, 
                 \$15181_modulo6685888_id\, 
                 \$12891_copy_root_in_ram6635884_id\, 
                 \$15556_modulo6685895_id\, \$17459_loop665_id\, 
                 \$15500_modulo6685896_id\, \$15093_modulo6685896_id\, 
                 \$17048_w16565937_id\, \$13927_branch_if648_id\, 
                 \$16662_fill6535928_id\, \$16811_compare6445898_id\, 
                 \$18634_aux664_id\, \$17505_forever6705894_id\, 
                 \$12857_forever6705883_id\, \$15413_modulo6685896_id\, 
                 \$18632_loop666_id\, \$13105_copy_root_in_ram6635884_id\, 
                 \$15021_modulo6685888_id\, \$16752_fill6545929_id\, 
                 \$15684_compare6445897_id\, \$14597_modulo6685888_id\, 
                 \$14644_binop_int6435901_id\, \$16881_compare6445898_id\, 
                 \$15792_compare6445897_id\, \$16858_compbranch6505932_id\, 
                 \$12803_loop666_id\, \$15614_forever6705914_id\, 
                 \$14693_modulo6685896_id\, \$15397_modulo6685888_id\, 
                 \$12804_loop665_id\, \$15661_binop_compare6455917_id\, 
                 \$16612_compare6445898_id\, \$15149_modulo6685895_id\, 
                 \$18793_copy_root_in_ram6635879_id\, \$12522_wait662_id\, 
                 \$14989_modulo6685895_id\, \$15173_modulo6685896_id\, 
                 \$14804_binop_int6435903_id\, \$12681_wait662_id\, 
                 \$13928_w652_id\, \$17509_forever6705890_id\, 
                 \$15333_modulo6685896_id\, \$16986_compare6445898_id\, 
                 \$12853_forever6705887_id\, \$14861_modulo6685888_id\, 
                 \$13920_loop666_id\, \$14564_binop_int6435900_id\, 
                 \$17458_loop666_id\, \$15077_modulo6685888_id\, 
                 \$15447_forever6705911_id\, \$15157_modulo6685888_id\, 
                 \$17547_copy_root_in_ram6635891_id\, 
                 \$14909_modulo6685895_id\, \$13926_make_block_n646_id\, 
                 \$16846_compare6445898_id\, 
                 \$12864_copy_root_in_ram6635886_id\, 
                 \$14757_modulo6685888_id\, \$14773_modulo6685896_id\, 
                 \$15389_modulo6685895_id\, \$16928_compbranch6505934_id\, 
                 \$18686_copy_root_in_ram6635880_id\, \$16063_w6515922_id\, 
                 \$13922_wait662_id\, \$15101_modulo6685888_id\, 
                 \$16158_forever6705923_id\, \$14837_modulo6685888_id\, 
                 \$15364_binop_int6435910_id\, \$15284_binop_int6435909_id\, 
                 \$15531_binop_int6435913_id\, \$16195_forever6705924_id\, 
                 \$16916_compare6445898_id\, \$15421_modulo6685888_id\, 
                 \$14917_modulo6685888_id\, \$12806_loop666_id\, 
                 \$15253_modulo6685896_id\, \$15341_modulo6685888_id\, 
                 \$15580_modulo6685896_id\, \$15476_modulo6685895_id\, 
                 \$17761_copy_root_in_ram6635891_id\, 
                 \$16823_compbranch6505931_id\, 
                 \$15769_binop_compare6455920_id\, 
                 \$15828_compare6445897_id\, \$14669_modulo6685895_id\, 
                 \$13078_copy_root_in_ram6635885_id\, 
                 \$14613_modulo6685896_id\, \$15648_compare6445897_id\, 
                 \$14964_binop_int6435905_id\, \$17513_forever6705889_id\, 
                 \$15204_binop_int6435908_id\, \$17018_w36575938_id\, 
                 \$17520_copy_root_in_ram6635893_id\, 
                 \$15484_modulo6685888_id\, \$14933_modulo6685896_id\, 
                 \$14724_binop_int6435902_id\, \$14749_modulo6685895_id\, 
                 \$12679_loop666_id\, \$17105_w06555936_id\, 
                 \$15069_modulo6685895_id\, \$12807_loop665_id\, 
                 \$17460_aux664_id\, \$16510_forever6705925_id\, 
                 \$16589_compbranch6505927_id\, \$12808_aux664_id\, 
                 \$15720_compare6445897_id\, \$18679_forever6705881_id\, 
                 \$15237_modulo6685888_id\, \$14677_modulo6685888_id\, 
                 \$14829_modulo6685895_id\, \$15625_binop_compare6455916_id\, 
                 \$18633_loop665_id\, \$15124_binop_int6435907_id\, 
                 \$16551_compbranch6505926_id\, \$12520_loop666_id\, 
                 \$16963_compbranch6505935_id\, \$15044_binop_int6435906_id\, 
                 \$16574_compare6445898_id\, \$17455_loop666_id\, 
                 \$17734_copy_root_in_ram6635892_id\, 
                 \$15261_modulo6685888_id\, \$14997_modulo6685888_id\, 
                 \$16893_compbranch6505933_id\ : value(0 to 11) := (others => '0');
        variable \$16893_compbranch6505933_arg\, 
                 \$16928_compbranch6505934_arg\, 
                 \$16589_compbranch6505927_arg\, 
                 \$16551_compbranch6505926_arg\, 
                 \$16963_compbranch6505935_arg\, 
                 \$16823_compbranch6505931_arg\, 
                 \$16788_compbranch6505930_arg\, 
                 \$16858_compbranch6505932_arg\ : value(0 to 215) := (others => '0');
        variable \$14690_r\, \$14770_r\, \$14662_res\, \$15226_r\, 
                 \$14822_res\, \$15549_res\, \$17062\, \$15146_r\, 
                 \$14850_r\, \$15157_modulo6685888_result\, \$15066_r\, 
                 \$14586_r\, \$14742_res\, \$v7329\, \$15469_res\, 
                 \$15222_res\, \$15149_modulo6685895_result\, \$14906_r\, 
                 \$15090_r\, \$15473_r\, \$15093_modulo6685896_result\, 
                 \$13965\, \$15013_modulo6685896_result\, \$16998_argument3\, 
                 \$14982_res\, \$15069_modulo6685895_result\, 
                 \$16624_argument2\, \$14669_modulo6685895_result\, 
                 \$15851_argument1\, \$15142_res\, \$15062_res\, \$15410_r\, 
                 \$17207_arg\, \$15497_r\, \$14693_modulo6685896_result\, 
                 \$14917_modulo6685888_result\, \$15306_r\, 
                 \$15173_modulo6685896_result\, \$14826_r\, 
                 \$14853_modulo6685896_result\, 
                 \$15421_modulo6685888_result\, 
                 \$14997_modulo6685888_result\, \$15250_r\, 
                 \$15588_modulo6685888_result\, 
                 \$14773_modulo6685896_result\, \$15302_res\, \$15170_r\, 
                 \$14902_res\, \$14701_modulo6685888_result\, \$15577_r\, 
                 \$15564_modulo6685888_result\, 
                 \$14989_modulo6685895_result\, 
                 \$15229_modulo6685895_result\, \$16203\, 
                 \$15508_modulo6685888_result\, 
                 \$15500_modulo6685896_result\, 
                 \$14909_modulo6685895_result\, 
                 \$14941_modulo6685888_result\, 
                 \$15261_modulo6685888_result\, \$14610_r\, 
                 \$15580_modulo6685896_result\, 
                 \$14757_modulo6685888_result\, 
                 \$15253_modulo6685896_result\, 
                 \$14621_modulo6685888_result\, \$14930_r\, \$v7283\, 
                 \$15309_modulo6685895_result\, \$17165\, \$15382_res\, 
                 \$14677_modulo6685888_result\, 
                 \$15341_modulo6685888_result\, 
                 \$15556_modulo6685895_result\, \$14746_r\, 
                 \$15413_modulo6685896_result\, 
                 \$14829_modulo6685895_result\, \$15010_r\, 
                 \$14933_modulo6685896_result\, \$14986_r\, 
                 \$15181_modulo6685888_result\, 
                 \$15333_modulo6685896_result\, 
                 \$15101_modulo6685888_result\, 
                 \$15317_modulo6685888_result\, \$15386_r\, \$v7290\, 
                 \$15476_modulo6685895_result\, 
                 \$15021_modulo6685888_result\, \$14582_res\, 
                 \$14597_modulo6685888_result\, 
                 \$14837_modulo6685888_result\, 
                 \$15389_modulo6685895_result\, \$v7300\, 
                 \$15397_modulo6685888_result\, \$15330_r\, 
                 \$14861_modulo6685888_result\, 
                 \$14781_modulo6685888_result\, 
                 \$14613_modulo6685896_result\, 
                 \$15237_modulo6685888_result\, \$15553_r\, 
                 \$15484_modulo6685888_result\, \$v7313\, 
                 \$14749_modulo6685895_result\, 
                 \$15077_modulo6685888_result\, 
                 \$14589_modulo6685895_result\, \$14666_r\ : value(0 to 30) := (others => '0');
        variable \$13925_offsetclosure_n639_arg\ : value(0 to 137) := (others => '0');
        variable \$13923_make_block579_arg\ : value(0 to 103) := (others => '0');
        variable result6147, result5974, \$12523_make_block579_arg\, 
                 result6503, \$12682_make_block579_arg\ : value(0 to 127) := (others => '0');
        variable \$v6311\, \$v7071\, \$13537\, \$15751_res\, \$17784\, 
                 \$12718\, \$14368\, \$v6028\, \$12812\, \$13465\, \$v6349\, 
                 \$13690\, \$v5971\, \$17965\, \$v6010\, \$v6592\, \$v6932\, 
                 \$13020\, \$12690\, \$v7316\, \$13128\, \$v7209\, \$17236\, 
                 \$v7239\, \$v7053\, \$v6168\, \$17810\, \$v6120\, \$v6063\, 
                 \$v6636\, \$v7312\, \$14355\, \$13622\, \$v7063\, \$v7384\, 
                 \$v7124\, \$v6630\, \$12661\, \$v6687\, \$18656\, \$12876\, 
                 \$v6944\, \$13699\, \$v6674\, \$v6923\, \$v7225\, \$18477\, 
                 \$12850\, \$v7043\, \$16910_b\, \$v6929\, \$v7152\, 
                 \$13534\, \$v7286\, \$18469\, \$19056\, \$13230\, \$13305\, 
                 \$v6612\, \$17806\, \$17396\, \$v7319\, \$v6226\, \$v7065\, 
                 \$17161\, \$18923\, \$19137\, \$15444\, \$18422\, 
                 \$18632_loop666_result\, \$v7148\, \$18840\, \$18847\, 
                 \$14561\, \$v7073\, \$v7173\, \$12940\, \$v6777\, \$18700\, 
                 \$18347\, \$v7394\, \$v6615\, \$v7325\, \$13819\, \$v6483\, 
                 \$v5864\, \$12711\, \$v6310\, \$17601\, \$18282\, \$18920\, 
                 \$12721\, \$v6210\, \$16951_compare6445898_result\, 
                 \$12700\, \$v6877\, \$15446\, \$v6145\, \$v6086\, \$13391\, 
                 \$v6141\, \$17756\, \$17352\, \$v7052\, \$16358\, \$v6018\, 
                 \$17757\, \$17571\, \$13448\, \$18039\, \$v6977\, \$13014\, 
                 \$18349\, \$16980_b\, \$17811\, \$v6540\, \$18195\, 
                 \$14015\, \$19072\, \$19148\, \$17672\, \$v6871\, \$18817\, 
                 \$16846_compare6445898_result\, \$18914\, \$15643_res\, 
                 \$v7309\, \$14260\, \$17483\, \$v7055\, \$16357\, \$18350\, 
                 \$v7266\, \$v6793\, \$18471\, \$13130\, \$v6024\, \$13231\, 
                 \$v5877\, \$19000\, \$18468\, \$v7001\, \$16296\, \$16706\, 
                 \$19141\, \$16413\, \$17596\, \$15620\, \$19073\, \$v6006\, 
                 \$v5979\, \$18710\, \$v6808\, \$15611\, \$v6039\, \$13015\, 
                 \$13953\, \$13159\, \$16293\, \$13920_loop666_result\, 
                 \$v7106\, \$12693\, \$16155\, \$13152\, \$v6486\, \$v6191\, 
                 \$17680\, \$v7040\, \$v6770\, \$v6886\, \$v6051\, \$v6250\, 
                 \$v6418\, \$v6671\, \$v7430\, \$v6850\, \$19270\, \$13462\, 
                 \$v7341\, \$v6539\, \$13306\, \$v7390\, \$v7131\, \$v7410\, 
                 \$v6331\, \$17486\, \$v6339\, \$v5968\, \$v7136\, \$16658\, 
                 \$12831\, \$v6747\, \$v7407\, \$v6412\, \$17061\, \$12687\, 
                 \$v6556\, \$13952\, \$v6497\, \$v7160\, 
                 \$15720_compare6445897_result\, \$v6215\, \$17481\, 
                 \$v6124\, \$18573\, \$13024\, \$v7075\, \$v6698\, \$v7026\, 
                 \$15908\, \$v6076\, \$18042\, \$v7270\, rdy5975, \$v6260\, 
                 \$19074\, \$18672\, \$v6032\, \$13118\, \$v6663\, \$v7257\, 
                 \$v6983\, \$17353\, \$v6620\, 
                 \$15648_compare6445897_result\, \$v7024\, \$13951\, 
                 \$13119\, \$12742\, \$v6244\, \$12916\, \$14265\, \$16462\, 
                 \$13091\, \$v6647\, \$16157\, \$18728\, \$v7423\, \$v6576\, 
                 \$v6675\, \$v7080\, \$v6566\, \$13698\, \$v7105\, \$16322\, 
                 \$13958\, \$v5871\, \$19338\, \$13394\, \$17172\, \$v6290\, 
                 \$13821\, \$v6220\, \$17807\, \$v7226\, \$18671\, \$18736\, 
                 \$v7122\, \$18345\, \$13017\, \$17589\, 
                 \$16195_forever6705924_arg\, \$v6895\, \$v7347\, \$18353\, 
                 \$17884\, \$15621_forever6705915_arg\, \$v6079\, \$v6439\, 
                 \$v6571\, \$v6194\, \$v6345\, \$17542\, rdy6113, \$13314\, 
                 \$19147\, \$v5989\, \$v6926\, \$17534\, \$v6980\, \$17599\, 
                 \$13813\, \$18589\, \$17533\, \$v6755\, \$v7036\, \$19139\, 
                 \$13228\, \$17184\, \$v6448\, \$v6524\, \$16724\, \$v6083\, 
                 \$v6528\, \$v6720\, \$v6762\, \$13022\, \$v6811\, \$v6774\, 
                 \$16461\, \$18678\, \$13025\, \$v6477\, \$17465\, \$13386\, 
                 \$18658\, \$v6267\, \$12905\, \$19146\, \$v7303\, \$18839\, 
                 \$16916_compare6445898_result\, \$16193\, \$v7130\, 
                 \$12657\, \$v6691\, \$14342\, \$v6264\, \$v6600\, \$v6582\, 
                 \$17545\, \$v6361\, \$12845\, \$v6280\, \$17969\, \$16404\, 
                 \$17809\, \$v7134\, \$v7276\, \$12803_loop666_result\, 
                 \$17970\, \$v6820\, \$17808\, \$13150\, \$v6457\, \$17499\, 
                 \$12813\, \$v7282\, \$v7012\, \$17011\, \$19265\, \$v5982\, 
                 \$v6415\, \$v7082\, \$v6294\, \$13533\, \$13820\, \$13812\, 
                 \$17895\, \$v7111\, \$15684_compare6445897_result\, 
                 \$12832\, \$v6358\, \$12703\, \$v6059\, \$17166\, \$v6011\, 
                 \$v6111\, \$12659\, \$18924\, \$v6295\, \$18190\, \$v7060\, 
                 \$v6639\, \$v7084\, \$v5960\, result6112, \$v7032\, 
                 \$18344\, \$18992\, \$13315\, \$16515\, \$16156\, \$17560\, 
                 \$17010\, \$12846\, \$12674\, \$v6315\, \$v7031\, \$12547\, 
                 \$v7070\, \$14471\, \$18991\, \$18708\, \$16508\, \$v7242\, 
                 \$v6769\, \$v6735\, \$19271\, \$v5983\, \$v7033\, \$13815\, 
                 \$v5973\, \$v6603\, \$13018\, \$v6144\, \$v6259\, \$13147\, 
                 \$17503\, \$v6781\, \$v6054\, \$13232\, \$v7113\, \$v7233\, 
                 \$17786\, \$18040\, \$v6704\, \$17544\, \$v7114\, \$v6159\, 
                 \$13229\, \$v6332\, \$v6968\, \$v7041\, \$19002\, \$v7191\, 
                 \$16534\, \$13390\, \$19261\, \$v7103\, \$18047\, rdy6148, 
                 \$v7072\, \$v6187\, \$12708\, \$13239\, \$v6476\, \$v6002\, 
                 \$17894\, \$v6322\, \$v7419\, \$v6814\, \$v6156\, \$v7254\, 
                 \$13528\, \$18640\, \$12933\, \$v6140\, \$13963\, \$18638\, 
                 \$17748\, \$v6045\, \$17310\, \$v7120\, \$v6787\, \$17966\, 
                 \$v7096\, \$19264\, \$13311\, \$12744\, \$16133\, \$16232\, 
                 \$18351\, \$18262\, \$v6527\, \$16568_b\, \$16840_b\, 
                 \$14552\, \$13313\, \$v6905\, \$v6098\, \$13023\, \$v6511\, 
                 \$v7182\, \$12842\, \$13536\, \$18049\, \$v7176\, \$16194\, 
                 \$12719\, \$17758\, \$17973\, \$13939\, \$v7104\, \$17747\, 
                 \$12520_loop666_result\, \$v6796\, \$12811\, \$v6536\, 
                 \$16510_forever6705925_arg\, \$16473\, \$18281\, \$v7126\, 
                 \$18735\, \$v6253\, \$v7061\, \$17482\, \$13535\, \$19143\, 
                 \$v7102\, \$18122\, \$v6705\, \$16457\, \$13538\, \$v7457\, 
                 \$18922\, \$v6759\, \$17598\, \$17972\, \$18842\, \$18740\, 
                 \$17677\, \$13021\, \$12713\, \$v6531\, \$14069\, \$17388\, 
                 \$v5867\, \$v7051\, \$13624\, \$v7267\, \$v6650\, \$14148\, 
                 \$17675\, \$v7112\, \$13383\, \$v6433\, \$v7095\, \$17320\, 
                 \$v7014\, \$14051\, \$13464\, \$13236\, \$17395\, \$v7296\, 
                 \$v6784\, \$18674\, \$19136\, \$v6436\, \$13814\, \$v5947\, 
                 \$13539\, \$12743\, \$v6133\, \$v5972\, \$18046\, \$17504\, 
                 \$18993\, \$v6353\, \$v6263\, \$v7115\, \$18676\, \$v5876\, 
                 \$18844\, \$v7194\, \$v7289\, \$v7397\, \$v6394\, \$13695\, 
                 \$17497\, \$19242\, \$12814\, \$17814\, \$v6409\, \$13227\, 
                 \$17673\, \$16300\, \$v6752\, \$18196\, \$17347\, \$19260\, 
                 \$v6335\, \$16811_compare6445898_result\, \$14024\, 
                 \$v6666\, \$15679_res\, \$v6956\, \$v7083\, \$13691\, 
                 \$18921\, \$18326\, \$v6606\, \$14033\, \$v6219\, \$18051\, 
                 \$12889\, \$v6859\, \$12847\, \$v7101\, \$17008\, \$17595\, 
                 \$18918\, \$18737\, \$12760\, \$v6072\, \$18119\, \$v7197\, 
                 \$17314\, \$v6247\, \$17759\, \$16288\, \$13117\, \$12696\, 
                 \$12705\, \$17572\, \$14281\, \$v6844\, \$v7213\, \$12709\, 
                 \$17967\, \$13626\, \$16403\, \$15618\, \$v7273\, \$v7116\, 
                 \$16507\, \$v6917\, \$15619\, \$18191\, \$v6493\, \$13529\, 
                 \$v6243\, \$17532\, \$v7046\, \$v7449\, \$18564\, \$v7010\, 
                 \$15860\, \$13766\, \$18639\, \$v5998\, \$17968\, \$v5967\, 
                 \$15787_res\, \$19214\, \$18673\, \$17458_loop666_result\, 
                 \$v7427\, \$13688\, \$12706\, \$17032\, \$v6256\, \$v6588\, 
                 \$12934\, \$v6236\, \$v6550\, \$v6325\, \$v6714\, \$13092\, 
                 \$v5948\, \$17393\, \$v6283\, \$13158\, \$18998\, 
                 \$15715_res\, \$v6889\, \$v6180\, \$v7021\, \$v5964\, 
                 \$v6190\, \$17594\, \$12720\, \$18044\, \$v7350\, \$18994\, 
                 \$v6152\, \$v6643\, \$v7260\, \$19266\, 
                 \$17048_w16565937_result\, \$v6379\, \$v7056\, \$v6829\, 
                 \$v7011\, \$v6880\, \$v6938\, rdy6504, \$14273\, \$12829\, 
                 \$13309\, \$v6684\, \$v6352\, \$v6031\, \$v6075\, \$18913\, 
                 \$12710\, \$v6176\, \$v7093\, \$18668\, \$17592\, \$13385\, 
                 \$18048\, \$17883\, \$v7229\, \$v7459\, \$18572\, \$19268\, 
                 \$v7156\, \$v6899\, \$16336\, \$17173\, \$v7387\, \$v6223\, 
                 \$v6790\, \$v6137\, \$18660\, \$18669\, \$v6521\, \$13818\, 
                 \$15613\, \$13019\, \$17164\, \$13149\, \$12830\, \$v6623\, 
                 \$16440\, \$18478\, \$v6616\, \$19267\, \$v6354\, \$v7445\, 
                 \$v6442\, \$17243\, \$v6155\, \$v6908\, \$12717\, \$v7167\, 
                 \$17804\, \$16626\, \$18476\, \$v6902\, \$15909\, \$18470\, 
                 \$v6184\, \$v6547\, \$18041\, \$12942\, \$17502\, \$v6036\, 
                 \$v6660\, \$17066\, \$18732\, \$v6535\, \$v6553\, \$v6109\, 
                 \$v6093\, \$12688\, \$16509\, \$18738\, \$13316\, \$18841\, 
                 \$v6766\, \$v7393\, \$v5872\, \$v7081\, \$v7020\, \$18546\, 
                 \$v6965\, \$v6319\, \$v7044\, \$v6328\, \$14008\, \$18845\, 
                 \$v7375\, \$v6742\, \$v7378\, \$13463\, \$v7426\, \$v6743\, 
                 \$v6562\, \$v7188\, \$v6692\, \$v6646\, \$v7332\, \$v6758\, 
                 \$18473\, \$v6171\, \$v6373\, \$v5995\, \$15910\, \$v6835\, 
                 \$17513_forever6705889_arg\, \$v7100\, \$v6862\, \$13540\, 
                 \$18118\, \$v7110\, \$12704\, \$17671\, \$v6585\, \$v6543\, 
                 \$17892\, \$18184\, \$18730\, \$v6765\, \$v6832\, \$v7365\, 
                 \$13384\, \$v5986\, \$16321\, \$v6989\, \$v6920\, \$17964\, 
                 rdy6469, \$18189\, \$15447_forever6705911_arg\, \$v6717\, 
                 \$13234\, \$v6042\, \$v6654\, \$12701\, \$12694\, \$19118\, 
                 \$17561\, \$v6096\, \$v6069\, \$13101\, \$18348\, \$16317\, 
                 \$v7245\, \$18843\, \$13700\, \$12938\, \$18806\, \$v7135\, 
                 \$16382\, \$12903\, \$v6287\, \$13317\, \$18657\, \$v7433\, 
                 \$13940\, \$13510\, \$v6421\, \$17805\, \$17500\, \$v6424\, 
                 \$12735\, \$v6403\, \$13822\, \$v7203\, \$v6097\, \$13100\, 
                 \$v6463\, \$17815\, \$14296\, \$v7092\, \$v6799\, \$v6080\, 
                 \$v6563\, \$v6062\, \$v6817\, \$13817\, \$v6670\, \$12886\, 
                 \$v7364\, \$v6232\, \$13148\, \$18280\, \$v6546\, \$v7206\, 
                 \$v5999\, \$v6971\, \$14311\, \$17889\, \$v6207\, \$v6911\, 
                 \$v6066\, \$14381\, \$18043\, \$v6179\, \$v6110\, \$18995\, 
                 \$13689\, \$v6121\, \$v6579\, \$17466\, \$v6003\, \$v6898\, 
                 \$16986_compare6445898_result\, \$17593\, \$v6515\, 
                 \$v6992\, \$v6624\, \$18571\, \$v7210\, \$17812\, \$18193\, 
                 \$18194\, \$13129\, \$14135\, \$12716\, \$17785\, \$v6998\, 
                 \$18187\, \$17775\, \$v6724\, \$12736\, \$v7232\, \$12660\, 
                 \$12936\, \$15828_compare6445897_result\, \$17890\, 
                 \$18475\, \$12913\, \$v6388\, \$v6400\, \$v7091\, \$v7015\, 
                 \$16231\, \$17774\, \$v6089\, \$12695\, \$v7054\, \$18356\, 
                 \$v7328\, \$13694\, \$17254\, \$19070\, \$v6286\, \$13238\, 
                 \$v6847\, \$19262\, \$12914\, \$13794\, \$17783\, \$12941\, 
                 \$v6048\, \$18679_forever6705881_arg\, \$17495\, \$17590\, 
                 \$13387\, \$13393\, \$17348\, \$18677\, \$13389\, \$14254\, 
                 \$18185\, \$18472\, \$v6012\, \$v6162\, \$v7458\, 
                 \$17455_loop666_result\, \$v6595\, \$v6947\, \$v6314\, 
                 \$v5992\, \$v6183\, \$18711\, \$v5878\, \$v7076\, 
                 \$15792_compare6445897_result\, \$13312\, \$12702\, 
                 \$v6364\, \$v6678\, \$v6738\, \$v7030\, \$18104\, \$v6165\, 
                 \$16767\, \$16292\, \$v6751\, \$17463\, \$v7322\, \$13466\, 
                 \$v6853\, \$12904\, \$12734\, \$v6229\, \$13693\, \$v7185\, 
                 \$v5874\, \$v6301\, \$18637\, \$18999\, \$v7086\, \$v6773\, 
                 \$v7219\, \$12857_forever6705883_arg\, \$18836\, \$16031\, 
                 \$12878\, \$v7133\, \$16126\, \$17377\, 
                 \$13928_w652_result\, \$16035\, \$18166\, \$v7416\, 
                 \$12939\, \$14042\, \$13307\, \$17315\, \$13946\, \$18818\, 
                 \$v6175\, \$v7121\, \$v6865\, \$v6102\, \$v6609\, \$14558\, 
                 \$v7335\, \$v6950\, \$v7453\, \$v6701\, \$13153\, \$v6055\, 
                 \$18734\, \$12806_loop666_result\, \$v6681\, \$v6271\, 
                 \$v7358\, \$18479\, \$13692\, \$v7023\, \$13103\, \$v6268\, 
                 \$v6307\, \$v7016\, \$13957\, \$v6214\, \$17600\, \$v6657\, 
                 \$v6995\, \$12943\, \$v6117\, \$v7368\, \$v7064\, \$12843\, 
                 \$14161\, \$13962\, \$v7441\, \$v6962\, \$v6277\, \$v7455\, 
                 \$12741\, \$v6445\, \$17681\, \$17961\, \$16805_b\, 
                 \$v6986\, \$v6935\, \$v6750\, \$v7066\, \$v6007\, \$v7140\, 
                 \$16234\, \$12679_loop666_result\, \$17167\, \$12834\, 
                 \$16192\, \$17349\, \$13013\, \$18450\, \$v5951\, \$v5866\, 
                 \$v6203\, \$v6868\, \$14222\, \$13530\, \$v6709\, \$v7090\, 
                 \$v7004\, \$13127\, \$v7179\, \$15847\, \$16606_b\, 
                 \$v5954\, \$v6342\, \$v7299\, \$16165\, \$16078\, \$13941\, 
                 \$17319\, \$v7361\, \$v6688\, 
                 \$16612_compare6445898_result\, \$v6200\, \$v6367\, 
                 \$17962\, \$12691\, \$v7013\, \$v6651\, \$v7372\, \$v6574\, 
                 \$v6874\, \$16158_forever6705923_arg\, \$v6695\, \$17394\, 
                 \$v6826\, \$12887\, \$v7042\, \$v7164\, \$17885\, \$18816\, 
                 \$v7045\, \$19263\, \$16399\, \$v7248\, \$13623\, \$18570\, 
                 \$v6856\, \$v6710\, \$12848\, \$19071\, \$19140\, \$15612\, 
                 \$v6883\, \$16875_b\, \$17678\, \$v7034\, \$16677\, 
                 \$19144\, \$13890\, \$18915\, \$v6914\, \$v6729\, \$17387\, 
                 \$v6892\, \$v6492\, \$18045\, \$v6136\, \$12915\, \$v6627\, 
                 \$17591\, \$18699\, \$12715\, \$16365\, 
                 \$16574_compare6445898_result\, \$17354\, \$12945\, 
                 \$12712\, \$17674\, \$13157\, \$v6708\, \$18346\, 
                 \$16945_b\, \$17498\, \$19001\, \$v6274\, 
                 \$17509_forever6705890_arg\, \$v6739\, \$v7434\, \$13625\, 
                 \$12935\, \$12692\, \$v6304\, \$13016\, \$18120\, \$v7025\, 
                 \$18279\, \$v6953\, \$v5957\, \$18733\, \$v6838\, \$18925\, 
                 \$v6746\, \$v6941\, \$v7007\, \$17412\, \$19269\, \$17559\, 
                 \$v6239\, \$16353\, \$13395\, \$13823\, \$18709\, \$v6397\, 
                 \$v7035\, \$v7216\, \$v6172\, \$18188\, \$12851\, \$14431\, 
                 \$v6460\, \$v7279\, \$18186\, \$v6501\, \$12685\, \$18919\, 
                 \$v7293\, \$v6532\, \$v6291\, \$19142\, \$17803\, \$17963\, 
                 \$v6480\, \$13388\, \$17505_forever6705894_arg\, \$v6235\, 
                 \$14012\, \$13310\, \$18563\, \$14122\, \$v6058\, \$v6633\, 
                 \$16327\, \$13606\, \$18731\, \$v7085\, \$12544\, \$18278\, 
                 \$v6518\, \$v6298\, \$v6732\, 
                 \$16881_compare6445898_result\, \$12707\, \$v7074\, 
                 \$v7306\, \$17891\, \$v5944\, \$v5963\, \$13950\, \$17746\, 
                 \$v6596\, \$15874\, \$v6211\, \$13816\, \$v6591\, \$v6508\, 
                 \$v7413\, \$v6667\, \$v6489\, \$v6406\, \$15893\, \$19145\, 
                 \$17888\, \$v7200\, \$v7132\, \$v7406\, \$v6218\, 
                 \$15823_res\, \$v6780\, \$v7144\, \$18480\, \$18698\, 
                 \$12877\, \$18565\, \$v6559\, \$18815\, \$v6015\, \$13696\, 
                 \$17669\, \$v6318\, \$v6430\, \$v6599\, \$17464\, \$v6802\, 
                 \$14555\, \$17670\, \$13233\, \$v6376\, \$13235\, \$13102\, 
                 rdy5940, \$18355\, \$v6466\, \$13697\, \$v6021\, \$16115\, 
                 \$12937\, \$13155\, \$12888\, \$v7344\, \$17773\, \$12697\, 
                 \$v6146\, \$13237\, \$v7454\, \$v6496\, \$v5869\, \$v6500\, 
                 \$v6728\, \$17543\, \$18805\, \$18837\, \$v6027\, \$18807\, 
                 \$12689\, \$v7050\, \$v7338\, \$v6721\, \$v6823\, \$13532\, 
                 \$15756_compare6445897_result\, \$17597\, \$17484\, 
                 \$12714\, \$18739\, \$v6370\, \$v6502\, \$v7420\, \$13964\, 
                 \$18352\, \$v6336\, \$13154\, \$17679\, \$18916\, \$v6092\, 
                 \$18917\, \$18846\, \$v7381\, \$12944\, \$v6035\, \$12698\, 
                 \$17569\, \$v6805\, \$13151\, \$17886\, \$18474\, \$v6974\, 
                 \$16748\, \$v6427\, \$v6619\, \$v7371\, \$18655\, \$16271\, 
                 \$16233\, \$18050\, \$v7353\, \$15445\, \$17386\, \$v6240\, 
                 \$14326\, \$v6385\, \$17494\, \$v7251\, 
                 \$12853_forever6705887_arg\, \$v6382\, \$17121\, \$v6348\, 
                 \$17971\, \$13531\, \$v6959\, \$13824\, \$18838\, \$v6391\, 
                 \$v7094\, \$13945\, \$19138\, \$v6575\, \$13156\, \$16141\, 
                 \$v7236\, \$15614_forever6705914_arg\, \$v7170\, \$v6206\, 
                 \$13308\, \$v6512\, \$v7222\, \$18121\, \$17676\, \$17570\, 
                 \$v7437\, \$17893\, \$19003\, \$13090\, \$v7125\, \$12699\, 
                 \$v6567\, \$18835\, \$18997\, \$17887\, \$v6473\, \$12852\, 
                 \$v7062\, \$12545_x\, \$v6451\, \$18354\, \$16182\, 
                 \$v6725\, \$v6127\, \$13670\, \$18192\, \$18729\, \$v6642\, 
                 \$v7123\, \$19272\, \$v6197\, \$v7263\, \$v6130\, 
                 \$12673_rdy\, \$18996\, \$13392\, \$v7022\, \$v6841\, 
                 \$17813\, \$v6570\, \$v6454\, \$14060\ : value(0 to 0) := (others => '0');
        variable \$13926_make_block_n646_arg\ : value(0 to 171) := (others => '0');
        variable \$13924_apply638_arg\ : value(0 to 165) := (others => '0');
        variable \$18793_copy_root_in_ram6635879_arg\, 
                 \$18686_copy_root_in_ram6635880_arg\, 
                 \$13078_copy_root_in_ram6635885_arg\, 
                 \$17520_copy_root_in_ram6635893_arg\, \$12824\, 
                 \$16662_fill6535928_arg\, \$12681_wait662_result\, 
                 \$17547_copy_root_in_ram6635891_arg\, 
                 \$17761_copy_root_in_ram6635891_arg\, \$17476\, \$12737\, 
                 \$13105_copy_root_in_ram6635884_arg\, 
                 \$12864_copy_root_in_ram6635886_arg\, \$17389\, 
                 \$13922_wait662_result\, \$17048_w16565937_arg\, 
                 \$12522_wait662_result\, 
                 \$17734_copy_root_in_ram6635892_arg\, 
                 \$12891_copy_root_in_ram6635884_arg\, \$18566\, \$18650\, 
                 \$16752_fill6545929_arg\, \$17018_w36575938_arg\ : value(0 to 79) := (others => '0');
        variable \$17444\, \$18611\, \$18621\, \$17434\, \$12792\, \$12782\ : value(0 to 128) := (others => '0');
        variable \$15625_binop_compare6455916_arg\, \$16301\, 
                 \$15044_binop_int6435906_arg\, \$16383\, \$16337\, 
                 \$14724_binop_int6435902_arg\, \$16272\, 
                 \$14964_binop_int6435905_arg\, 
                 \$15451_binop_int6435912_arg\, 
                 \$14884_binop_int6435904_arg\, 
                 \$15364_binop_int6435910_arg\, 
                 \$15204_binop_int6435908_arg\, 
                 \$15284_binop_int6435909_arg\, 
                 \$14644_binop_int6435901_arg\, 
                 \$14804_binop_int6435903_arg\, 
                 \$15124_binop_int6435907_arg\, 
                 \$15733_binop_compare6455919_arg\, 
                 \$15805_binop_compare6455921_arg\, \$16441\, 
                 \$15697_binop_compare6455918_arg\, 
                 \$15769_binop_compare6455920_arg\, 
                 \$15661_binop_compare6455917_arg\, 
                 \$15531_binop_int6435913_arg\, \$14564_binop_int6435900_arg\ : value(0 to 153) := (others => '0');
        variable \$12654\, \$13374_w\, \$13628\, \$13093\, \$15465_v\, 
                 \$13803_w\, \$18340_hd\, \$16437_v\, \$14025_v\, \$v7087\, 
                 \$13120\, \$14493_v\, \$v7141\, \$14393_hd\, \$16041_v\, 
                 \$16335_v\, \$14002_v\, \$13889\, \$18545\, \$14081\, 
                 \$17660_w\, \$13987_v\, \$16313_v\, \$19132_hd\, 
                 \$17799_hd\, \$v7067\, \$15138_v\, \$18284\, \$14034_v\, 
                 \$18553\, \$16725\, \$16381_v\, \$14377_v\, \$16334_v\, 
                 \$19076\, \$13972_v\, \$13143_hd\, \$19111\, \$13684_hd\, 
                 \$17562\, \$17368_v\, \$18035_hd\, \$15747_v\, \$v7097\, 
                 \$15639_v\, \$v7149\, \$14103\, \$v7401\, \$v7037\, 
                 \$14464_v\, \$18180_hd\, \$13787\, \$v7157\, \$13977_v\, 
                 \$17952_w\, \$14185_next_env\, \$16380_v\, \$18030_w\, 
                 \$17183\, \$18261\, \$14300_v\, \$14512_v\, \$14898_v\, 
                 \$14016_v\, \$v7047\, \$16074_v\, \$16709\, \$v7127\, 
                 \$13004_w\, \$15711_v\, \$14423_v\, \$14413_v\, \$18459_w\, 
                 \$15545_v\, \$12929_hd\, \$13992_v\, \$18464_hd\, \$18701\, 
                 \$14446_v\, \$18808\, \$19127_w\, \$14578_v\, \$14043_v\, 
                 \$15819_v\, \$17117_v\, \$18335_w\, \$18175_w\, \$17874_w\, 
                 \$17585_hd\, \$13605\, \$14165\, \$14406_v\, \$19213\, 
                 \$14738_v\, \$14070_v\, \$16673_v\, \$16349_v\, \$12553\, 
                 \$14139\, \$17371_v\, \$15883\, \$v7107\, \$17749\, 
                 \$17239_v\, \$13524_hd\, \$13223_hd\, \$15861_v\, \$v7117\, 
                 \$16763_v\, \$17535\, \$14463_v\, \$15980_v\, \$14508_v\, 
                 \$18443\, \$17374_v\, \$18826_w\, \$17337\, \$14092\, 
                 \$13009_hd\, \$14152\, \$12879\, \$v7355\, \$13765\, 
                 \$v7399\, \$12549\, \$13379_hd\, \$18124\, \$14315_v\, 
                 \$18319\, \$v7145\, \$15897\, \$16121_v\, \$13808_hd\, 
                 \$14221\, \$12924_w\, \$17957_hd\, \$12906\, \$12546_dur\, 
                 \$19251_w\, \$19235\, \$13138_w\, \$17879_hd\, 
                 \$14453_next_acc\, \$17580_w\, \$16630\, \$18724_hd\, 
                 \$16217_hd\, \$15378_v\, \$12538_cy\, \$16379_v\, \$v7398\, 
                 \$14424_v\, \$v7057\, \$15981_v\, \$16395_v\, \$18904_w\, 
                 \$v7077\, \$14285_v\, \$14114\, \$16127_v\, \$14658_v\, 
                 \$v7354\, \$16436_v\, \$14517_v\, \$18982_w\, \$16439_v\, 
                 \$14338_v\, \$15976_v\, \$14818_v\, \$16042_v\, \$v7400\, 
                 \$13296_w\, \$13301_hd\, \$14330_v\, \$15853_v\, \$v7017\, 
                 \$17250_v\, \$16713_v\, \$17794_w\, \$13468\, \$18831_hd\, 
                 \$16438_v\, \$15218_v\, \$18909_hd\, \$15298_v\, \$16037_v\, 
                 \$15783_v\, \$14351_v\, \$14177_hd\, \$v7403\, \$15961\, 
                 \$18159\, \$17665_hd\, \$16169_v\, \$17776\, \$13519_w\, 
                 \$v7402\, \$15932\, \$13218_w\, \$13663\, \$13679_w\, 
                 \$v7027\, \$16284_v\, \$14364_v\, \$19337\, \$19256_hd\, 
                 \$13967_v\, \$v7161\, \$15058_v\, \$16729_v\, \$14061_v\, 
                 \$14978_v\, \$13997_v\, \$16299_v\, \$v7137\, \$16527_f0\, 
                 \$18987_hd\, \$18719_w\, \$13982_v\, \$16178_v\, \$v7153\, 
                 \$16453_v\, \$14126\, \$13503\, \$14052_v\, \$15675_v\, 
                 \$18421\, \$14516_v\ : value(0 to 31) := (others => '0');
        variable \$15364_binop_int6435910_result\, 
                 \$16551_compbranch6505926_result\, 
                 \$15733_binop_compare6455919_result\, 
                 \$16858_compbranch6505932_result\, 
                 \$15124_binop_int6435907_result\, 
                 \$14884_binop_int6435904_result\, 
                 \$15769_binop_compare6455920_result\, 
                 \$15531_binop_int6435913_result\, 
                 \$14964_binop_int6435905_result\, 
                 \$15805_binop_compare6455921_result\, 
                 \$15451_binop_int6435912_result\, 
                 \$16788_compbranch6505930_result\, 
                 \$16963_compbranch6505935_result\, 
                 \$16589_compbranch6505927_result\, 
                 \$13925_offsetclosure_n639_result\, 
                 \$15044_binop_int6435906_result\, \$13924_apply638_result\, 
                 \$13926_make_block_n646_result\, 
                 \$15661_binop_compare6455917_result\, 
                 \$15284_binop_int6435909_result\, 
                 \$14804_binop_int6435903_result\, 
                 \$15204_binop_int6435908_result\, 
                 \$16928_compbranch6505934_result\, 
                 \$16823_compbranch6505931_result\, 
                 \$15625_binop_compare6455916_result\, 
                 \$15697_binop_compare6455918_result\, result6468, 
                 \$14644_binop_int6435901_result\, 
                 \$13927_branch_if648_result\, 
                 \$16893_compbranch6505933_result\, 
                 \$14564_binop_int6435900_result\, 
                 \$14724_binop_int6435902_result\ : value(0 to 121) := (others => '0');
        variable state : t_state;
        variable state_var7464 : t_state_var7464;
        variable state_var7463 : t_state_var7463;
        variable state_var7462 : t_state_var7462;
        variable state_var7461 : t_state_var7461;
        variable state_var7460 : t_state_var7460;
        variable \$ram_lock\ : value(0 to 0);
        variable \$global_end_lock\ : value(0 to 0);
        variable \$code_lock\ : value(0 to 0);
        
    begin
      \$12559\ := \$12559%now\;
      \$14060\ := \$14060%now\;
      \$v6454\ := \$v6454%now\;
      \$14516_v\ := \$14516_v%now\;
      \$15069_modulo6685895_arg\ := \$15069_modulo6685895_arg%now\;
      \$18421\ := \$18421%now\;
      \$v6570\ := \$v6570%now\;
      \$14564_binop_int6435900_arg\ := \$14564_binop_int6435900_arg%now\;
      \$17813\ := \$17813%now\;
      \$v6841\ := \$v6841%now\;
      \$14666_r\ := \$14666_r%now\;
      \$v7022\ := \$v7022%now\;
      \$14589_modulo6685895_result\ := \$14589_modulo6685895_result%now\;
      \$13392\ := \$13392%now\;
      \$18996\ := \$18996%now\;
      \$12673_rdy\ := \$12673_rdy%now\;
      \$v6130\ := \$v6130%now\;
      \$v7263\ := \$v7263%now\;
      \$14917_modulo6685888_arg\ := \$14917_modulo6685888_arg%now\;
      \$v6197\ := \$v6197%now\;
      \$19272\ := \$19272%now\;
      \$v7123\ := \$v7123%now\;
      \$v6642\ := \$v6642%now\;
      \$18729\ := \$18729%now\;
      \$18192\ := \$18192%now\;
      \$13670\ := \$13670%now\;
      \$v6127\ := \$v6127%now\;
      \$15675_v\ := \$15675_v%now\;
      \$15077_modulo6685888_result\ := \$15077_modulo6685888_result%now\;
      \$v6725\ := \$v6725%now\;
      \$16182\ := \$16182%now\;
      \$14052_v\ := \$14052_v%now\;
      \$18354\ := \$18354%now\;
      \$14749_modulo6685895_result\ := \$14749_modulo6685895_result%now\;
      \$v6451\ := \$v6451%now\;
      \$12545_x\ := \$12545_x%now\;
      \$v7062\ := \$v7062%now\;
      \$17496_next\ := \$17496_next%now\;
      \$12852\ := \$12852%now\;
      \$13503\ := \$13503%now\;
      \$v6473\ := \$v6473%now\;
      \$15531_binop_int6435913_arg\ := \$15531_binop_int6435913_arg%now\;
      \$17887\ := \$17887%now\;
      \$18997\ := \$18997%now\;
      \$18835\ := \$18835%now\;
      \$v6567\ := \$v6567%now\;
      \$v7313\ := \$v7313%now\;
      \$14724_binop_int6435902_result\ := \$14724_binop_int6435902_result%now\;
      \$12699\ := \$12699%now\;
      \$v7125\ := \$v7125%now\;
      \$14989_modulo6685895_arg\ := \$14989_modulo6685895_arg%now\;
      \$13090\ := \$13090%now\;
      \$19003\ := \$19003%now\;
      \$12522_wait662_arg\ := \$12522_wait662_arg%now\;
      \$16811_compare6445898_arg\ := \$16811_compare6445898_arg%now\;
      \$17893\ := \$17893%now\;
      \$15661_binop_compare6455917_arg\ := \$15661_binop_compare6455917_arg%now\;
      \$14126\ := \$14126%now\;
      \$v7437\ := \$v7437%now\;
      \$17570\ := \$17570%now\;
      \$16453_v\ := \$16453_v%now\;
      \$17676\ := \$17676%now\;
      \$18121\ := \$18121%now\;
      \$v7222\ := \$v7222%now\;
      \$v6512\ := \$v6512%now\;
      \$13308\ := \$13308%now\;
      \$17018_w36575938_arg\ := \$17018_w36575938_arg%now\;
      \$v6206\ := \$v6206%now\;
      \$15484_modulo6685888_result\ := \$15484_modulo6685888_result%now\;
      \$v7170\ := \$v7170%now\;
      \$15614_forever6705914_arg\ := \$15614_forever6705914_arg%now\;
      \$16858_compbranch6505932_arg\ := \$16858_compbranch6505932_arg%now\;
      \$v7236\ := \$v7236%now\;
      \$v7153\ := \$v7153%now\;
      \$16893_compbranch6505933_id\ := \$16893_compbranch6505933_id%now\;
      \$14597_modulo6685888_arg\ := \$14597_modulo6685888_arg%now\;
      \$16141\ := \$16141%now\;
      \$v6105\ := \$v6105%now\;
      \$v7446\ := \$v7446%now\;
      \$13156\ := \$13156%now\;
      \$v6575\ := \$v6575%now\;
      \$19138\ := \$19138%now\;
      \$16178_v\ := \$16178_v%now\;
      \$13945\ := \$13945%now\;
      \$v7094\ := \$v7094%now\;
      \$v6391\ := \$v6391%now\;
      \$18838\ := \$18838%now\;
      \$13824\ := \$13824%now\;
      \$v6959\ := \$v6959%now\;
      \$13531\ := \$13531%now\;
      \$16788_compbranch6505930_arg\ := \$16788_compbranch6505930_arg%now\;
      \$17971\ := \$17971%now\;
      \$v6348\ := \$v6348%now\;
      \$17121\ := \$17121%now\;
      \$16752_fill6545929_arg\ := \$16752_fill6545929_arg%now\;
      \$v6382\ := \$v6382%now\;
      \$12853_forever6705887_arg\ := \$12853_forever6705887_arg%now\;
      \$v7251\ := \$v7251%now\;
      \$15769_binop_compare6455920_arg\ := \$15769_binop_compare6455920_arg%now\;
      \$17494\ := \$17494%now\;
      \$v6385\ := \$v6385%now\;
      \$14326\ := \$14326%now\;
      \$v6240\ := \$v6240%now\;
      \$19080_next\ := \$19080_next%now\;
      \$17386\ := \$17386%now\;
      \$13982_v\ := \$13982_v%now\;
      \$17459_loop665_arg\ := \$17459_loop665_arg%now\;
      \$18719_w\ := \$18719_w%now\;
      \$15445\ := \$15445%now\;
      \$v7353\ := \$v7353%now\;
      \$16752_fill6545929_result\ := \$16752_fill6545929_result%now\;
      \$14997_modulo6685888_id\ := \$14997_modulo6685888_id%now\;
      \$18050\ := \$18050%now\;
      \$12883\ := \$12883%now\;
      \$16823_compbranch6505931_arg\ := \$16823_compbranch6505931_arg%now\;
      \$16233\ := \$16233%now\;
      \$16271\ := \$16271%now\;
      \$12682_make_block579_arg\ := \$12682_make_block579_arg%now\;
      \$18655\ := \$18655%now\;
      \$v7371\ := \$v7371%now\;
      \$18987_hd\ := \$18987_hd%now\;
      \$v6619\ := \$v6619%now\;
      \$v6427\ := \$v6427%now\;
      \$16748\ := \$16748%now\;
      \$v6974\ := \$v6974%now\;
      \$18474\ := \$18474%now\;
      \$17886\ := \$17886%now\;
      \$15756_compare6445897_arg\ := \$15756_compare6445897_arg%now\;
      \$13151\ := \$13151%now\;
      \$v6805\ := \$v6805%now\;
      \$17569\ := \$17569%now\;
      \$12698\ := \$12698%now\;
      \$15389_modulo6685895_arg\ := \$15389_modulo6685895_arg%now\;
      \$v6035\ := \$v6035%now\;
      \$15553_r\ := \$15553_r%now\;
      \$15237_modulo6685888_result\ := \$15237_modulo6685888_result%now\;
      \$12944\ := \$12944%now\;
      \$14613_modulo6685896_result\ := \$14613_modulo6685896_result%now\;
      \$v7381\ := \$v7381%now\;
      \$18846\ := \$18846%now\;
      \$18917\ := \$18917%now\;
      \$v6092\ := \$v6092%now\;
      \$18916\ := \$18916%now\;
      \$15261_modulo6685888_id\ := \$15261_modulo6685888_id%now\;
      \$17679\ := \$17679%now\;
      \$13154\ := \$13154%now\;
      \$v6336\ := \$v6336%now\;
      \$16527_f0\ := \$16527_f0%now\;
      \$18352\ := \$18352%now\;
      \$13964\ := \$13964%now\;
      \$v7420\ := \$v7420%now\;
      \$13632_next\ := \$13632_next%now\;
      \$v6502\ := \$v6502%now\;
      \$v6370\ := \$v6370%now\;
      \$18739\ := \$18739%now\;
      \$12714\ := \$12714%now\;
      \$17484\ := \$17484%now\;
      \$17597\ := \$17597%now\;
      \$15756_compare6445897_result\ := \$15756_compare6445897_result%now\;
      \$v7137\ := \$v7137%now\;
      \$13532\ := \$13532%now\;
      \$v6823\ := \$v6823%now\;
      \$14781_modulo6685888_result\ := \$14781_modulo6685888_result%now\;
      \$v6721\ := \$v6721%now\;
      \$17734_copy_root_in_ram6635892_id\ := \$17734_copy_root_in_ram6635892_id%now\;
      \$v7338\ := \$v7338%now\;
      \$14749_modulo6685895_arg\ := \$14749_modulo6685895_arg%now\;
      \$v7050\ := \$v7050%now\;
      \$16299_v\ := \$16299_v%now\;
      \$12689\ := \$12689%now\;
      \$18807\ := \$18807%now\;
      \$13920_loop666_arg\ := \$13920_loop666_arg%now\;
      \$17455_loop666_id\ := \$17455_loop666_id%now\;
      \$v6027\ := \$v6027%now\;
      \$18650\ := \$18650%now\;
      \$18837\ := \$18837%now\;
      \$16951_compare6445898_arg\ := \$16951_compare6445898_arg%now\;
      \$14861_modulo6685888_result\ := \$14861_modulo6685888_result%now\;
      \$18805\ := \$18805%now\;
      \$17543\ := \$17543%now\;
      \$13997_v\ := \$13997_v%now\;
      \$16574_compare6445898_id\ := \$16574_compare6445898_id%now\;
      \$v6728\ := \$v6728%now\;
      \$v6500\ := \$v6500%now\;
      \$v5869\ := \$v5869%now\;
      \$v6496\ := \$v6496%now\;
      \$14978_v\ := \$14978_v%now\;
      \$v7454\ := \$v7454%now\;
      \$13237\ := \$13237%now\;
      \$v6146\ := \$v6146%now\;
      \$15330_r\ := \$15330_r%now\;
      \$12839\ := \$12839%now\;
      \$14061_v\ := \$14061_v%now\;
      \$14701_modulo6685888_arg\ := \$14701_modulo6685888_arg%now\;
      \$12697\ := \$12697%now\;
      \$17773\ := \$17773%now\;
      \$v7344\ := \$v7344%now\;
      \$12888\ := \$12888%now\;
      \$13155\ := \$13155%now\;
      \$12937\ := \$12937%now\;
      \$16115\ := \$16115%now\;
      \$12805_aux664_result\ := \$12805_aux664_result%now\;
      \$v6021\ := \$v6021%now\;
      \$13697\ := \$13697%now\;
      \$v6466\ := \$v6466%now\;
      \$18355\ := \$18355%now\;
      rdy5940 := \rdy5940%now\;
      \$13102\ := \$13102%now\;
      \$13235\ := \$13235%now\;
      \$15044_binop_int6435906_id\ := \$15044_binop_int6435906_id%now\;
      \$16729_v\ := \$16729_v%now\;
      \$v6376\ := \$v6376%now\;
      \$13233\ := \$13233%now\;
      \$17670\ := \$17670%now\;
      \$14555\ := \$14555%now\;
      \$14564_binop_int6435900_result\ := \$14564_binop_int6435900_result%now\;
      \$v6802\ := \$v6802%now\;
      \$15058_v\ := \$15058_v%now\;
      \$17464\ := \$17464%now\;
      \$v6599\ := \$v6599%now\;
      \$v6430\ := \$v6430%now\;
      \$v6318\ := \$v6318%now\;
      \$v7161\ := \$v7161%now\;
      \$17669\ := \$17669%now\;
      \$16963_compbranch6505935_id\ := \$16963_compbranch6505935_id%now\;
      \$13967_v\ := \$13967_v%now\;
      \$13696\ := \$13696%now\;
      \$v6015\ := \$v6015%now\;
      \$15476_modulo6685895_arg\ := \$15476_modulo6685895_arg%now\;
      \$17470\ := \$17470%now\;
      \$12520_loop666_id\ := \$12520_loop666_id%now\;
      \$18815\ := \$18815%now\;
      \$v6559\ := \$v6559%now\;
      \$18565\ := \$18565%now\;
      \$16551_compbranch6505926_id\ := \$16551_compbranch6505926_id%now\;
      \$15397_modulo6685888_result\ := \$15397_modulo6685888_result%now\;
      \$12877\ := \$12877%now\;
      \$18698\ := \$18698%now\;
      \$18480\ := \$18480%now\;
      \$v7300\ := \$v7300%now\;
      \$15389_modulo6685895_result\ := \$15389_modulo6685895_result%now\;
      \$v7144\ := \$v7144%now\;
      \$v6780\ := \$v6780%now\;
      \$19256_hd\ := \$19256_hd%now\;
      \$15823_res\ := \$15823_res%now\;
      \$15124_binop_int6435907_id\ := \$15124_binop_int6435907_id%now\;
      \$v6218\ := \$v6218%now\;
      \$v7406\ := \$v7406%now\;
      \$16963_compbranch6505935_arg\ := \$16963_compbranch6505935_arg%now\;
      \$v7132\ := \$v7132%now\;
      \$v7200\ := \$v7200%now\;
      \$18633_loop665_id\ := \$18633_loop665_id%now\;
      \$17888\ := \$17888%now\;
      \$19145\ := \$19145%now\;
      \$15625_binop_compare6455916_id\ := \$15625_binop_compare6455916_id%now\;
      \$19337\ := \$19337%now\;
      \$15893\ := \$15893%now\;
      \$14364_v\ := \$14364_v%now\;
      \$16893_compbranch6505933_result\ := \$16893_compbranch6505933_result%now\;
      \$v6406\ := \$v6406%now\;
      \$v6489\ := \$v6489%now\;
      \$14837_modulo6685888_result\ := \$14837_modulo6685888_result%now\;
      \$14677_modulo6685888_arg\ := \$14677_modulo6685888_arg%now\;
      \$v6667\ := \$v6667%now\;
      \$v7413\ := \$v7413%now\;
      \$v6508\ := \$v6508%now\;
      \$v6591\ := \$v6591%now\;
      \$16284_v\ := \$16284_v%now\;
      \$12808_aux664_result\ := \$12808_aux664_result%now\;
      \$13816\ := \$13816%now\;
      \$v6211\ := \$v6211%now\;
      \$15874\ := \$15874%now\;
      \$14829_modulo6685895_id\ := \$14829_modulo6685895_id%now\;
      \$v7027\ := \$v7027%now\;
      \$v6596\ := \$v6596%now\;
      \$17746\ := \$17746%now\;
      \$13950\ := \$13950%now\;
      \$v5963\ := \$v5963%now\;
      \$v5944\ := \$v5944%now\;
      \$14597_modulo6685888_result\ := \$14597_modulo6685888_result%now\;
      \$14582_res\ := \$14582_res%now\;
      \$17891\ := \$17891%now\;
      \$15397_modulo6685888_arg\ := \$15397_modulo6685888_arg%now\;
      \$13927_branch_if648_result\ := \$13927_branch_if648_result%now\;
      \$v7306\ := \$v7306%now\;
      \$v7074\ := \$v7074%now\;
      \$15021_modulo6685888_result\ := \$15021_modulo6685888_result%now\;
      \$12707\ := \$12707%now\;
      \$16881_compare6445898_result\ := \$16881_compare6445898_result%now\;
      \$13679_w\ := \$13679_w%now\;
      \$13663\ := \$13663%now\;
      \$18447\ := \$18447%now\;
      \$v6732\ := \$v6732%now\;
      \$v6298\ := \$v6298%now\;
      \$v6518\ := \$v6518%now\;
      \$18278\ := \$18278%now\;
      \$12544\ := \$12544%now\;
      \$13218_w\ := \$13218_w%now\;
      \$15932\ := \$15932%now\;
      \$v7402\ := \$v7402%now\;
      \$v7085\ := \$v7085%now\;
      \$18731\ := \$18731%now\;
      \$13519_w\ := \$13519_w%now\;
      \$13606\ := \$13606%now\;
      \$17776\ := \$17776%now\;
      \$18644\ := \$18644%now\;
      \$16327\ := \$16327%now\;
      \$16169_v\ := \$16169_v%now\;
      \$16551_compbranch6505926_arg\ := \$16551_compbranch6505926_arg%now\;
      \$15229_modulo6685895_arg\ := \$15229_modulo6685895_arg%now\;
      \$17457_aux664_result\ := \$17457_aux664_result%now\;
      \$v6633\ := \$v6633%now\;
      \$17665_hd\ := \$17665_hd%now\;
      \$18159\ := \$18159%now\;
      \$v6058\ := \$v6058%now\;
      \$14122\ := \$14122%now\;
      \$18563\ := \$18563%now\;
      \$13310\ := \$13310%now\;
      \$14012\ := \$14012%now\;
      \$14677_modulo6685888_id\ := \$14677_modulo6685888_id%now\;
      \$14181_sp\ := \$14181_sp%now\;
      \$v6235\ := \$v6235%now\;
      \$15961\ := \$15961%now\;
      \$15476_modulo6685895_result\ := \$15476_modulo6685895_result%now\;
      \$15237_modulo6685888_id\ := \$15237_modulo6685888_id%now\;
      \$17505_forever6705894_arg\ := \$17505_forever6705894_arg%now\;
      \$13388\ := \$13388%now\;
      \$v6480\ := \$v6480%now\;
      \$17001\ := \$17001%now\;
      \$17963\ := \$17963%now\;
      \$17803\ := \$17803%now\;
      \$19142\ := \$19142%now\;
      \$18679_forever6705881_id\ := \$18679_forever6705881_id%now\;
      \$v6291\ := \$v6291%now\;
      \$v6532\ := \$v6532%now\;
      \$v7293\ := \$v7293%now\;
      \$18919\ := \$18919%now\;
      \$12685\ := \$12685%now\;
      \$v6501\ := \$v6501%now\;
      \$17238_sp\ := \$17238_sp%now\;
      \$18186\ := \$18186%now\;
      \$v7279\ := \$v7279%now\;
      \$v6460\ := \$v6460%now\;
      \$14431\ := \$14431%now\;
      \$13667\ := \$13667%now\;
      \$17455_loop666_arg\ := \$17455_loop666_arg%now\;
      \$12851\ := \$12851%now\;
      \$18188\ := \$18188%now\;
      \$v6172\ := \$v6172%now\;
      \$v7403\ := \$v7403%now\;
      \$v7216\ := \$v7216%now\;
      \$v7035\ := \$v7035%now\;
      \$v6397\ := \$v6397%now\;
      \$18709\ := \$18709%now\;
      \$15720_compare6445897_id\ := \$15720_compare6445897_id%now\;
      \$13823\ := \$13823%now\;
      \$14177_hd\ := \$14177_hd%now\;
      result6503 := \result6503%now\;
      \$13395\ := \$13395%now\;
      \$16353\ := \$16353%now\;
      \$v6239\ := \$v6239%now\;
      \$17559\ := \$17559%now\;
      \$14351_v\ := \$14351_v%now\;
      \$12808_aux664_id\ := \$12808_aux664_id%now\;
      \$19269\ := \$19269%now\;
      \$17412\ := \$17412%now\;
      \$v7007\ := \$v7007%now\;
      \$v6941\ := \$v6941%now\;
      \$v6746\ := \$v6746%now\;
      \$18925\ := \$18925%now\;
      \$v6838\ := \$v6838%now\;
      \$18733\ := \$18733%now\;
      \$v5957\ := \$v5957%now\;
      \$v6953\ := \$v6953%now\;
      \$15783_v\ := \$15783_v%now\;
      \$18279\ := \$18279%now\;
      \$14207_loop_push6495899_result\ := \$14207_loop_push6495899_result%now\;
      \$v6108\ := \$v6108%now\;
      \$v7025\ := \$v7025%now\;
      \$18120\ := \$18120%now\;
      \$18566\ := \$18566%now\;
      \$13016\ := \$13016%now\;
      \$v6304\ := \$v6304%now\;
      \$12692\ := \$12692%now\;
      \$16037_v\ := \$16037_v%now\;
      \$12935\ := \$12935%now\;
      \$13625\ := \$13625%now\;
      \$v7434\ := \$v7434%now\;
      \$v6739\ := \$v6739%now\;
      \$17509_forever6705890_arg\ := \$17509_forever6705890_arg%now\;
      \$v6274\ := \$v6274%now\;
      \$19001\ := \$19001%now\;
      \$v7290\ := \$v7290%now\;
      \$17498\ := \$17498%now\;
      \$16945_b\ := \$16945_b%now\;
      \$15298_v\ := \$15298_v%now\;
      \$18346\ := \$18346%now\;
      \$16589_compbranch6505927_id\ := \$16589_compbranch6505927_id%now\;
      \$v6708\ := \$v6708%now\;
      \$13157\ := \$13157%now\;
      \$18909_hd\ := \$18909_hd%now\;
      \$17674\ := \$17674%now\;
      \$12712\ := \$12712%now\;
      \$12945\ := \$12945%now\;
      \$17354\ := \$17354%now\;
      \$16574_compare6445898_result\ := \$16574_compare6445898_result%now\;
      \$16365\ := \$16365%now\;
      \$12715\ := \$12715%now\;
      \$16510_forever6705925_id\ := \$16510_forever6705925_id%now\;
      \$15218_v\ := \$15218_v%now\;
      \$18699\ := \$18699%now\;
      \$17591\ := \$17591%now\;
      \$v6627\ := \$v6627%now\;
      \$12915\ := \$12915%now\;
      \$v6136\ := \$v6136%now\;
      \$18045\ := \$18045%now\;
      \$17460_aux664_id\ := \$17460_aux664_id%now\;
      \$12807_loop665_id\ := \$12807_loop665_id%now\;
      \$15069_modulo6685895_id\ := \$15069_modulo6685895_id%now\;
      \$v6492\ := \$v6492%now\;
      \$17487\ := \$17487%now\;
      \$v6892\ := \$v6892%now\;
      \$17387\ := \$17387%now\;
      \$15386_r\ := \$15386_r%now\;
      \$v6729\ := \$v6729%now\;
      \$v6914\ := \$v6914%now\;
      \$18915\ := \$18915%now\;
      \$17105_w06555936_id\ := \$17105_w06555936_id%now\;
      \$16589_compbranch6505927_arg\ := \$16589_compbranch6505927_arg%now\;
      \$13890\ := \$13890%now\;
      \$19144\ := \$19144%now\;
      \$16677\ := \$16677%now\;
      \$v7034\ := \$v7034%now\;
      \$17678\ := \$17678%now\;
      \$16875_b\ := \$16875_b%now\;
      \$13927_branch_if648_arg\ := \$13927_branch_if648_arg%now\;
      \$v6883\ := \$v6883%now\;
      \$16438_v\ := \$16438_v%now\;
      \$15612\ := \$15612%now\;
      \$14773_modulo6685896_arg\ := \$14773_modulo6685896_arg%now\;
      \$19140\ := \$19140%now\;
      \$19071\ := \$19071%now\;
      \$12848\ := \$12848%now\;
      \$18831_hd\ := \$18831_hd%now\;
      \$v6710\ := \$v6710%now\;
      \$13468\ := \$13468%now\;
      \$v6856\ := \$v6856%now\;
      \$15317_modulo6685888_result\ := \$15317_modulo6685888_result%now\;
      \$18570\ := \$18570%now\;
      \$13623\ := \$13623%now\;
      \$18128_next\ := \$18128_next%now\;
      \$v7248\ := \$v7248%now\;
      \$14644_binop_int6435901_result\ := \$14644_binop_int6435901_result%now\;
      \$12679_loop666_id\ := \$12679_loop666_id%now\;
      \$16399\ := \$16399%now\;
      \$19263\ := \$19263%now\;
      \$14749_modulo6685895_id\ := \$14749_modulo6685895_id%now\;
      \$17794_w\ := \$17794_w%now\;
      result6468 := \result6468%now\;
      \$v7045\ := \$v7045%now\;
      \$18816\ := \$18816%now\;
      \$17885\ := \$17885%now\;
      \$v7164\ := \$v7164%now\;
      \$15101_modulo6685888_result\ := \$15101_modulo6685888_result%now\;
      \$v7042\ := \$v7042%now\;
      \$15500_modulo6685896_arg\ := \$15500_modulo6685896_arg%now\;
      \$15333_modulo6685896_result\ := \$15333_modulo6685896_result%now\;
      \$17761_copy_root_in_ram6635891_result\ := \$17761_copy_root_in_ram6635891_result%now\;
      \$15720_compare6445897_arg\ := \$15720_compare6445897_arg%now\;
      \$16713_v\ := \$16713_v%now\;
      \$15697_binop_compare6455918_arg\ := \$15697_binop_compare6455918_arg%now\;
      \$17250_v\ := \$17250_v%now\;
      \$12887\ := \$12887%now\;
      \$v6826\ := \$v6826%now\;
      \$17394\ := \$17394%now\;
      \$v6695\ := \$v6695%now\;
      \$17333_sp\ := \$17333_sp%now\;
      \$v7017\ := \$v7017%now\;
      \$16158_forever6705923_arg\ := \$16158_forever6705923_arg%now\;
      \$v6874\ := \$v6874%now\;
      \$v6574\ := \$v6574%now\;
      \$15853_v\ := \$15853_v%now\;
      \$v7372\ := \$v7372%now\;
      \$v6651\ := \$v6651%now\;
      \$v7013\ := \$v7013%now\;
      \$15181_modulo6685888_result\ := \$15181_modulo6685888_result%now\;
      \$12691\ := \$12691%now\;
      \$17962\ := \$17962%now\;
      \$v6367\ := \$v6367%now\;
      \$v6200\ := \$v6200%now\;
      \$16612_compare6445898_result\ := \$16612_compare6445898_result%now\;
      \$v6688\ := \$v6688%now\;
      \$14330_v\ := \$14330_v%now\;
      \$v7361\ := \$v7361%now\;
      \$17319\ := \$17319%now\;
      \$13941\ := \$13941%now\;
      \$16078\ := \$16078%now\;
      \$16165\ := \$16165%now\;
      \$v7299\ := \$v7299%now\;
      \$17012_sp\ := \$17012_sp%now\;
      \$15261_modulo6685888_arg\ := \$15261_modulo6685888_arg%now\;
      \$v6342\ := \$v6342%now\;
      \$v5954\ := \$v5954%now\;
      \$16606_b\ := \$16606_b%now\;
      \$14986_r\ := \$14986_r%now\;
      \$13301_hd\ := \$13301_hd%now\;
      \$15847\ := \$15847%now\;
      \$v7179\ := \$v7179%now\;
      \$15021_modulo6685888_arg\ := \$15021_modulo6685888_arg%now\;
      \$13127\ := \$13127%now\;
      \$v7004\ := \$v7004%now\;
      \$v7090\ := \$v7090%now\;
      \$v6709\ := \$v6709%now\;
      \$17321\ := \$17321%now\;
      \$13530\ := \$13530%now\;
      \$14222\ := \$14222%now\;
      \$v6868\ := \$v6868%now\;
      \$v6203\ := \$v6203%now\;
      \$v5866\ := \$v5866%now\;
      \$v5951\ := \$v5951%now\;
      \$18450\ := \$18450%now\;
      \$13296_w\ := \$13296_w%now\;
      \$14724_binop_int6435902_id\ := \$14724_binop_int6435902_id%now\;
      \$v7400\ := \$v7400%now\;
      \$13013\ := \$13013%now\;
      \$17349\ := \$17349%now\;
      \$16192\ := \$16192%now\;
      \$12834\ := \$12834%now\;
      \$16441\ := \$16441%now\;
      \$17167\ := \$17167%now\;
      \$16042_v\ := \$16042_v%now\;
      \$15697_binop_compare6455918_result\ := \$15697_binop_compare6455918_result%now\;
      \$12679_loop666_result\ := \$12679_loop666_result%now\;
      \$16234\ := \$16234%now\;
      \$15625_binop_compare6455916_result\ := \$15625_binop_compare6455916_result%now\;
      \$v7140\ := \$v7140%now\;
      \$18163\ := \$18163%now\;
      \$v6007\ := \$v6007%now\;
      \$14933_modulo6685896_result\ := \$14933_modulo6685896_result%now\;
      \$v7066\ := \$v7066%now\;
      \$14818_v\ := \$14818_v%now\;
      \$v6750\ := \$v6750%now\;
      \$15976_v\ := \$15976_v%now\;
      \$v6935\ := \$v6935%now\;
      \$14338_v\ := \$14338_v%now\;
      \$v6986\ := \$v6986%now\;
      \$16805_b\ := \$16805_b%now\;
      \$17961\ := \$17961%now\;
      \$16439_v\ := \$16439_v%now\;
      \$14933_modulo6685896_id\ := \$14933_modulo6685896_id%now\;
      \$17681\ := \$17681%now\;
      \$12910\ := \$12910%now\;
      \$v6445\ := \$v6445%now\;
      \$12741\ := \$12741%now\;
      \$v7455\ := \$v7455%now\;
      \$v6277\ := \$v6277%now\;
      \$v6962\ := \$v6962%now\;
      \$v7441\ := \$v7441%now\;
      \$13962\ := \$13962%now\;
      \$15010_r\ := \$15010_r%now\;
      \$14829_modulo6685895_result\ := \$14829_modulo6685895_result%now\;
      \$12521_loop665_arg\ := \$12521_loop665_arg%now\;
      \$14161\ := \$14161%now\;
      \$15805_binop_compare6455921_arg\ := \$15805_binop_compare6455921_arg%now\;
      \$12843\ := \$12843%now\;
      \$15413_modulo6685896_result\ := \$15413_modulo6685896_result%now\;
      \$v7064\ := \$v7064%now\;
      \$15484_modulo6685888_arg\ := \$15484_modulo6685888_arg%now\;
      \$v7368\ := \$v7368%now\;
      \$v6117\ := \$v6117%now\;
      \$18634_aux664_result\ := \$18634_aux664_result%now\;
      \$12943\ := \$12943%now\;
      \$v6995\ := \$v6995%now\;
      \$v6657\ := \$v6657%now\;
      \$17600\ := \$17600%now\;
      \$v6214\ := \$v6214%now\;
      \$13957\ := \$13957%now\;
      \$v7016\ := \$v7016%now\;
      \$v6307\ := \$v6307%now\;
      \$v6268\ := \$v6268%now\;
      \$18982_w\ := \$18982_w%now\;
      \$13103\ := \$13103%now\;
      \$14517_v\ := \$14517_v%now\;
      \$v7023\ := \$v7023%now\;
      \$13692\ := \$13692%now\;
      \$18479\ := \$18479%now\;
      \$v7358\ := \$v7358%now\;
      \$v6271\ := \$v6271%now\;
      \$v6681\ := \$v6681%now\;
      \$12806_loop666_result\ := \$12806_loop666_result%now\;
      \$12680_loop665_result\ := \$12680_loop665_result%now\;
      \$18734\ := \$18734%now\;
      \$15484_modulo6685888_id\ := \$15484_modulo6685888_id%now\;
      \$v6055\ := \$v6055%now\;
      \$14746_r\ := \$14746_r%now\;
      \$17327\ := \$17327%now\;
      \$13153\ := \$13153%now\;
      \$v6701\ := \$v6701%now\;
      \$v7453\ := \$v7453%now\;
      \$v6950\ := \$v6950%now\;
      \$15733_binop_compare6455919_arg\ := \$15733_binop_compare6455919_arg%now\;
      \$16436_v\ := \$16436_v%now\;
      \$v7335\ := \$v7335%now\;
      \$14837_modulo6685888_arg\ := \$14837_modulo6685888_arg%now\;
      \$14558\ := \$14558%now\;
      \$v6609\ := \$v6609%now\;
      \$v6102\ := \$v6102%now\;
      \$v6865\ := \$v6865%now\;
      \$v7121\ := \$v7121%now\;
      \$v6175\ := \$v6175%now\;
      \$17520_copy_root_in_ram6635893_id\ := \$17520_copy_root_in_ram6635893_id%now\;
      \$18818\ := \$18818%now\;
      \$17018_w36575938_id\ := \$17018_w36575938_id%now\;
      \$13946\ := \$13946%now\;
      \$v7354\ := \$v7354%now\;
      \$17315\ := \$17315%now\;
      \$15204_binop_int6435908_id\ := \$15204_binop_int6435908_id%now\;
      \$14658_v\ := \$14658_v%now\;
      \$13307\ := \$13307%now\;
      \$14042\ := \$14042%now\;
      \$12939\ := \$12939%now\;
      \$12891_copy_root_in_ram6635884_arg\ := \$12891_copy_root_in_ram6635884_arg%now\;
      \$v7416\ := \$v7416%now\;
      \$18166\ := \$18166%now\;
      \$15556_modulo6685895_result\ := \$15556_modulo6685895_result%now\;
      \$16035\ := \$16035%now\;
      \$14853_modulo6685896_arg\ := \$14853_modulo6685896_arg%now\;
      \$15124_binop_int6435907_arg\ := \$15124_binop_int6435907_arg%now\;
      \$13928_w652_result\ := \$13928_w652_result%now\;
      \$15317_modulo6685888_arg\ := \$15317_modulo6685888_arg%now\;
      \$17377\ := \$17377%now\;
      \$16126\ := \$16126%now\;
      \$v7133\ := \$v7133%now\;
      \$16127_v\ := \$16127_v%now\;
      \$12878\ := \$12878%now\;
      \$16031\ := \$16031%now\;
      \$18836\ := \$18836%now\;
      \$12857_forever6705883_arg\ := \$12857_forever6705883_arg%now\;
      \$v7219\ := \$v7219%now\;
      \$v6773\ := \$v6773%now\;
      \$14114\ := \$14114%now\;
      \$v7086\ := \$v7086%now\;
      \$18999\ := \$18999%now\;
      \$18637\ := \$18637%now\;
      \$v6301\ := \$v6301%now\;
      \$17734_copy_root_in_ram6635892_arg\ := \$17734_copy_root_in_ram6635892_arg%now\;
      \$v5874\ := \$v5874%now\;
      \$v7185\ := \$v7185%now\;
      \$13693\ := \$13693%now\;
      \$v6229\ := \$v6229%now\;
      \$14285_v\ := \$14285_v%now\;
      \$12734\ := \$12734%now\;
      \$15341_modulo6685888_arg\ := \$15341_modulo6685888_arg%now\;
      \$12904\ := \$12904%now\;
      \$v7077\ := \$v7077%now\;
      \$17513_forever6705889_id\ := \$17513_forever6705889_id%now\;
      \$v6853\ := \$v6853%now\;
      \$13466\ := \$13466%now\;
      \$v7322\ := \$v7322%now\;
      \$14804_binop_int6435903_arg\ := \$14804_binop_int6435903_arg%now\;
      \$17463\ := \$17463%now\;
      \$19115\ := \$19115%now\;
      \$18904_w\ := \$18904_w%now\;
      \$12818\ := \$12818%now\;
      \$v6751\ := \$v6751%now\;
      \$16292\ := \$16292%now\;
      \$12844_next\ := \$12844_next%now\;
      \$16395_v\ := \$16395_v%now\;
      \$14964_binop_int6435905_id\ := \$14964_binop_int6435905_id%now\;
      \$16767\ := \$16767%now\;
      \$15093_modulo6685896_arg\ := \$15093_modulo6685896_arg%now\;
      \$v6103\ := \$v6103%now\;
      \$15648_compare6445897_id\ := \$15648_compare6445897_id%now\;
      \$v6165\ := \$v6165%now\;
      \$18104\ := \$18104%now\;
      \$v7030\ := \$v7030%now\;
      \$14613_modulo6685896_id\ := \$14613_modulo6685896_id%now\;
      \$v6738\ := \$v6738%now\;
      \$v6678\ := \$v6678%now\;
      \$17491\ := \$17491%now\;
      \$13078_copy_root_in_ram6635885_id\ := \$13078_copy_root_in_ram6635885_id%now\;
      \$15981_v\ := \$15981_v%now\;
      \$12560\ := \$12560%now\;
      \$v7057\ := \$v7057%now\;
      \$v6364\ := \$v6364%now\;
      \$12702\ := \$12702%now\;
      \$13312\ := \$13312%now\;
      \$12520_loop666_arg\ := \$12520_loop666_arg%now\;
      \$15792_compare6445897_result\ := \$15792_compare6445897_result%now\;
      \$15341_modulo6685888_result\ := \$15341_modulo6685888_result%now\;
      \$v7076\ := \$v7076%now\;
      \$14669_modulo6685895_id\ := \$14669_modulo6685895_id%now\;
      \$v5878\ := \$v5878%now\;
      \$18711\ := \$18711%now\;
      \$15828_compare6445897_id\ := \$15828_compare6445897_id%now\;
      \$15237_modulo6685888_arg\ := \$15237_modulo6685888_arg%now\;
      \$v6183\ := \$v6183%now\;
      \$v5992\ := \$v5992%now\;
      \$v6314\ := \$v6314%now\;
      \$12522_wait662_result\ := \$12522_wait662_result%now\;
      \$v6947\ := \$v6947%now\;
      \$v6595\ := \$v6595%now\;
      \$17455_loop666_result\ := \$17455_loop666_result%now\;
      \$v7458\ := \$v7458%now\;
      \$v6162\ := \$v6162%now\;
      \$12838_next\ := \$12838_next%now\;
      \$v6012\ := \$v6012%now\;
      \$18472\ := \$18472%now\;
      \$16036_sp\ := \$16036_sp%now\;
      \$18185\ := \$18185%now\;
      \$14424_v\ := \$14424_v%now\;
      \$14254\ := \$14254%now\;
      \$13389\ := \$13389%now\;
      \$18677\ := \$18677%now\;
      \$17348\ := \$17348%now\;
      \$13393\ := \$13393%now\;
      \$15769_binop_compare6455920_id\ := \$15769_binop_compare6455920_id%now\;
      \$13387\ := \$13387%now\;
      \$17590\ := \$17590%now\;
      \$v7398\ := \$v7398%now\;
      \$16823_compbranch6505931_id\ := \$16823_compbranch6505931_id%now\;
      \$17495\ := \$17495%now\;
      \$16379_v\ := \$16379_v%now\;
      \$16881_compare6445898_arg\ := \$16881_compare6445898_arg%now\;
      \$18679_forever6705881_arg\ := \$18679_forever6705881_arg%now\;
      \$v6048\ := \$v6048%now\;
      \$14677_modulo6685888_result\ := \$14677_modulo6685888_result%now\;
      \$18288_next\ := \$18288_next%now\;
      \$12538_cy\ := \$12538_cy%now\;
      \$15378_v\ := \$15378_v%now\;
      \$12941\ := \$12941%now\;
      \$17783\ := \$17783%now\;
      \$13794\ := \$13794%now\;
      \$14693_modulo6685896_arg\ := \$14693_modulo6685896_arg%now\;
      \$12914\ := \$12914%now\;
      \$19262\ := \$19262%now\;
      \$v6847\ := \$v6847%now\;
      \$15382_res\ := \$15382_res%now\;
      \$12521_loop665_result\ := \$12521_loop665_result%now\;
      \$13238\ := \$13238%now\;
      \$v6286\ := \$v6286%now\;
      \$19070\ := \$19070%now\;
      \$17254\ := \$17254%now\;
      \$13694\ := \$13694%now\;
      \$14941_modulo6685888_arg\ := \$14941_modulo6685888_arg%now\;
      \$v7328\ := \$v7328%now\;
      \$18356\ := \$18356%now\;
      \$v7054\ := \$v7054%now\;
      \$17761_copy_root_in_ram6635891_id\ := \$17761_copy_root_in_ram6635891_id%now\;
      \$12695\ := \$12695%now\;
      \$v6089\ := \$v6089%now\;
      \$17774\ := \$17774%now\;
      \$16231\ := \$16231%now\;
      \$v7015\ := \$v7015%now\;
      \$16202_ofs\ := \$16202_ofs%now\;
      \$v7091\ := \$v7091%now\;
      \$16217_hd\ := \$16217_hd%now\;
      \$v6400\ := \$v6400%now\;
      \$v6388\ := \$v6388%now\;
      \$16024\ := \$16024%now\;
      \$12913\ := \$12913%now\;
      \$17048_w16565937_arg\ := \$17048_w16565937_arg%now\;
      \$15476_modulo6685895_id\ := \$15476_modulo6685895_id%now\;
      \$16823_compbranch6505931_result\ := \$16823_compbranch6505931_result%now\;
      \$16928_compbranch6505934_result\ := \$16928_compbranch6505934_result%now\;
      \$18475\ := \$18475%now\;
      \$17890\ := \$17890%now\;
      \$15580_modulo6685896_id\ := \$15580_modulo6685896_id%now\;
      \$15828_compare6445897_result\ := \$15828_compare6445897_result%now\;
      \$12936\ := \$12936%now\;
      \$17165\ := \$17165%now\;
      \$12660\ := \$12660%now\;
      \$v7232\ := \$v7232%now\;
      \$12736\ := \$12736%now\;
      \$v6724\ := \$v6724%now\;
      \$18724_hd\ := \$18724_hd%now\;
      \$17775\ := \$17775%now\;
      \$16630\ := \$16630%now\;
      \$15341_modulo6685888_id\ := \$15341_modulo6685888_id%now\;
      \$18187\ := \$18187%now\;
      \$v6998\ := \$v6998%now\;
      \$17580_w\ := \$17580_w%now\;
      \$17785\ := \$17785%now\;
      \$12716\ := \$12716%now\;
      \$15253_modulo6685896_id\ := \$15253_modulo6685896_id%now\;
      \$14135\ := \$14135%now\;
      \$15828_compare6445897_arg\ := \$15828_compare6445897_arg%now\;
      \$13129\ := \$13129%now\;
      \$18194\ := \$18194%now\;
      \$18193\ := \$18193%now\;
      \$16916_compare6445898_arg\ := \$16916_compare6445898_arg%now\;
      \$17812\ := \$17812%now\;
      \$12806_loop666_id\ := \$12806_loop666_id%now\;
      \$15204_binop_int6435908_result\ := \$15204_binop_int6435908_result%now\;
      \$v7210\ := \$v7210%now\;
      \$17457_aux664_arg\ := \$17457_aux664_arg%now\;
      \$14453_next_acc\ := \$14453_next_acc%now\;
      \$18571\ := \$18571%now\;
      \$15309_modulo6685895_result\ := \$15309_modulo6685895_result%now\;
      \$17879_hd\ := \$17879_hd%now\;
      \$13138_w\ := \$13138_w%now\;
      \$v6624\ := \$v6624%now\;
      \$v6992\ := \$v6992%now\;
      \$14644_binop_int6435901_arg\ := \$14644_binop_int6435901_arg%now\;
      \$v6515\ := \$v6515%now\;
      \$13507\ := \$13507%now\;
      \$19235\ := \$19235%now\;
      \$17593\ := \$17593%now\;
      \$17460_aux664_result\ := \$17460_aux664_result%now\;
      \$v7283\ := \$v7283%now\;
      \$16986_compare6445898_result\ := \$16986_compare6445898_result%now\;
      \$14930_r\ := \$14930_r%now\;
      \$v6898\ := \$v6898%now\;
      \$v6003\ := \$v6003%now\;
      \$17466\ := \$17466%now\;
      \$v6579\ := \$v6579%now\;
      \$v6121\ := \$v6121%now\;
      \$14621_modulo6685888_result\ := \$14621_modulo6685888_result%now\;
      \$13689\ := \$13689%now\;
      \$14804_binop_int6435903_result\ := \$14804_binop_int6435903_result%now\;
      \$12782\ := \$12782%now\;
      \$18995\ := \$18995%now\;
      \$v6110\ := \$v6110%now\;
      \$v6179\ := \$v6179%now\;
      \$18043\ := \$18043%now\;
      \$19251_w\ := \$19251_w%now\;
      \$14381\ := \$14381%now\;
      \$v6066\ := \$v6066%now\;
      \$12546_dur\ := \$12546_dur%now\;
      \$v6911\ := \$v6911%now\;
      \$v6207\ := \$v6207%now\;
      \$15253_modulo6685896_result\ := \$15253_modulo6685896_result%now\;
      \$17889\ := \$17889%now\;
      \$14311\ := \$14311%now\;
      \$v6971\ := \$v6971%now\;
      \$v5999\ := \$v5999%now\;
      \$12906\ := \$12906%now\;
      \$v7206\ := \$v7206%now\;
      \$14917_modulo6685888_id\ := \$14917_modulo6685888_id%now\;
      \$18661\ := \$18661%now\;
      \$17957_hd\ := \$17957_hd%now\;
      \$12924_w\ := \$12924_w%now\;
      \$v6546\ := \$v6546%now\;
      \$18280\ := \$18280%now\;
      \$13148\ := \$13148%now\;
      \$v6232\ := \$v6232%now\;
      \$18633_loop665_arg\ := \$18633_loop665_arg%now\;
      \$14757_modulo6685888_result\ := \$14757_modulo6685888_result%now\;
      \$13922_wait662_result\ := \$13922_wait662_result%now\;
      \$v7364\ := \$v7364%now\;
      \$15580_modulo6685896_result\ := \$15580_modulo6685896_result%now\;
      \$15421_modulo6685888_id\ := \$15421_modulo6685888_id%now\;
      \$14610_r\ := \$14610_r%now\;
      \$16916_compare6445898_id\ := \$16916_compare6445898_id%now\;
      \$12886\ := \$12886%now\;
      \$16195_forever6705924_id\ := \$16195_forever6705924_id%now\;
      \$v6670\ := \$v6670%now\;
      \$13817\ := \$13817%now\;
      \$v6817\ := \$v6817%now\;
      \$14221\ := \$14221%now\;
      \$v6062\ := \$v6062%now\;
      \$17389\ := \$17389%now\;
      \$v6563\ := \$v6563%now\;
      \$v6080\ := \$v6080%now\;
      \$v6799\ := \$v6799%now\;
      \$v7092\ := \$v7092%now\;
      \$14296\ := \$14296%now\;
      \$17815\ := \$17815%now\;
      \$v6463\ := \$v6463%now\;
      \$13100\ := \$13100%now\;
      \$v6097\ := \$v6097%now\;
      \$v7203\ := \$v7203%now\;
      \$13808_hd\ := \$13808_hd%now\;
      \$13822\ := \$13822%now\;
      \$16121_v\ := \$16121_v%now\;
      \$v6403\ := \$v6403%now\;
      \$17000_sp\ := \$17000_sp%now\;
      \$12735\ := \$12735%now\;
      \$v6424\ := \$v6424%now\;
      \$15261_modulo6685888_result\ := \$15261_modulo6685888_result%now\;
      \$17500\ := \$17500%now\;
      \$17805\ := \$17805%now\;
      \$v6421\ := \$v6421%now\;
      \$13510\ := \$13510%now\;
      \$13940\ := \$13940%now\;
      \$v7433\ := \$v7433%now\;
      \$15309_modulo6685895_arg\ := \$15309_modulo6685895_arg%now\;
      \$18657\ := \$18657%now\;
      \$16574_compare6445898_arg\ := \$16574_compare6445898_arg%now\;
      \$13317\ := \$13317%now\;
      \$v6287\ := \$v6287%now\;
      \$12903\ := \$12903%now\;
      \$16382\ := \$16382%now\;
      \$15897\ := \$15897%now\;
      \$14941_modulo6685888_result\ := \$14941_modulo6685888_result%now\;
      \$14909_modulo6685895_result\ := \$14909_modulo6685895_result%now\;
      \$v7135\ := \$v7135%now\;
      \$18806\ := \$18806%now\;
      \$17458_loop666_arg\ := \$17458_loop666_arg%now\;
      \$12938\ := \$12938%now\;
      \$15531_binop_int6435913_id\ := \$15531_binop_int6435913_id%now\;
      \$15284_binop_int6435909_id\ := \$15284_binop_int6435909_id%now\;
      \$13700\ := \$13700%now\;
      \$18843\ := \$18843%now\;
      \$15364_binop_int6435910_id\ := \$15364_binop_int6435910_id%now\;
      \$12523_make_block579_arg\ := \$12523_make_block579_arg%now\;
      \$v7245\ := \$v7245%now\;
      \$16317\ := \$16317%now\;
      \$18348\ := \$18348%now\;
      \$13101\ := \$13101%now\;
      \$v6069\ := \$v6069%now\;
      \$16063_w6515922_result\ := \$16063_w6515922_result%now\;
      \$v6096\ := \$v6096%now\;
      \$12864_copy_root_in_ram6635886_arg\ := \$12864_copy_root_in_ram6635886_arg%now\;
      \$14669_modulo6685895_arg\ := \$14669_modulo6685895_arg%now\;
      \$17561\ := \$17561%now\;
      \$19118\ := \$19118%now\;
      \$14837_modulo6685888_id\ := \$14837_modulo6685888_id%now\;
      \$12694\ := \$12694%now\;
      \$15284_binop_int6435909_arg\ := \$15284_binop_int6435909_arg%now\;
      \$12701\ := \$12701%now\;
      \$v7450\ := \$v7450%now\;
      \$16158_forever6705923_id\ := \$16158_forever6705923_id%now\;
      \$15101_modulo6685888_id\ := \$15101_modulo6685888_id%now\;
      \$v7145\ := \$v7145%now\;
      \$v6654\ := \$v6654%now\;
      \$v6042\ := \$v6042%now\;
      \$13234\ := \$13234%now\;
      \$v6717\ := \$v6717%now\;
      \$15580_modulo6685896_arg\ := \$15580_modulo6685896_arg%now\;
      \$15500_modulo6685896_result\ := \$15500_modulo6685896_result%now\;
      \$15447_forever6705911_arg\ := \$15447_forever6705911_arg%now\;
      \$18189\ := \$18189%now\;
      rdy6469 := \rdy6469%now\;
      \$17964\ := \$17964%now\;
      \$18319\ := \$18319%now\;
      \$v6920\ := \$v6920%now\;
      \$v6989\ := \$v6989%now\;
      \$14315_v\ := \$14315_v%now\;
      \$18124\ := \$18124%now\;
      \$16321\ := \$16321%now\;
      \$v5986\ := \$v5986%now\;
      \$13384\ := \$13384%now\;
      \$13379_hd\ := \$13379_hd%now\;
      \$15421_modulo6685888_arg\ := \$15421_modulo6685888_arg%now\;
      \$v7365\ := \$v7365%now\;
      \$13922_wait662_id\ := \$13922_wait662_id%now\;
      \$12549\ := \$12549%now\;
      \$v6832\ := \$v6832%now\;
      \$v6765\ := \$v6765%now\;
      \$v6104\ := \$v6104%now\;
      \$18730\ := \$18730%now\;
      \$18184\ := \$18184%now\;
      \$17892\ := \$17892%now\;
      \$v6543\ := \$v6543%now\;
      \$v6585\ := \$v6585%now\;
      \$17671\ := \$17671%now\;
      \$v6106\ := \$v6106%now\;
      \$12704\ := \$12704%now\;
      \$v7399\ := \$v7399%now\;
      \$v7110\ := \$v7110%now\;
      \$18118\ := \$18118%now\;
      \$13540\ := \$13540%now\;
      \$v6862\ := \$v6862%now\;
      \$15508_modulo6685888_result\ := \$15508_modulo6685888_result%now\;
      \$v7100\ := \$v7100%now\;
      \$17513_forever6705889_arg\ := \$17513_forever6705889_arg%now\;
      \$v6835\ := \$v6835%now\;
      \$16203\ := \$16203%now\;
      \$15229_modulo6685895_result\ := \$15229_modulo6685895_result%now\;
      \$15910\ := \$15910%now\;
      \$17456_loop665_result\ := \$17456_loop665_result%now\;
      \$v5995\ := \$v5995%now\;
      \$13765\ := \$13765%now\;
      \$12807_loop665_result\ := \$12807_loop665_result%now\;
      \$v6373\ := \$v6373%now\;
      \$v6171\ := \$v6171%now\;
      \$18473\ := \$18473%now\;
      \$v6758\ := \$v6758%now\;
      \$v7332\ := \$v7332%now\;
      \$v6646\ := \$v6646%now\;
      \$v6692\ := \$v6692%now\;
      \$v7188\ := \$v7188%now\;
      \$16063_w6515922_id\ := \$16063_w6515922_id%now\;
      \$v6562\ := \$v6562%now\;
      \$v6743\ := \$v6743%now\;
      \$v7426\ := \$v7426%now\;
      \$13463\ := \$13463%now\;
      \$18686_copy_root_in_ram6635880_id\ := \$18686_copy_root_in_ram6635880_id%now\;
      \$v7378\ := \$v7378%now\;
      \$v6742\ := \$v6742%now\;
      \$14989_modulo6685895_result\ := \$14989_modulo6685895_result%now\;
      \$v7375\ := \$v7375%now\;
      \$15204_binop_int6435908_arg\ := \$15204_binop_int6435908_arg%now\;
      \$18845\ := \$18845%now\;
      \$14008\ := \$14008%now\;
      \$v6328\ := \$v6328%now\;
      \$v7355\ := \$v7355%now\;
      \$v7044\ := \$v7044%now\;
      \$v6319\ := \$v6319%now\;
      \$15364_binop_int6435910_arg\ := \$15364_binop_int6435910_arg%now\;
      \$v6965\ := \$v6965%now\;
      \$12879\ := \$12879%now\;
      \$15284_binop_int6435909_result\ := \$15284_binop_int6435909_result%now\;
      \$12804_loop665_result\ := \$12804_loop665_result%now\;
      \$18546\ := \$18546%now\;
      \$v7020\ := \$v7020%now\;
      \$15564_modulo6685888_result\ := \$15564_modulo6685888_result%now\;
      \$v7081\ := \$v7081%now\;
      \$v5872\ := \$v5872%now\;
      \$v7393\ := \$v7393%now\;
      \$14152\ := \$14152%now\;
      \$v6766\ := \$v6766%now\;
      \$18841\ := \$18841%now\;
      \$15661_binop_compare6455917_result\ := \$15661_binop_compare6455917_result%now\;
      \$13316\ := \$13316%now\;
      \$13009_hd\ := \$13009_hd%now\;
      \$14909_modulo6685895_arg\ := \$14909_modulo6685895_arg%now\;
      \$12682_make_block579_result\ := \$12682_make_block579_result%now\;
      \$18738\ := \$18738%now\;
      \$16509\ := \$16509%now\;
      \$12688\ := \$12688%now\;
      \$15577_r\ := \$15577_r%now\;
      \$v6093\ := \$v6093%now\;
      \$v6109\ := \$v6109%now\;
      \$15564_modulo6685888_arg\ := \$15564_modulo6685888_arg%now\;
      \$16928_compbranch6505934_id\ := \$16928_compbranch6505934_id%now\;
      \$14884_binop_int6435904_arg\ := \$14884_binop_int6435904_arg%now\;
      \$v6553\ := \$v6553%now\;
      \$14092\ := \$14092%now\;
      \$v6535\ := \$v6535%now\;
      \$18732\ := \$18732%now\;
      \$17066\ := \$17066%now\;
      \$15389_modulo6685895_id\ := \$15389_modulo6685895_id%now\;
      \$v6660\ := \$v6660%now\;
      \$17337\ := \$17337%now\;
      \$18826_w\ := \$18826_w%now\;
      \$v6036\ := \$v6036%now\;
      \$17374_v\ := \$17374_v%now\;
      \$17502\ := \$17502%now\;
      \$12942\ := \$12942%now\;
      \$14773_modulo6685896_id\ := \$14773_modulo6685896_id%now\;
      \$14757_modulo6685888_id\ := \$14757_modulo6685888_id%now\;
      \$18041\ := \$18041%now\;
      \$v6547\ := \$v6547%now\;
      \$v6184\ := \$v6184%now\;
      \$12864_copy_root_in_ram6635886_id\ := \$12864_copy_root_in_ram6635886_id%now\;
      \$18470\ := \$18470%now\;
      \$12835\ := \$12835%now\;
      \$15909\ := \$15909%now\;
      \$v6902\ := \$v6902%now\;
      \$17009_sp\ := \$17009_sp%now\;
      \$18476\ := \$18476%now\;
      \$16626\ := \$16626%now\;
      \$17804\ := \$17804%now\;
      \$18443\ := \$18443%now\;
      \$14701_modulo6685888_result\ := \$14701_modulo6685888_result%now\;
      \$v7167\ := \$v7167%now\;
      \$14902_res\ := \$14902_res%now\;
      \$12717\ := \$12717%now\;
      \$v6908\ := \$v6908%now\;
      \$13917\ := \$13917%now\;
      \$16749_sp\ := \$16749_sp%now\;
      \$v6155\ := \$v6155%now\;
      \$17243\ := \$17243%now\;
      \$v6442\ := \$v6442%now\;
      \$13923_make_block579_result\ := \$13923_make_block579_result%now\;
      \$v7445\ := \$v7445%now\;
      \$v6354\ := \$v6354%now\;
      \$14508_v\ := \$14508_v%now\;
      \$15157_modulo6685888_arg\ := \$15157_modulo6685888_arg%now\;
      \$19267\ := \$19267%now\;
      \$16846_compare6445898_id\ := \$16846_compare6445898_id%now\;
      \$15170_r\ := \$15170_r%now\;
      \$v6616\ := \$v6616%now\;
      \$13926_make_block_n646_id\ := \$13926_make_block_n646_id%now\;
      \$18478\ := \$18478%now\;
      \$16440\ := \$16440%now\;
      \$15451_binop_int6435912_arg\ := \$15451_binop_int6435912_arg%now\;
      \$15980_v\ := \$15980_v%now\;
      \$v6623\ := \$v6623%now\;
      \$14909_modulo6685895_id\ := \$14909_modulo6685895_id%now\;
      \$12830\ := \$12830%now\;
      \$13149\ := \$13149%now\;
      \$17164\ := \$17164%now\;
      \$14463_v\ := \$14463_v%now\;
      \$13019\ := \$13019%now\;
      \$15613\ := \$15613%now\;
      \$17535\ := \$17535%now\;
      \$13818\ := \$13818%now\;
      \$v6521\ := \$v6521%now\;
      \$16763_v\ := \$16763_v%now\;
      \$18669\ := \$18669%now\;
      \$18660\ := \$18660%now\;
      \$v6137\ := \$v6137%now\;
      \$v6790\ := \$v6790%now\;
      \$v7117\ := \$v7117%now\;
      \$v6223\ := \$v6223%now\;
      \$13105_copy_root_in_ram6635884_arg\ := \$13105_copy_root_in_ram6635884_arg%now\;
      \$v7387\ := \$v7387%now\;
      \$17547_copy_root_in_ram6635891_id\ := \$17547_copy_root_in_ram6635891_id%now\;
      \$15157_modulo6685888_id\ := \$15157_modulo6685888_id%now\;
      \$18632_loop666_arg\ := \$18632_loop666_arg%now\;
      \$17173\ := \$17173%now\;
      \$15447_forever6705911_id\ := \$15447_forever6705911_id%now\;
      \$15861_v\ := \$15861_v%now\;
      \$13223_hd\ := \$13223_hd%now\;
      \$13524_hd\ := \$13524_hd%now\;
      \$16336\ := \$16336%now\;
      \$v6899\ := \$v6899%now\;
      \$v7156\ := \$v7156%now\;
      \$15302_res\ := \$15302_res%now\;
      \$19268\ := \$19268%now\;
      \$18572\ := \$18572%now\;
      \$v7459\ := \$v7459%now\;
      \$v7229\ := \$v7229%now\;
      \$17883\ := \$17883%now\;
      \$18048\ := \$18048%now\;
      \$13385\ := \$13385%now\;
      \$17239_v\ := \$17239_v%now\;
      \$14773_modulo6685896_result\ := \$14773_modulo6685896_result%now\;
      \$17592\ := \$17592%now\;
      \$13926_make_block_n646_result\ := \$13926_make_block_n646_result%now\;
      \$17749\ := \$17749%now\;
      \$18668\ := \$18668%now\;
      \$v7093\ := \$v7093%now\;
      \$v6176\ := \$v6176%now\;
      \$12710\ := \$12710%now\;
      \$18913\ := \$18913%now\;
      \$v7107\ := \$v7107%now\;
      \$v6075\ := \$v6075%now\;
      \$v6031\ := \$v6031%now\;
      \$14861_modulo6685888_arg\ := \$14861_modulo6685888_arg%now\;
      \$v6352\ := \$v6352%now\;
      \$13924_apply638_result\ := \$13924_apply638_result%now\;
      \$15883\ := \$15883%now\;
      \$v6684\ := \$v6684%now\;
      \$13309\ := \$13309%now\;
      \$12829\ := \$12829%now\;
      \$14273\ := \$14273%now\;
      rdy6504 := \rdy6504%now\;
      \$v6938\ := \$v6938%now\;
      \$17371_v\ := \$17371_v%now\;
      \$v6880\ := \$v6880%now\;
      \$v7011\ := \$v7011%now\;
      \$17232\ := \$17232%now\;
      \$12864_copy_root_in_ram6635886_result\ := \$12864_copy_root_in_ram6635886_result%now\;
      \$v6829\ := \$v6829%now\;
      \$v7056\ := \$v7056%now\;
      \$14139\ := \$14139%now\;
      \$v6379\ := \$v6379%now\;
      \$17332_sp\ := \$17332_sp%now\;
      \$17048_w16565937_result\ := \$17048_w16565937_result%now\;
      \$19266\ := \$19266%now\;
      \$15588_modulo6685888_result\ := \$15588_modulo6685888_result%now\;
      \$v7260\ := \$v7260%now\;
      \$14621_modulo6685888_arg\ := \$14621_modulo6685888_arg%now\;
      \$13924_apply638_arg\ := \$13924_apply638_arg%now\;
      \$v6643\ := \$v6643%now\;
      \$v6152\ := \$v6152%now\;
      \$18994\ := \$18994%now\;
      \$15250_r\ := \$15250_r%now\;
      \$15044_binop_int6435906_result\ := \$15044_binop_int6435906_result%now\;
      \$16650_sp\ := \$16650_sp%now\;
      \$v7350\ := \$v7350%now\;
      \$18633_loop665_result\ := \$18633_loop665_result%now\;
      \$12553\ := \$12553%now\;
      \$18044\ := \$18044%now\;
      \$12720\ := \$12720%now\;
      \$17594\ := \$17594%now\;
      \$v6190\ := \$v6190%now\;
      \$v5964\ := \$v5964%now\;
      \$13926_make_block_n646_arg\ := \$13926_make_block_n646_arg%now\;
      \$15077_modulo6685888_id\ := \$15077_modulo6685888_id%now\;
      \$v7021\ := \$v7021%now\;
      \$17018_w36575938_result\ := \$17018_w36575938_result%now\;
      \$v6180\ := \$v6180%now\;
      \$v6889\ := \$v6889%now\;
      \$15715_res\ := \$15715_res%now\;
      \$16349_v\ := \$16349_v%now\;
      \$14964_binop_int6435905_arg\ := \$14964_binop_int6435905_arg%now\;
      \$18998\ := \$18998%now\;
      \$13158\ := \$13158%now\;
      \$v6283\ := \$v6283%now\;
      \$17393\ := \$17393%now\;
      \$v5948\ := \$v5948%now\;
      \$13092\ := \$13092%now\;
      \$v6714\ := \$v6714%now\;
      \$v6325\ := \$v6325%now\;
      \$14997_modulo6685888_result\ := \$14997_modulo6685888_result%now\;
      \$v6550\ := \$v6550%now\;
      \$v6236\ := \$v6236%now\;
      \$12934\ := \$12934%now\;
      \$v6588\ := \$v6588%now\;
      \$v6256\ := \$v6256%now\;
      \$17458_loop666_id\ := \$17458_loop666_id%now\;
      \$17032\ := \$17032%now\;
      \$12706\ := \$12706%now\;
      \$16673_v\ := \$16673_v%now\;
      \$13688\ := \$13688%now\;
      \$v7427\ := \$v7427%now\;
      \$17458_loop666_result\ := \$17458_loop666_result%now\;
      \$12681_wait662_arg\ := \$12681_wait662_arg%now\;
      \$18673\ := \$18673%now\;
      \$17324\ := \$17324%now\;
      \$14070_v\ := \$14070_v%now\;
      \$12737\ := \$12737%now\;
      \$19214\ := \$19214%now\;
      \$15787_res\ := \$15787_res%now\;
      \$14589_modulo6685895_arg\ := \$14589_modulo6685895_arg%now\;
      \$v5967\ := \$v5967%now\;
      \$17968\ := \$17968%now\;
      \$14738_v\ := \$14738_v%now\;
      \$v5998\ := \$v5998%now\;
      \$18639\ := \$18639%now\;
      \$13766\ := \$13766%now\;
      \$15413_modulo6685896_arg\ := \$15413_modulo6685896_arg%now\;
      \$15860\ := \$15860%now\;
      \$v7010\ := \$v7010%now\;
      \$18564\ := \$18564%now\;
      \$v7449\ := \$v7449%now\;
      \$v7046\ := \$v7046%now\;
      \$17532\ := \$17532%now\;
      \$v6243\ := \$v6243%now\;
      \$19213\ := \$19213%now\;
      \$13529\ := \$13529%now\;
      \$v6493\ := \$v6493%now\;
      \$15421_modulo6685888_result\ := \$15421_modulo6685888_result%now\;
      \$18191\ := \$18191%now\;
      \$14564_binop_int6435900_id\ := \$14564_binop_int6435900_id%now\;
      \$12679_loop666_arg\ := \$12679_loop666_arg%now\;
      \$14406_v\ := \$14406_v%now\;
      \$15619\ := \$15619%now\;
      \$v6917\ := \$v6917%now\;
      \$16507\ := \$16507%now\;
      \$v7116\ := \$v7116%now\;
      \$v7273\ := \$v7273%now\;
      \$14165\ := \$14165%now\;
      \$13920_loop666_id\ := \$13920_loop666_id%now\;
      \$15618\ := \$15618%now\;
      \$16403\ := \$16403%now\;
      \$17476\ := \$17476%now\;
      \$13626\ := \$13626%now\;
      \$17967\ := \$17967%now\;
      \$12709\ := \$12709%now\;
      \$v7213\ := \$v7213%now\;
      \$14861_modulo6685888_id\ := \$14861_modulo6685888_id%now\;
      \$v6844\ := \$v6844%now\;
      \$12804_loop665_arg\ := \$12804_loop665_arg%now\;
      \$14281\ := \$14281%now\;
      \$16272\ := \$16272%now\;
      \$17572\ := \$17572%now\;
      \$12705\ := \$12705%now\;
      \$12696\ := \$12696%now\;
      \$13117\ := \$13117%now\;
      \$13605\ := \$13605%now\;
      \$16288\ := \$16288%now\;
      \$12853_forever6705887_id\ := \$12853_forever6705887_id%now\;
      \$17734_copy_root_in_ram6635892_result\ := \$17734_copy_root_in_ram6635892_result%now\;
      \$17759\ := \$17759%now\;
      \$v6247\ := \$v6247%now\;
      \$16986_compare6445898_id\ := \$16986_compare6445898_id%now\;
      \$17314\ := \$17314%now\;
      \$v7197\ := \$v7197%now\;
      \$12680_loop665_arg\ := \$12680_loop665_arg%now\;
      \$18119\ := \$18119%now\;
      \$v6072\ := \$v6072%now\;
      \$12760\ := \$12760%now\;
      \$12548_dis\ := \$12548_dis%now\;
      \$15077_modulo6685888_arg\ := \$15077_modulo6685888_arg%now\;
      \$14853_modulo6685896_result\ := \$14853_modulo6685896_result%now\;
      \$18737\ := \$18737%now\;
      \$18918\ := \$18918%now\;
      \$17237_sp\ := \$17237_sp%now\;
      \$15173_modulo6685896_arg\ := \$15173_modulo6685896_arg%now\;
      \$17595\ := \$17595%now\;
      \$17008\ := \$17008%now\;
      \$17761_copy_root_in_ram6635891_arg\ := \$17761_copy_root_in_ram6635891_arg%now\;
      \$v7101\ := \$v7101%now\;
      \$12847\ := \$12847%now\;
      \$v6859\ := \$v6859%now\;
      \$12889\ := \$12889%now\;
      \$18051\ := \$18051%now\;
      \$v6219\ := \$v6219%now\;
      \$14826_r\ := \$14826_r%now\;
      \$14033\ := \$14033%now\;
      \$v6606\ := \$v6606%now\;
      \$18326\ := \$18326%now\;
      \$18921\ := \$18921%now\;
      \$13691\ := \$13691%now\;
      \$v7083\ := \$v7083%now\;
      \$v6956\ := \$v6956%now\;
      \$15679_res\ := \$15679_res%now\;
      \$v6666\ := \$v6666%now\;
      \$19239\ := \$19239%now\;
      \$14024\ := \$14024%now\;
      \$v7442\ := \$v7442%now\;
      \$16811_compare6445898_result\ := \$16811_compare6445898_result%now\;
      \$14781_modulo6685888_arg\ := \$14781_modulo6685888_arg%now\;
      \$v6335\ := \$v6335%now\;
      \$19260\ := \$19260%now\;
      \$17347\ := \$17347%now\;
      \$15333_modulo6685896_id\ := \$15333_modulo6685896_id%now\;
      \$18196\ := \$18196%now\;
      \$v6752\ := \$v6752%now\;
      \$16300\ := \$16300%now\;
      \$17673\ := \$17673%now\;
      \$13227\ := \$13227%now\;
      \$16612_compare6445898_arg\ := \$16612_compare6445898_arg%now\;
      \$13925_offsetclosure_n639_result\ := \$13925_offsetclosure_n639_result%now\;
      \$v6409\ := \$v6409%now\;
      \$17814\ := \$17814%now\;
      \$17585_hd\ := \$17585_hd%now\;
      \$17509_forever6705890_id\ := \$17509_forever6705890_id%now\;
      \$17566\ := \$17566%now\;
      \$12814\ := \$12814%now\;
      \$19242\ := \$19242%now\;
      \$17497\ := \$17497%now\;
      \$13695\ := \$13695%now\;
      \$v6394\ := \$v6394%now\;
      \$v7397\ := \$v7397%now\;
      \$v7289\ := \$v7289%now\;
      \$v7194\ := \$v7194%now\;
      \$17874_w\ := \$17874_w%now\;
      \$18844\ := \$18844%now\;
      \$15181_modulo6685888_arg\ := \$15181_modulo6685888_arg%now\;
      \$18175_w\ := \$18175_w%now\;
      \$v5876\ := \$v5876%now\;
      \$18676\ := \$18676%now\;
      \$17539\ := \$17539%now\;
      \$v7115\ := \$v7115%now\;
      \$v6263\ := \$v6263%now\;
      \$v6353\ := \$v6353%now\;
      \$18335_w\ := \$18335_w%now\;
      \$18993\ := \$18993%now\;
      \$13928_w652_id\ := \$13928_w652_id%now\;
      \$17504\ := \$17504%now\;
      \$18046\ := \$18046%now\;
      \$12670\ := \$12670%now\;
      \$v5972\ := \$v5972%now\;
      \$v6133\ := \$v6133%now\;
      \$12743\ := \$12743%now\;
      \$13539\ := \$13539%now\;
      \$v5947\ := \$v5947%now\;
      \$17117_v\ := \$17117_v%now\;
      \$15173_modulo6685896_result\ := \$15173_modulo6685896_result%now\;
      \$15819_v\ := \$15819_v%now\;
      \$17547_copy_root_in_ram6635891_arg\ := \$17547_copy_root_in_ram6635891_arg%now\;
      \$12681_wait662_id\ := \$12681_wait662_id%now\;
      \$14043_v\ := \$14043_v%now\;
      \$13814\ := \$13814%now\;
      \$12803_loop666_arg\ := \$12803_loop666_arg%now\;
      \$v6436\ := \$v6436%now\;
      \$19136\ := \$19136%now\;
      \$18674\ := \$18674%now\;
      \$v6784\ := \$v6784%now\;
      \$v7296\ := \$v7296%now\;
      \$17395\ := \$17395%now\;
      \$13236\ := \$13236%now\;
      \$13464\ := \$13464%now\;
      \$14051\ := \$14051%now\;
      \$v7014\ := \$v7014%now\;
      \$17320\ := \$17320%now\;
      \$v7095\ := \$v7095%now\;
      \$v6433\ := \$v6433%now\;
      \$12681_wait662_result\ := \$12681_wait662_result%now\;
      \$13383\ := \$13383%now\;
      \$14578_v\ := \$14578_v%now\;
      \$v7112\ := \$v7112%now\;
      \$17675\ := \$17675%now\;
      \$19127_w\ := \$19127_w%now\;
      \$18808\ := \$18808%now\;
      \$14148\ := \$14148%now\;
      \$18705\ := \$18705%now\;
      \$14804_binop_int6435903_id\ := \$14804_binop_int6435903_id%now\;
      \$v6650\ := \$v6650%now\;
      \$v7267\ := \$v7267%now\;
      \$13624\ := \$13624%now\;
      \$15588_modulo6685888_arg\ := \$15588_modulo6685888_arg%now\;
      \$v7051\ := \$v7051%now\;
      \$v5867\ := \$v5867%now\;
      \$17388\ := \$17388%now\;
      \$15173_modulo6685896_id\ := \$15173_modulo6685896_id%now\;
      \$16589_compbranch6505927_result\ := \$16589_compbranch6505927_result%now\;
      \$14069\ := \$14069%now\;
      \$v6531\ := \$v6531%now\;
      \$12713\ := \$12713%now\;
      \$13021\ := \$13021%now\;
      \$18666_next\ := \$18666_next%now\;
      \$14446_v\ := \$14446_v%now\;
      \$17677\ := \$17677%now\;
      \$18740\ := \$18740%now\;
      \$18842\ := \$18842%now\;
      \$17972\ := \$17972%now\;
      \$14989_modulo6685895_id\ := \$14989_modulo6685895_id%now\;
      \$17598\ := \$17598%now\;
      \$12522_wait662_id\ := \$12522_wait662_id%now\;
      \$18701\ := \$18701%now\;
      \$16662_fill6535928_arg\ := \$16662_fill6535928_arg%now\;
      \$17490_next\ := \$17490_next%now\;
      \$v6759\ := \$v6759%now\;
      \$16928_compbranch6505934_arg\ := \$16928_compbranch6505934_arg%now\;
      \$18922\ := \$18922%now\;
      \$18464_hd\ := \$18464_hd%now\;
      \$16963_compbranch6505935_result\ := \$16963_compbranch6505935_result%now\;
      \$13992_v\ := \$13992_v%now\;
      \$15508_modulo6685888_arg\ := \$15508_modulo6685888_arg%now\;
      \$12929_hd\ := \$12929_hd%now\;
      \$v7457\ := \$v7457%now\;
      \$13538\ := \$13538%now\;
      \$16457\ := \$16457%now\;
      \$15306_r\ := \$15306_r%now\;
      \$v6705\ := \$v6705%now\;
      \$18122\ := \$18122%now\;
      \$v7102\ := \$v7102%now\;
      \$19143\ := \$19143%now\;
      \$18670_next\ := \$18670_next%now\;
      \$18634_aux664_arg\ := \$18634_aux664_arg%now\;
      \$18793_copy_root_in_ram6635879_id\ := \$18793_copy_root_in_ram6635879_id%now\;
      \$15149_modulo6685895_id\ := \$15149_modulo6685895_id%now\;
      \$16788_compbranch6505930_result\ := \$16788_compbranch6505930_result%now\;
      \$13535\ := \$13535%now\;
      \$15545_v\ := \$15545_v%now\;
      \$17482\ := \$17482%now\;
      \$v7061\ := \$v7061%now\;
      \$v6253\ := \$v6253%now\;
      \$13897\ := \$13897%now\;
      \$18735\ := \$18735%now\;
      \$v7126\ := \$v7126%now\;
      \$18281\ := \$18281%now\;
      \$16473\ := \$16473%now\;
      \$14917_modulo6685888_result\ := \$14917_modulo6685888_result%now\;
      \$16741\ := \$16741%now\;
      \$16510_forever6705925_arg\ := \$16510_forever6705925_arg%now\;
      \$v6536\ := \$v6536%now\;
      \$12811\ := \$12811%now\;
      \$v6796\ := \$v6796%now\;
      \$18459_w\ := \$18459_w%now\;
      \$14413_v\ := \$14413_v%now\;
      \$12520_loop666_result\ := \$12520_loop666_result%now\;
      \$16612_compare6445898_id\ := \$16612_compare6445898_id%now\;
      \$17747\ := \$17747%now\;
      \$v7104\ := \$v7104%now\;
      \$13939\ := \$13939%now\;
      \$15661_binop_compare6455917_id\ := \$15661_binop_compare6455917_id%now\;
      \$17973\ := \$17973%now\;
      \$12804_loop665_id\ := \$12804_loop665_id%now\;
      \$17758\ := \$17758%now\;
      \$12719\ := \$12719%now\;
      \$15397_modulo6685888_id\ := \$15397_modulo6685888_id%now\;
      \$17105_w06555936_arg\ := \$17105_w06555936_arg%now\;
      \$12792\ := \$12792%now\;
      \$16194\ := \$16194%now\;
      \$v7176\ := \$v7176%now\;
      \$14829_modulo6685895_arg\ := \$14829_modulo6685895_arg%now\;
      \$18049\ := \$18049%now\;
      \$13536\ := \$13536%now\;
      \$12842\ := \$12842%now\;
      \$v7182\ := \$v7182%now\;
      \$v6511\ := \$v6511%now\;
      \$14693_modulo6685896_id\ := \$14693_modulo6685896_id%now\;
      \$13023\ := \$13023%now\;
      \$v6098\ := \$v6098%now\;
      \$15792_compare6445897_arg\ := \$15792_compare6445897_arg%now\;
      \$v6905\ := \$v6905%now\;
      \$13313\ := \$13313%now\;
      \$14552\ := \$14552%now\;
      \$16840_b\ := \$16840_b%now\;
      \$16568_b\ := \$16568_b%now\;
      \$14423_v\ := \$14423_v%now\;
      \$v6527\ := \$v6527%now\;
      \$18262\ := \$18262%now\;
      \$13078_copy_root_in_ram6635885_result\ := \$13078_copy_root_in_ram6635885_result%now\;
      \$18351\ := \$18351%now\;
      \$16232\ := \$16232%now\;
      \$16133\ := \$16133%now\;
      \$15711_v\ := \$15711_v%now\;
      \$15614_forever6705914_id\ := \$15614_forever6705914_id%now\;
      \$13004_w\ := \$13004_w%now\;
      \$12803_loop666_id\ := \$12803_loop666_id%now\;
      \$12744\ := \$12744%now\;
      \$13311\ := \$13311%now\;
      \$18664_next\ := \$18664_next%now\;
      \$19264\ := \$19264%now\;
      \$13472_next\ := \$13472_next%now\;
      \$16858_compbranch6505932_id\ := \$16858_compbranch6505932_id%now\;
      \$v7096\ := \$v7096%now\;
      \$17966\ := \$17966%now\;
      \$v6787\ := \$v6787%now\;
      \$17459_loop665_result\ := \$17459_loop665_result%now\;
      \$v7120\ := \$v7120%now\;
      \$17310\ := \$17310%now\;
      \$17492_next\ := \$17492_next%now\;
      \$v6045\ := \$v6045%now\;
      \$17748\ := \$17748%now\;
      \$18638\ := \$18638%now\;
      \$15792_compare6445897_id\ := \$15792_compare6445897_id%now\;
      \$13963\ := \$13963%now\;
      \$v6140\ := \$v6140%now\;
      \$12933\ := \$12933%now\;
      \$18640\ := \$18640%now\;
      \$13528\ := \$13528%now\;
      \$v7254\ := \$v7254%now\;
      \$16881_compare6445898_id\ := \$16881_compare6445898_id%now\;
      \$17460_aux664_arg\ := \$17460_aux664_arg%now\;
      \$12523_make_block579_result\ := \$12523_make_block579_result%now\;
      \$13922_wait662_arg\ := \$13922_wait662_arg%now\;
      \$v6156\ := \$v6156%now\;
      \$v6814\ := \$v6814%now\;
      \$v7419\ := \$v7419%now\;
      \$15451_binop_int6435912_result\ := \$15451_binop_int6435912_result%now\;
      \$v6322\ := \$v6322%now\;
      \$17331_sp\ := \$17331_sp%now\;
      \$17894\ := \$17894%now\;
      \$v6002\ := \$v6002%now\;
      \$v6476\ := \$v6476%now\;
      \$13239\ := \$13239%now\;
      \$12708\ := \$12708%now\;
      \$18812\ := \$18812%now\;
      \$v6187\ := \$v6187%now\;
      \$v7072\ := \$v7072%now\;
      rdy6148 := \rdy6148%now\;
      \$18047\ := \$18047%now\;
      \$14644_binop_int6435901_id\ := \$14644_binop_int6435901_id%now\;
      \$14597_modulo6685888_id\ := \$14597_modulo6685888_id%now\;
      \$v7103\ := \$v7103%now\;
      \$19261\ := \$19261%now\;
      \$16893_compbranch6505933_arg\ := \$16893_compbranch6505933_arg%now\;
      \$13390\ := \$13390%now\;
      \$16534\ := \$16534%now\;
      \$v7191\ := \$v7191%now\;
      \$19002\ := \$19002%now\;
      \$v7041\ := \$v7041%now\;
      \$v6968\ := \$v6968%now\;
      \$v7127\ := \$v7127%now\;
      \$17520_copy_root_in_ram6635893_result\ := \$17520_copy_root_in_ram6635893_result%now\;
      \$v6332\ := \$v6332%now\;
      \$13229\ := \$13229%now\;
      \$v6159\ := \$v6159%now\;
      \$15684_compare6445897_id\ := \$15684_compare6445897_id%now\;
      \$v7114\ := \$v7114%now\;
      \$17544\ := \$17544%now\;
      \$v6704\ := \$v6704%now\;
      \$18040\ := \$18040%now\;
      \$17786\ := \$17786%now\;
      \$v7233\ := \$v7233%now\;
      \$14207_loop_push6495899_arg\ := \$14207_loop_push6495899_arg%now\;
      \$16709\ := \$16709%now\;
      \$v7113\ := \$v7113%now\;
      \$14724_binop_int6435902_arg\ := \$14724_binop_int6435902_arg%now\;
      \$13232\ := \$13232%now\;
      \$16986_compare6445898_arg\ := \$16986_compare6445898_arg%now\;
      \$v6054\ := \$v6054%now\;
      \$16074_v\ := \$16074_v%now\;
      \$v6781\ := \$v6781%now\;
      \$v7047\ := \$v7047%now\;
      \$17503\ := \$17503%now\;
      \$13147\ := \$13147%now\;
      \$v6259\ := \$v6259%now\;
      \$v6144\ := \$v6144%now\;
      \$13018\ := \$13018%now\;
      \$v6603\ := \$v6603%now\;
      \$14016_v\ := \$14016_v%now\;
      \$16752_fill6545929_id\ := \$16752_fill6545929_id%now\;
      \$v5973\ := \$v5973%now\;
      \$13815\ := \$13815%now\;
      \$v7033\ := \$v7033%now\;
      \$v5983\ := \$v5983%now\;
      \$19271\ := \$19271%now\;
      \$v6735\ := \$v6735%now\;
      \$v6769\ := \$v6769%now\;
      \$v7242\ := \$v7242%now\;
      \$16508\ := \$16508%now\;
      \$12808_aux664_arg\ := \$12808_aux664_arg%now\;
      \$18708\ := \$18708%now\;
      \$18991\ := \$18991%now\;
      \$14471\ := \$14471%now\;
      \$v7070\ := \$v7070%now\;
      \$12547\ := \$12547%now\;
      \$v7031\ := \$v7031%now\;
      \$v6315\ := \$v6315%now\;
      \$12674\ := \$12674%now\;
      \$12846\ := \$12846%now\;
      \$17010\ := \$17010%now\;
      \$17560\ := \$17560%now\;
      \$16156\ := \$16156%now\;
      \$15021_modulo6685888_id\ := \$15021_modulo6685888_id%now\;
      \$13925_offsetclosure_n639_arg\ := \$13925_offsetclosure_n639_arg%now\;
      \$14898_v\ := \$14898_v%now\;
      \$14693_modulo6685896_result\ := \$14693_modulo6685896_result%now\;
      \$15497_r\ := \$15497_r%now\;
      \$13105_copy_root_in_ram6635884_id\ := \$13105_copy_root_in_ram6635884_id%now\;
      \$17434\ := \$17434%now\;
      \$16515\ := \$16515%now\;
      \$14512_v\ := \$14512_v%now\;
      \$14300_v\ := \$14300_v%now\;
      \$18261\ := \$18261%now\;
      \$17207_arg\ := \$17207_arg%now\;
      \$13315\ := \$13315%now\;
      \$18992\ := \$18992%now\;
      \$18344\ := \$18344%now\;
      \$17183\ := \$17183%now\;
      \$v7032\ := \$v7032%now\;
      result6112 := \result6112%now\;
      \$v5960\ := \$v5960%now\;
      \$v7084\ := \$v7084%now\;
      \$v6639\ := \$v6639%now\;
      \$v7060\ := \$v7060%now\;
      \$18030_w\ := \$18030_w%now\;
      \$18190\ := \$18190%now\;
      \$16380_v\ := \$16380_v%now\;
      \$v6295\ := \$v6295%now\;
      \$18924\ := \$18924%now\;
      \$12659\ := \$12659%now\;
      \$v6111\ := \$v6111%now\;
      \$v6011\ := \$v6011%now\;
      \$12891_copy_root_in_ram6635884_result\ := \$12891_copy_root_in_ram6635884_result%now\;
      \$18621\ := \$18621%now\;
      \$14185_next_env\ := \$14185_next_env%now\;
      \$17166\ := \$17166%now\;
      \$v6059\ := \$v6059%now\;
      \$12703\ := \$12703%now\;
      \$v6358\ := \$v6358%now\;
      \$12832\ := \$12832%now\;
      \$15684_compare6445897_result\ := \$15684_compare6445897_result%now\;
      \$v7111\ := \$v7111%now\;
      \$17895\ := \$17895%now\;
      \$13812\ := \$13812%now\;
      \$18632_loop666_id\ := \$18632_loop666_id%now\;
      \$17952_w\ := \$17952_w%now\;
      \$13820\ := \$13820%now\;
      \$13533\ := \$13533%now\;
      \$15805_binop_compare6455921_result\ := \$15805_binop_compare6455921_result%now\;
      \$15413_modulo6685896_id\ := \$15413_modulo6685896_id%now\;
      \$13977_v\ := \$13977_v%now\;
      \$v6294\ := \$v6294%now\;
      \$12857_forever6705883_id\ := \$12857_forever6705883_id%now\;
      \$v7438\ := \$v7438%now\;
      \$v7082\ := \$v7082%now\;
      \$v6415\ := \$v6415%now\;
      \$v5982\ := \$v5982%now\;
      \$19265\ := \$19265%now\;
      \$17011\ := \$17011%now\;
      \$v7012\ := \$v7012%now\;
      \$17505_forever6705894_id\ := \$17505_forever6705894_id%now\;
      \$v7282\ := \$v7282%now\;
      \$12813\ := \$12813%now\;
      \$17499\ := \$17499%now\;
      \$v6457\ := \$v6457%now\;
      \$13150\ := \$13150%now\;
      \$17808\ := \$17808%now\;
      \$v6820\ := \$v6820%now\;
      \$17970\ := \$17970%now\;
      \$12803_loop666_result\ := \$12803_loop666_result%now\;
      \$v7276\ := \$v7276%now\;
      \$14964_binop_int6435905_result\ := \$14964_binop_int6435905_result%now\;
      \$v7134\ := \$v7134%now\;
      \$17809\ := \$17809%now\;
      \$16404\ := \$16404%now\;
      \$v7157\ := \$v7157%now\;
      \$17969\ := \$17969%now\;
      \$v6280\ := \$v6280%now\;
      \$12845\ := \$12845%now\;
      \$v6361\ := \$v6361%now\;
      \$12561\ := \$12561%now\;
      \$17545\ := \$17545%now\;
      \$18634_aux664_id\ := \$18634_aux664_id%now\;
      \$15410_r\ := \$15410_r%now\;
      \$v6582\ := \$v6582%now\;
      \$v6600\ := \$v6600%now\;
      \$15062_res\ := \$15062_res%now\;
      \$v6264\ := \$v6264%now\;
      \$14342\ := \$14342%now\;
      \$v6691\ := \$v6691%now\;
      \$12562\ := \$12562%now\;
      result5939 := \result5939%now\;
      \$12657\ := \$12657%now\;
      \$v7130\ := \$v7130%now\;
      \$16193\ := \$16193%now\;
      \$16916_compare6445898_result\ := \$16916_compare6445898_result%now\;
      \$18839\ := \$18839%now\;
      \$13787\ := \$13787%now\;
      \$v7303\ := \$v7303%now\;
      \$19146\ := \$19146%now\;
      \$15684_compare6445897_arg\ := \$15684_compare6445897_arg%now\;
      \$15142_res\ := \$15142_res%now\;
      \$12905\ := \$12905%now\;
      \$v6267\ := \$v6267%now\;
      \$18658\ := \$18658%now\;
      \$13386\ := \$13386%now\;
      \$17465\ := \$17465%now\;
      \$v6477\ := \$v6477%now\;
      \$13025\ := \$13025%now\;
      \$18678\ := \$18678%now\;
      \$16461\ := \$16461%now\;
      \$v6774\ := \$v6774%now\;
      \$18180_hd\ := \$18180_hd%now\;
      \$v6811\ := \$v6811%now\;
      \$13791\ := \$13791%now\;
      \$14464_v\ := \$14464_v%now\;
      \$15851_argument1\ := \$15851_argument1%now\;
      \$13022\ := \$13022%now\;
      \$15101_modulo6685888_arg\ := \$15101_modulo6685888_arg%now\;
      \$13124\ := \$13124%now\;
      \$v6762\ := \$v6762%now\;
      \$v6720\ := \$v6720%now\;
      \$v6528\ := \$v6528%now\;
      \$v6083\ := \$v6083%now\;
      \$16724\ := \$16724%now\;
      \$v6524\ := \$v6524%now\;
      \$v6448\ := \$v6448%now\;
      \$17184\ := \$17184%now\;
      \$13228\ := \$13228%now\;
      \$19139\ := \$19139%now\;
      \$v7036\ := \$v7036%now\;
      \$v6755\ := \$v6755%now\;
      \$17533\ := \$17533%now\;
      result5974 := \result5974%now\;
      \$v7037\ := \$v7037%now\;
      \$18589\ := \$18589%now\;
      \$14669_modulo6685895_result\ := \$14669_modulo6685895_result%now\;
      \$13813\ := \$13813%now\;
      \$17105_w06555936_result\ := \$17105_w06555936_result%now\;
      \$13921_loop665_arg\ := \$13921_loop665_arg%now\;
      \$17599\ := \$17599%now\;
      \$13921_loop665_result\ := \$13921_loop665_result%now\;
      \$v7401\ := \$v7401%now\;
      \$v6980\ := \$v6980%now\;
      \$16337\ := \$16337%now\;
      \$17534\ := \$17534%now\;
      \$12558\ := \$12558%now\;
      \$v6926\ := \$v6926%now\;
      \$16811_compare6445898_id\ := \$16811_compare6445898_id%now\;
      \$v5989\ := \$v5989%now\;
      \$14103\ := \$14103%now\;
      \$15556_modulo6685895_arg\ := \$15556_modulo6685895_arg%now\;
      \$19147\ := \$19147%now\;
      \$16383\ := \$16383%now\;
      \$v7149\ := \$v7149%now\;
      \$13314\ := \$13314%now\;
      \$15639_v\ := \$15639_v%now\;
      \$16624_argument2\ := \$16624_argument2%now\;
      \$15069_modulo6685895_result\ := \$15069_modulo6685895_result%now\;
      \$16662_fill6535928_id\ := \$16662_fill6535928_id%now\;
      rdy6113 := \rdy6113%now\;
      \$17542\ := \$17542%now\;
      \$v6345\ := \$v6345%now\;
      \$v6194\ := \$v6194%now\;
      \$v6571\ := \$v6571%now\;
      \$15531_binop_int6435913_result\ := \$15531_binop_int6435913_result%now\;
      \$v6439\ := \$v6439%now\;
      \$v6079\ := \$v6079%now\;
      \$15621_forever6705915_arg\ := \$15621_forever6705915_arg%now\;
      \$17884\ := \$17884%now\;
      \$v7097\ := \$v7097%now\;
      \$13927_branch_if648_id\ := \$13927_branch_if648_id%now\;
      \$14982_res\ := \$14982_res%now\;
      \$18353\ := \$18353%now\;
      \$v7347\ := \$v7347%now\;
      \$16846_compare6445898_arg\ := \$16846_compare6445898_arg%now\;
      \$v6895\ := \$v6895%now\;
      \$16195_forever6705924_arg\ := \$16195_forever6705924_arg%now\;
      \$17589\ := \$17589%now\;
      \$13017\ := \$13017%now\;
      \$15747_v\ := \$15747_v%now\;
      \$16662_fill6535928_result\ := \$16662_fill6535928_result%now\;
      \$18345\ := \$18345%now\;
      \$v7122\ := \$v7122%now\;
      \$17048_w16565937_id\ := \$17048_w16565937_id%now\;
      \$18686_copy_root_in_ram6635880_result\ := \$18686_copy_root_in_ram6635880_result%now\;
      \$15093_modulo6685896_id\ := \$15093_modulo6685896_id%now\;
      \$18736\ := \$18736%now\;
      \$18671\ := \$18671%now\;
      \$15500_modulo6685896_id\ := \$15500_modulo6685896_id%now\;
      \$v7226\ := \$v7226%now\;
      \$17459_loop665_id\ := \$17459_loop665_id%now\;
      \$15333_modulo6685896_arg\ := \$15333_modulo6685896_arg%now\;
      \$17807\ := \$17807%now\;
      \$v6220\ := \$v6220%now\;
      \$13821\ := \$13821%now\;
      \$18035_hd\ := \$18035_hd%now\;
      \$v6290\ := \$v6290%now\;
      \$17172\ := \$17172%now\;
      \$13394\ := \$13394%now\;
      \$19338\ := \$19338%now\;
      \$17368_v\ := \$17368_v%now\;
      \$v5871\ := \$v5871%now\;
      \$13958\ := \$13958%now\;
      \$12824\ := \$12824%now\;
      \$17562\ := \$17562%now\;
      \$16322\ := \$16322%now\;
      \$v7105\ := \$v7105%now\;
      \$13698\ := \$13698%now\;
      \$17520_copy_root_in_ram6635893_arg\ := \$17520_copy_root_in_ram6635893_arg%now\;
      \$15556_modulo6685895_id\ := \$15556_modulo6685895_id%now\;
      \$13105_copy_root_in_ram6635884_result\ := \$13105_copy_root_in_ram6635884_result%now\;
      \$12891_copy_root_in_ram6635884_id\ := \$12891_copy_root_in_ram6635884_id%now\;
      \$12806_loop666_arg\ := \$12806_loop666_arg%now\;
      \$v6566\ := \$v6566%now\;
      \$15181_modulo6685888_id\ := \$15181_modulo6685888_id%now\;
      \$v7080\ := \$v7080%now\;
      \$v6675\ := \$v6675%now\;
      \$v6576\ := \$v6576%now\;
      \$16998_argument3\ := \$16998_argument3%now\;
      \$v7423\ := \$v7423%now\;
      \$18728\ := \$18728%now\;
      \$16157\ := \$16157%now\;
      \$13684_hd\ := \$13684_hd%now\;
      \$19111\ := \$19111%now\;
      \$v6647\ := \$v6647%now\;
      \$13091\ := \$13091%now\;
      \$13143_hd\ := \$13143_hd%now\;
      \$18793_copy_root_in_ram6635879_result\ := \$18793_copy_root_in_ram6635879_result%now\;
      \$15769_binop_compare6455920_result\ := \$15769_binop_compare6455920_result%now\;
      \$16462\ := \$16462%now\;
      \$14265\ := \$14265%now\;
      \$12916\ := \$12916%now\;
      \$v6244\ := \$v6244%now\;
      \$12742\ := \$12742%now\;
      \$13119\ := \$13119%now\;
      \$13972_v\ := \$13972_v%now\;
      \$14884_binop_int6435904_result\ := \$14884_binop_int6435904_result%now\;
      \$13951\ := \$13951%now\;
      \$v7024\ := \$v7024%now\;
      \$13923_make_block579_arg\ := \$13923_make_block579_arg%now\;
      \$15648_compare6445897_result\ := \$15648_compare6445897_result%now\;
      \$17330_sp\ := \$17330_sp%now\;
      \$v6620\ := \$v6620%now\;
      \$17353\ := \$17353%now\;
      \$v6983\ := \$v6983%now\;
      \$v7257\ := \$v7257%now\;
      \$v6663\ := \$v6663%now\;
      \$13118\ := \$13118%now\;
      \$v6032\ := \$v6032%now\;
      \$18672\ := \$18672%now\;
      \$19074\ := \$19074%now\;
      \$15309_modulo6685895_id\ := \$15309_modulo6685895_id%now\;
      \$v6260\ := \$v6260%now\;
      \$19076\ := \$19076%now\;
      rdy5975 := \rdy5975%now\;
      \$15124_binop_int6435907_result\ := \$15124_binop_int6435907_result%now\;
      \$16334_v\ := \$16334_v%now\;
      \$v7270\ := \$v7270%now\;
      \$18042\ := \$18042%now\;
      \$18611\ := \$18611%now\;
      \$14377_v\ := \$14377_v%now\;
      \$16381_v\ := \$16381_v%now\;
      \$v6076\ := \$v6076%now\;
      \$15908\ := \$15908%now\;
      \$12563\ := \$12563%now\;
      \$v7026\ := \$v7026%now\;
      \$v6698\ := \$v6698%now\;
      \$15013_modulo6685896_result\ := \$15013_modulo6685896_result%now\;
      \$12805_aux664_arg\ := \$12805_aux664_arg%now\;
      \$v7075\ := \$v7075%now\;
      \$13024\ := \$13024%now\;
      \$13965\ := \$13965%now\;
      \$18573\ := \$18573%now\;
      \$v6124\ := \$v6124%now\;
      \$17481\ := \$17481%now\;
      \$v6215\ := \$v6215%now\;
      \$15720_compare6445897_result\ := \$15720_compare6445897_result%now\;
      \$v7160\ := \$v7160%now\;
      \$v6497\ := \$v6497%now\;
      \$15044_binop_int6435906_arg\ := \$15044_binop_int6435906_arg%now\;
      \$13097\ := \$13097%now\;
      \$17456_loop665_arg\ := \$17456_loop665_arg%now\;
      \$13952\ := \$13952%now\;
      \$15093_modulo6685896_result\ := \$15093_modulo6685896_result%now\;
      \$13924_apply638_id\ := \$13924_apply638_id%now\;
      \$v6556\ := \$v6556%now\;
      \$14701_modulo6685888_id\ := \$14701_modulo6685888_id%now\;
      \$12687\ := \$12687%now\;
      \$15473_r\ := \$15473_r%now\;
      \$17061\ := \$17061%now\;
      \$16725\ := \$16725%now\;
      \$v6412\ := \$v6412%now\;
      \$v7407\ := \$v7407%now\;
      \$v6747\ := \$v6747%now\;
      \$12831\ := \$12831%now\;
      \$16651\ := \$16651%now\;
      \$14781_modulo6685888_id\ := \$14781_modulo6685888_id%now\;
      \$16658\ := \$16658%now\;
      \$v7136\ := \$v7136%now\;
      \$14589_modulo6685895_id\ := \$14589_modulo6685895_id%now\;
      \$v5968\ := \$v5968%now\;
      \$v6339\ := \$v6339%now\;
      \$16788_compbranch6505930_id\ := \$16788_compbranch6505930_id%now\;
      \$17486\ := \$17486%now\;
      \$v6331\ := \$v6331%now\;
      \$18553\ := \$18553%now\;
      \$14034_v\ := \$14034_v%now\;
      \$v7410\ := \$v7410%now\;
      \$v7131\ := \$v7131%now\;
      \$18284\ := \$18284%now\;
      \$v7390\ := \$v7390%now\;
      \$13306\ := \$13306%now\;
      \$v6539\ := \$v6539%now\;
      \$v7341\ := \$v7341%now\;
      \$15090_r\ := \$15090_r%now\;
      \$14906_r\ := \$14906_r%now\;
      \$13462\ := \$13462%now\;
      \$19270\ := \$19270%now\;
      \$v6850\ := \$v6850%now\;
      \$v7430\ := \$v7430%now\;
      \$v6671\ := \$v6671%now\;
      \$15149_modulo6685895_result\ := \$15149_modulo6685895_result%now\;
      \$15756_compare6445897_id\ := \$15756_compare6445897_id%now\;
      \$v6418\ := \$v6418%now\;
      \$v6250\ := \$v6250%now\;
      \$v6051\ := \$v6051%now\;
      \$15621_forever6705915_id\ := \$15621_forever6705915_id%now\;
      \$v6886\ := \$v6886%now\;
      \$16858_compbranch6505932_result\ := \$16858_compbranch6505932_result%now\;
      \$15222_res\ := \$15222_res%now\;
      \$v6770\ := \$v6770%now\;
      \$v7040\ := \$v7040%now\;
      \$16301\ := \$16301%now\;
      \$13911\ := \$13911%now\;
      \$17680\ := \$17680%now\;
      \$v6191\ := \$v6191%now\;
      \$15138_v\ := \$15138_v%now\;
      \$v6486\ := \$v6486%now\;
      \$13152\ := \$13152%now\;
      \$16155\ := \$16155%now\;
      \$14933_modulo6685896_arg\ := \$14933_modulo6685896_arg%now\;
      \$12693\ := \$12693%now\;
      \$v7106\ := \$v7106%now\;
      \$v7067\ := \$v7067%now\;
      \$13920_loop666_result\ := \$13920_loop666_result%now\;
      \$16293\ := \$16293%now\;
      \$13159\ := \$13159%now\;
      \$13953\ := \$13953%now\;
      \$15625_binop_compare6455916_arg\ := \$15625_binop_compare6455916_arg%now\;
      \$13015\ := \$13015%now\;
      \$17799_hd\ := \$17799_hd%now\;
      \$v6039\ := \$v6039%now\;
      \$15611\ := \$15611%now\;
      \$v6808\ := \$v6808%now\;
      \$17444\ := \$17444%now\;
      \$14853_modulo6685896_id\ := \$14853_modulo6685896_id%now\;
      \$18665\ := \$18665%now\;
      \$19132_hd\ := \$19132_hd%now\;
      \$16313_v\ := \$16313_v%now\;
      \$14757_modulo6685888_arg\ := \$14757_modulo6685888_arg%now\;
      \$18710\ := \$18710%now\;
      \$v5979\ := \$v5979%now\;
      \$v6006\ := \$v6006%now\;
      \$14621_modulo6685888_id\ := \$14621_modulo6685888_id%now\;
      \$14941_modulo6685888_id\ := \$14941_modulo6685888_id%now\;
      \$19073\ := \$19073%now\;
      \$15733_binop_compare6455919_id\ := \$15733_binop_compare6455919_id%now\;
      \$15620\ := \$15620%now\;
      \$17596\ := \$17596%now\;
      \$16413\ := \$16413%now\;
      \$19141\ := \$19141%now\;
      \$17753\ := \$17753%now\;
      \$16706\ := \$16706%now\;
      \$16296\ := \$16296%now\;
      \$v7001\ := \$v7001%now\;
      \$18468\ := \$18468%now\;
      \$19000\ := \$19000%now\;
      \$v5877\ := \$v5877%now\;
      \$16951_compare6445898_id\ := \$16951_compare6445898_id%now\;
      \$13231\ := \$13231%now\;
      \$v6024\ := \$v6024%now\;
      \$13130\ := \$13130%now\;
      \$15469_res\ := \$15469_res%now\;
      \$18471\ := \$18471%now\;
      \$v6793\ := \$v6793%now\;
      \$v7266\ := \$v7266%now\;
      \$18350\ := \$18350%now\;
      \$16357\ := \$16357%now\;
      \$15149_modulo6685895_arg\ := \$15149_modulo6685895_arg%now\;
      \$13987_v\ := \$13987_v%now\;
      \$v7055\ := \$v7055%now\;
      \$17483\ := \$17483%now\;
      \$14260\ := \$14260%now\;
      \$15588_modulo6685888_id\ := \$15588_modulo6685888_id%now\;
      \$v7309\ := \$v7309%now\;
      \$15643_res\ := \$15643_res%now\;
      \$13078_copy_root_in_ram6635885_arg\ := \$13078_copy_root_in_ram6635885_arg%now\;
      \$18914\ := \$18914%now\;
      \$17660_w\ := \$17660_w%now\;
      \$16846_compare6445898_result\ := \$16846_compare6445898_result%now\;
      \$18817\ := \$18817%now\;
      \$v6871\ := \$v6871%now\;
      \$17672\ := \$17672%now\;
      \$19148\ := \$19148%now\;
      \$v7329\ := \$v7329%now\;
      \$19072\ := \$19072%now\;
      \$15733_binop_compare6455919_result\ := \$15733_binop_compare6455919_result%now\;
      \$14081\ := \$14081%now\;
      \$18545\ := \$18545%now\;
      \$13889\ := \$13889%now\;
      \$14015\ := \$14015%now\;
      \$12840_next\ := \$12840_next%now\;
      \$18686_copy_root_in_ram6635880_arg\ := \$18686_copy_root_in_ram6635880_arg%now\;
      \$14742_res\ := \$14742_res%now\;
      \$14586_r\ := \$14586_r%now\;
      \$18195\ := \$18195%now\;
      \$v6540\ := \$v6540%now\;
      \$18793_copy_root_in_ram6635879_arg\ := \$18793_copy_root_in_ram6635879_arg%now\;
      \$15317_modulo6685888_id\ := \$15317_modulo6685888_id%now\;
      \$16551_compbranch6505926_result\ := \$16551_compbranch6505926_result%now\;
      \$17811\ := \$17811%now\;
      \$16980_b\ := \$16980_b%now\;
      \$18349\ := \$18349%now\;
      \$15451_binop_int6435912_id\ := \$15451_binop_int6435912_id%now\;
      \$14002_v\ := \$14002_v%now\;
      \$14997_modulo6685888_arg\ := \$14997_modulo6685888_arg%now\;
      \$16335_v\ := \$16335_v%now\;
      \$13014\ := \$13014%now\;
      \$v6977\ := \$v6977%now\;
      \$18039\ := \$18039%now\;
      \$13448\ := \$13448%now\;
      \$17571\ := \$17571%now\;
      \$17757\ := \$17757%now\;
      \$v6018\ := \$v6018%now\;
      \$16358\ := \$16358%now\;
      \$v7052\ := \$v7052%now\;
      \$17352\ := \$17352%now\;
      \$17756\ := \$17756%now\;
      \$v6141\ := \$v6141%now\;
      \$13391\ := \$13391%now\;
      \$v6086\ := \$v6086%now\;
      \$v6145\ := \$v6145%now\;
      \$15066_r\ := \$15066_r%now\;
      result6147 := \result6147%now\;
      \$15446\ := \$15446%now\;
      \$v6877\ := \$v6877%now\;
      \$16041_v\ := \$16041_v%now\;
      \$16063_w6515922_arg\ := \$16063_w6515922_arg%now\;
      \$12700\ := \$12700%now\;
      \$16951_compare6445898_result\ := \$16951_compare6445898_result%now\;
      \$v6210\ := \$v6210%now\;
      \$15564_modulo6685888_id\ := \$15564_modulo6685888_id%now\;
      \$12721\ := \$12721%now\;
      \$18920\ := \$18920%now\;
      \$14393_hd\ := \$14393_hd%now\;
      \$18282\ := \$18282%now\;
      \$v7141\ := \$v7141%now\;
      \$15157_modulo6685888_result\ := \$15157_modulo6685888_result%now\;
      \$14850_r\ := \$14850_r%now\;
      \$17601\ := \$17601%now\;
      \$v6310\ := \$v6310%now\;
      \$14493_v\ := \$14493_v%now\;
      \$12711\ := \$12711%now\;
      \$v5864\ := \$v5864%now\;
      \$v6483\ := \$v6483%now\;
      \$13819\ := \$13819%now\;
      \$v7325\ := \$v7325%now\;
      \$13120\ := \$13120%now\;
      \$v7087\ := \$v7087%now\;
      \$v6615\ := \$v6615%now\;
      \$15146_r\ := \$15146_r%now\;
      \$v7394\ := \$v7394%now\;
      \$18347\ := \$18347%now\;
      \$18700\ := \$18700%now\;
      \$v6777\ := \$v6777%now\;
      \$12940\ := \$12940%now\;
      \$v7173\ := \$v7173%now\;
      \$17062\ := \$17062%now\;
      \$v7073\ := \$v7073%now\;
      \$14025_v\ := \$14025_v%now\;
      \$14561\ := \$14561%now\;
      \$16437_v\ := \$16437_v%now\;
      \$15549_res\ := \$15549_res%now\;
      \$15253_modulo6685896_arg\ := \$15253_modulo6685896_arg%now\;
      \$15013_modulo6685896_arg\ := \$15013_modulo6685896_arg%now\;
      \$14822_res\ := \$14822_res%now\;
      \$18847\ := \$18847%now\;
      \$18840\ := \$18840%now\;
      \$18340_hd\ := \$18340_hd%now\;
      \$v7148\ := \$v7148%now\;
      \$14884_binop_int6435904_id\ := \$14884_binop_int6435904_id%now\;
      \$18632_loop666_result\ := \$18632_loop666_result%now\;
      \$15226_r\ := \$15226_r%now\;
      \$18422\ := \$18422%now\;
      \$15444\ := \$15444%now\;
      \$19137\ := \$19137%now\;
      \$18923\ := \$18923%now\;
      \$17161\ := \$17161%now\;
      \$12662\ := \$12662%now\;
      \$v7065\ := \$v7065%now\;
      \$14662_res\ := \$14662_res%now\;
      \$v6226\ := \$v6226%now\;
      \$v7319\ := \$v7319%now\;
      \$17396\ := \$17396%now\;
      \$17806\ := \$17806%now\;
      \$v6612\ := \$v6612%now\;
      \$15805_binop_compare6455921_id\ := \$15805_binop_compare6455921_id%now\;
      \$13305\ := \$13305%now\;
      \$13230\ := \$13230%now\;
      \$19056\ := \$19056%now\;
      \$18469\ := \$18469%now\;
      \$v7286\ := \$v7286%now\;
      \$13534\ := \$13534%now\;
      \$v7152\ := \$v7152%now\;
      \$v6929\ := \$v6929%now\;
      \$16910_b\ := \$16910_b%now\;
      \$v7043\ := \$v7043%now\;
      \$12850\ := \$12850%now\;
      \$17456_loop665_id\ := \$17456_loop665_id%now\;
      \$18477\ := \$18477%now\;
      \$v7225\ := \$v7225%now\;
      \$v6923\ := \$v6923%now\;
      \$v6674\ := \$v6674%now\;
      \$13699\ := \$13699%now\;
      \$v6944\ := \$v6944%now\;
      \$13923_make_block579_id\ := \$13923_make_block579_id%now\;
      \$14207_loop_push6495899_id\ := \$14207_loop_push6495899_id%now\;
      \$15648_compare6445897_arg\ := \$15648_compare6445897_arg%now\;
      \$13803_w\ := \$13803_w%now\;
      \$17780\ := \$17780%now\;
      \$12876\ := \$12876%now\;
      \$18656\ := \$18656%now\;
      \$v6687\ := \$v6687%now\;
      \$v6107\ := \$v6107%now\;
      \$12661\ := \$12661%now\;
      \$v6630\ := \$v6630%now\;
      \$15697_binop_compare6455918_id\ := \$15697_binop_compare6455918_id%now\;
      \$v7124\ := \$v7124%now\;
      \$v7384\ := \$v7384%now\;
      \$v7063\ := \$v7063%now\;
      \$13928_w652_arg\ := \$13928_w652_arg%now\;
      \$15465_v\ := \$15465_v%now\;
      \$13622\ := \$13622%now\;
      \$14355\ := \$14355%now\;
      \$v7312\ := \$v7312%now\;
      \$v6636\ := \$v6636%now\;
      \$14770_r\ := \$14770_r%now\;
      \$v6063\ := \$v6063%now\;
      \$15013_modulo6685896_id\ := \$15013_modulo6685896_id%now\;
      \$14690_r\ := \$14690_r%now\;
      \$12807_loop665_arg\ := \$12807_loop665_arg%now\;
      \$v6120\ := \$v6120%now\;
      \$17810\ := \$17810%now\;
      \$v6168\ := \$v6168%now\;
      \$v7053\ := \$v7053%now\;
      \$v7239\ := \$v7239%now\;
      \$17236\ := \$17236%now\;
      \$v7209\ := \$v7209%now\;
      \$13128\ := \$13128%now\;
      \$15229_modulo6685895_id\ := \$15229_modulo6685895_id%now\;
      \$v7316\ := \$v7316%now\;
      \$12690\ := \$12690%now\;
      \$13925_offsetclosure_n639_id\ := \$13925_offsetclosure_n639_id%now\;
      \$13020\ := \$13020%now\;
      \$v6932\ := \$v6932%now\;
      \$12539\ := \$12539%now\;
      \$v6592\ := \$v6592%now\;
      \$v6010\ := \$v6010%now\;
      \$13093\ := \$13093%now\;
      \$18323\ := \$18323%now\;
      \$17965\ := \$17965%now\;
      \$v5971\ := \$v5971%now\;
      \$16659_sp\ := \$16659_sp%now\;
      \$17547_copy_root_in_ram6635891_result\ := \$17547_copy_root_in_ram6635891_result%now\;
      \$13690\ := \$13690%now\;
      \$13628\ := \$13628%now\;
      \$v6349\ := \$v6349%now\;
      \$13465\ := \$13465%now\;
      \$12812\ := \$12812%now\;
      \$v6028\ := \$v6028%now\;
      \$13374_w\ := \$13374_w%now\;
      \$14368\ := \$14368%now\;
      \$12718\ := \$12718%now\;
      \$17784\ := \$17784%now\;
      \$15508_modulo6685888_id\ := \$15508_modulo6685888_id%now\;
      \$15364_binop_int6435910_result\ := \$15364_binop_int6435910_result%now\;
      \$14613_modulo6685896_arg\ := \$14613_modulo6685896_arg%now\;
      \$15751_res\ := \$15751_res%now\;
      \$13537\ := \$13537%now\;
      \$12654\ := \$12654%now\;
      \$v7071\ := \$v7071%now\;
      \$v6311\ := \$v6311%now\;
      \$ram_lock\ := \$ram_lock%now\;
      \$global_end_lock\ := \$global_end_lock%now\;
      \$code_lock\ := \$code_lock%now\;
      state := \state%now\;
      state_var7464 := \state_var7464%now\;
      state_var7463 := \state_var7463%now\;
      state_var7462 := \state_var7462%now\;
      state_var7461 := \state_var7461%now\;
      state_var7460 := \state_var7460%now\;
      case state is
      when \$12520_LOOP666\ =>
        \$v5948\ := work.Int.ge(\$12520_loop666_arg\(0 to 15), work.Int.add(
                                                               \$12520_loop666_arg\(48 to 63), X"000" & X"1"));
        if \$v5948\(0) = '1' then
          \$12520_loop666_result\ := eclat_unit;
          \$19270\ := \$12520_loop666_result\;
          \$v5957\ := \$ram_lock\;
          if \$v5957\(0) = '1' then
            state := Q_WAIT5956;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$19235\(0 to 30),16)));
            \$ram_write\ <= eclat_resize(\$12521_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
            state := PAUSE_SET5955;
          end if;
        else
          \$v5947\ := \$ram_lock\;
          if \$v5947\(0) = '1' then
            state := Q_WAIT5946;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$12520_loop666_arg\(32 to 47), \$12520_loop666_arg\(0 to 15))));
            state := PAUSE_GET5945;
          end if;
        end if;
      when \$12521_LOOP665\ =>
        \$v5972\ := work.Int.ge(\$12521_loop665_arg\(0 to 15), work.Int.add(
                                                               \$12521_loop665_arg\(80 to 95), X"000" & X"1"));
        if \$v5972\(0) = '1' then
          \$12521_loop665_result\ := \$12521_loop665_arg\(16 to 31);
          state := \$12521_LOOP665\;
        else
          \$v5971\ := \$ram_lock\;
          if \$v5971\(0) = '1' then
            state := Q_WAIT5970;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$12521_loop665_arg\(64 to 79), \$12521_loop665_arg\(0 to 15))));
            state := PAUSE_GET5969;
          end if;
        end if;
      when \$12522_WAIT662\ =>
        if \$v5864\(0) = '1' then
          
        else
          \$v5864\ := eclat_true;
          \$18621\ := \$12522_wait662_arg\(1 to 32) & \$12522_wait662_arg\(33 to 64) & X"0" & X"fa0" & X"0" & X"fa0" & X"0" & X"fa0" & 
          work.Int.add(X"0" & X"fa0", X"1770") & eclat_false;
        end if;
        case state_var7464 is
        when \$18632_LOOP666\ =>
          \$v5983\ := work.Int.ge(\$18632_loop666_arg\(0 to 15), work.Int.add(
                                                                 \$18632_loop666_arg\(48 to 63), X"000" & X"1"));
          if \$v5983\(0) = '1' then
            \$18632_loop666_result\ := eclat_unit;
            case \$18632_loop666_id\ is
            when "000000000010" =>
              \$19146\ := \$18632_loop666_result\;
              \$v5992\ := \$ram_lock\;
              if \$v5992\(0) = '1' then
                state_var7464 := Q_WAIT5991;
              else
                acquire(\$ram_lock\);
                \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$19111\(0 to 30),16)));
                \$ram_write\ <= eclat_resize(\$18633_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                state_var7464 := PAUSE_SET5990;
              end if;
            when "000000000110" =>
              \$18738\ := \$18632_loop666_result\;
              \$v6021\ := \$ram_lock\;
              if \$v6021\(0) = '1' then
                state_var7464 := Q_WAIT6020;
              else
                acquire(\$ram_lock\);
                \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18701\(0 to 30),16)));
                \$ram_write\ <= eclat_resize(\$18686_copy_root_in_ram6635880_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                state_var7464 := PAUSE_SET6019;
              end if;
            when "000000001000" =>
              \$18845\ := \$18632_loop666_result\;
              \$v6048\ := \$ram_lock\;
              if \$v6048\(0) = '1' then
                state_var7464 := Q_WAIT6047;
              else
                acquire(\$ram_lock\);
                \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18808\(0 to 30),16)));
                \$ram_write\ <= eclat_resize(\$18793_copy_root_in_ram6635879_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                state_var7464 := PAUSE_SET6046;
              end if;
            when "000000001010" =>
              \$18923\ := \$18632_loop666_result\;
              \$v6069\ := \$ram_lock\;
              if \$v6069\(0) = '1' then
                state_var7464 := Q_WAIT6068;
              else
                acquire(\$ram_lock\);
                \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$12522_wait662_arg\(33 to 63),16)));
                \$ram_write\ <= eclat_resize(\$18644\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                state_var7464 := PAUSE_SET6067;
              end if;
            when "000000001011" =>
              \$19001\ := \$18632_loop666_result\;
              \$v6086\ := \$ram_lock\;
              if \$v6086\(0) = '1' then
                state_var7464 := Q_WAIT6085;
              else
                acquire(\$ram_lock\);
                \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$12522_wait662_arg\(1 to 31),16)));
                \$ram_write\ <= eclat_resize(\$18621\(112 to 127),31) & eclat_false; \$ram_write_request\ <= '1';
                state_var7464 := PAUSE_SET6084;
              end if;
            when others =>
              
            end case;
          else
            \$v5982\ := \$ram_lock\;
            if \$v5982\(0) = '1' then
              state_var7464 := Q_WAIT5981;
            else
              acquire(\$ram_lock\);
              \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$18632_loop666_arg\(32 to 47), \$18632_loop666_arg\(0 to 15))));
              state_var7464 := PAUSE_GET5980;
            end if;
          end if;
        when \$18633_LOOP665\ =>
          \$v6007\ := work.Int.ge(\$18633_loop665_arg\(0 to 15), work.Int.add(
                                                                 \$18633_loop665_arg\(80 to 95), X"000" & X"1"));
          if \$v6007\(0) = '1' then
            \$18633_loop665_result\ := \$18633_loop665_arg\(16 to 31);
            \$19080_next\ := \$18633_loop665_result\;
            \$18634_aux664_arg\ := work.Int.add(\$18634_aux664_arg\(0 to 15), 
                                                work.Int.add(eclat_resize(
                                                             work.Int.lsr(
                                                             eclat_resize(eclat_resize(\$19076\(0 to 30),16),31), X"0000000" & X"2"),16), X"000" & X"1")) & \$19080_next\ & \$18634_aux664_arg\(32 to 47) & \$18634_aux664_arg\(48 to 63);
            state_var7464 := \$18634_AUX664\;
          else
            \$v6006\ := \$ram_lock\;
            if \$v6006\(0) = '1' then
              state_var7464 := Q_WAIT6005;
            else
              acquire(\$ram_lock\);
              \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$18633_loop665_arg\(64 to 79), \$18633_loop665_arg\(0 to 15))));
              state_var7464 := PAUSE_GET6004;
            end if;
          end if;
        when \$18634_AUX664\ =>
          \$19070\ := work.Print.print_string(clk,of_string("     scan="));
          \$19071\ := work.Int.print(clk,\$18634_aux664_arg\(0 to 15));
          \$19072\ := work.Print.print_string(clk,of_string(" | next="));
          \$19073\ := work.Int.print(clk,\$18634_aux664_arg\(16 to 31));
          \$19074\ := work.Print.print_newline(clk,eclat_unit);
          \$v6011\ := work.Int.ge(\$18634_aux664_arg\(0 to 15), \$18634_aux664_arg\(16 to 31));
          if \$v6011\(0) = '1' then
            \$18634_aux664_result\ := \$18634_aux664_arg\(16 to 31);
            \$18670_next\ := \$18634_aux664_result\;
            \$18671\ := work.Print.print_string(clk,of_string("memory copied in to_space : "));
            \$18672\ := work.Int.print(clk,work.Int.sub(\$18670_next\, \$18621\(112 to 127)));
            \$18673\ := work.Print.print_string(clk,of_string(" words"));
            \$18674\ := work.Print.print_newline(clk,eclat_unit);
            \$v6012\ := work.Int.gt(work.Int.sub(\$18670_next\, \$18621\(112 to 127)), X"1770");
            if \$v6012\(0) = '1' then
              \$18676\ := work.Print.print_string(clk,of_string("fatal error: "));
              \$18677\ := work.Print.print_string(clk,of_string("Out of memory"));
              \$18678\ := work.Print.print_newline(clk,eclat_unit);
              \$18679_forever6705881_id\ := "000000000100";
              \$18679_forever6705881_arg\ := eclat_unit;
              state_var7464 := \$18679_FOREVER6705881\;
            else
              \$18650\ := \$18644\(0 to 31) & \$18661\(0 to 31) & \$18670_next\;
              \$18655\ := work.Print.print_newline(clk,eclat_unit);
              \$18656\ := work.Print.print_newline(clk,eclat_unit);
              \$18657\ := work.Print.print_string(clk,of_string("[================= GC END ======================]"));
              \$18660\ := work.Print.print_newline(clk,eclat_unit);
              \$18658\ := work.Print.print_newline(clk,eclat_unit);
              result5974 := \$18650\(0 to 31) & \$18650\(32 to 63) & \$18650\(64 to 79) & 
              work.Int.add(\$18650\(64 to 79), \$12522_wait662_arg\(81 to 96)) & \$18621\(112 to 127) & \$18621\(96 to 111);
              rdy5975 := eclat_true;
              state_var7464 := IDLE5976;
            end if;
          else
            \$v6010\ := \$ram_lock\;
            if \$v6010\(0) = '1' then
              state_var7464 := Q_WAIT6009;
            else
              acquire(\$ram_lock\);
              \$ram_ptr\ <= to_integer(unsigned(\$18634_aux664_arg\(0 to 15)));
              state_var7464 := PAUSE_GET6008;
            end if;
          end if;
        when \$18679_FOREVER6705881\ =>
          \$18679_forever6705881_arg\ := eclat_unit;
          state_var7464 := \$18679_FOREVER6705881\;
        when \$18686_COPY_ROOT_IN_RAM6635880\ =>
          \$v6036\ := work.Int.ge(\$18686_copy_root_in_ram6635880_arg\(0 to 15), \$18686_copy_root_in_ram6635880_arg\(16 to 31));
          if \$v6036\(0) = '1' then
            \$18686_copy_root_in_ram6635880_result\ := \$18686_copy_root_in_ram6635880_arg\(32 to 47);
            \$18666_next\ := \$18686_copy_root_in_ram6635880_result\;
            \$18668\ := work.Print.print_string(clk,of_string("======================================="));
            \$18669\ := work.Print.print_newline(clk,eclat_unit);
            \$18634_aux664_id\ := "000000000101";
            \$18634_aux664_arg\ := \$18621\(112 to 127) & \$18666_next\ & \$18621\(96 to 111) & \$18621\(112 to 127);
            state_var7464 := \$18634_AUX664\;
          else
            \$18698\ := work.Print.print_string(clk,of_string("racine:"));
            \$18699\ := work.Int.print(clk,\$18686_copy_root_in_ram6635880_arg\(0 to 15));
            \$18700\ := work.Print.print_newline(clk,eclat_unit);
            \$v6035\ := \$ram_lock\;
            if \$v6035\(0) = '1' then
              state_var7464 := Q_WAIT6034;
            else
              acquire(\$ram_lock\);
              \$ram_ptr\ <= to_integer(unsigned(\$18686_copy_root_in_ram6635880_arg\(0 to 15)));
              state_var7464 := PAUSE_GET6033;
            end if;
          end if;
        when \$18793_COPY_ROOT_IN_RAM6635879\ =>
          \$v6063\ := work.Int.ge(\$18793_copy_root_in_ram6635879_arg\(0 to 15), \$18793_copy_root_in_ram6635879_arg\(16 to 31));
          if \$v6063\(0) = '1' then
            \$18793_copy_root_in_ram6635879_result\ := \$18793_copy_root_in_ram6635879_arg\(32 to 47);
            \$18664_next\ := \$18793_copy_root_in_ram6635879_result\;
            \$v6039\ := \$global_end_lock\;
            if \$v6039\(0) = '1' then
              state_var7464 := Q_WAIT6038;
            else
              acquire(\$global_end_lock\);
              \$global_end_ptr\ <= 0;
              state_var7464 := PAUSE_GET6037;
            end if;
          else
            \$18805\ := work.Print.print_string(clk,of_string("racine:"));
            \$18806\ := work.Int.print(clk,\$18793_copy_root_in_ram6635879_arg\(0 to 15));
            \$18807\ := work.Print.print_newline(clk,eclat_unit);
            \$v6062\ := \$ram_lock\;
            if \$v6062\(0) = '1' then
              state_var7464 := Q_WAIT6061;
            else
              acquire(\$ram_lock\);
              \$ram_ptr\ <= to_integer(unsigned(\$18793_copy_root_in_ram6635879_arg\(0 to 15)));
              state_var7464 := PAUSE_GET6060;
            end if;
          end if;
        when PAUSE_GET5980 =>
          \$19213\ := \$ram_value\;
          release(\$ram_lock\);
          \$v5979\ := \$ram_lock\;
          if \$v5979\(0) = '1' then
            state_var7464 := Q_WAIT5978;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(\$18632_loop666_arg\(16 to 31), \$18632_loop666_arg\(0 to 15))));
            \$ram_write\ <= \$19213\; \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET5977;
          end if;
        when PAUSE_GET5996 =>
          \$19132_hd\ := \$ram_value\;
          release(\$ram_lock\);
          \$19136\ := work.Print.print_string(clk,of_string("bloc "));
          \$19137\ := work.Int.print(clk,eclat_resize(\$19111\(0 to 30),16));
          \$19138\ := work.Print.print_string(clk,of_string(" of size "));
          \$19139\ := work.Int.print(clk,work.Int.add(eclat_resize(work.Int.lsr(
                                                                   \$19132_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
          \$19140\ := work.Print.print_string(clk,of_string(" from "));
          \$19141\ := work.Int.print(clk,eclat_resize(\$19111\(0 to 30),16));
          \$19142\ := work.Print.print_string(clk,of_string(" to "));
          \$19143\ := work.Int.print(clk,\$18633_loop665_arg\(16 to 31));
          \$19144\ := work.Print.print_newline(clk,eclat_unit);
          \$v5995\ := \$ram_lock\;
          if \$v5995\(0) = '1' then
            state_var7464 := Q_WAIT5994;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(\$18633_loop665_arg\(16 to 31)));
            \$ram_write\ <= \$19132_hd\; \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET5993;
          end if;
        when PAUSE_GET6000 =>
          \$19127_w\ := \$ram_value\;
          release(\$ram_lock\);
          \$v5999\ := eclat_if(work.Bool.lnot(""&\$19127_w\(31)) & eclat_if(
                                                                   work.Int.le(
                                                                   \$18633_loop665_arg\(48 to 63), eclat_resize(\$19127_w\(0 to 30),16)) & 
                                                                   work.Int.lt(
                                                                   eclat_resize(\$19127_w\(0 to 30),16), 
                                                                   work.Int.add(
                                                                   \$18633_loop665_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false);
          if \$v5999\(0) = '1' then
            \$19115\ := \$19127_w\ & \$18633_loop665_arg\(16 to 31);
            \$v5986\ := \$ram_lock\;
            if \$v5986\(0) = '1' then
              state_var7464 := Q_WAIT5985;
            else
              acquire(\$ram_lock\);
              \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(\$18633_loop665_arg\(64 to 79), \$18633_loop665_arg\(0 to 15))));
              \$ram_write\ <= \$19115\(0 to 31); \$ram_write_request\ <= '1';
              state_var7464 := PAUSE_SET5984;
            end if;
          else
            \$v5998\ := \$ram_lock\;
            if \$v5998\(0) = '1' then
              state_var7464 := Q_WAIT5997;
            else
              acquire(\$ram_lock\);
              \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$19111\(0 to 30),16)));
              state_var7464 := PAUSE_GET5996;
            end if;
          end if;
        when PAUSE_GET6004 =>
          \$19111\ := \$ram_value\;
          release(\$ram_lock\);
          \$v6003\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$19111\(31)) & 
                                     eclat_if(work.Int.le(\$18633_loop665_arg\(32 to 47), eclat_resize(\$19111\(0 to 30),16)) & 
                                     work.Int.lt(eclat_resize(\$19111\(0 to 30),16), 
                                                 work.Int.add(\$18633_loop665_arg\(32 to 47), X"1770")) & eclat_false) & eclat_false));
          if \$v6003\(0) = '1' then
            \$19115\ := \$19111\ & \$18633_loop665_arg\(16 to 31);
            \$v5986\ := \$ram_lock\;
            if \$v5986\(0) = '1' then
              state_var7464 := Q_WAIT5985;
            else
              acquire(\$ram_lock\);
              \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(\$18633_loop665_arg\(64 to 79), \$18633_loop665_arg\(0 to 15))));
              \$ram_write\ <= \$19115\(0 to 31); \$ram_write_request\ <= '1';
              state_var7464 := PAUSE_SET5984;
            end if;
          else
            \$v6002\ := \$ram_lock\;
            if \$v6002\(0) = '1' then
              state_var7464 := Q_WAIT6001;
            else
              acquire(\$ram_lock\);
              \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19111\(0 to 30),16), X"000" & X"1")));
              state_var7464 := PAUSE_GET6000;
            end if;
          end if;
        when PAUSE_GET6008 =>
          \$19076\ := \$ram_value\;
          release(\$ram_lock\);
          \$18633_loop665_id\ := "000000000011";
          \$18633_loop665_arg\ := X"000" & X"1" & \$18634_aux664_arg\(16 to 31) & \$18634_aux664_arg\(32 to 47) & \$18634_aux664_arg\(48 to 63) & \$18634_aux664_arg\(0 to 15) & eclat_resize(
          work.Int.lsr(eclat_resize(eclat_resize(\$19076\(0 to 30),16),31), X"0000000" & X"2"),16);
          state_var7464 := \$18633_LOOP665\;
        when PAUSE_GET6025 =>
          \$18724_hd\ := \$ram_value\;
          release(\$ram_lock\);
          \$18728\ := work.Print.print_string(clk,of_string("bloc "));
          \$18729\ := work.Int.print(clk,eclat_resize(\$18701\(0 to 30),16));
          \$18730\ := work.Print.print_string(clk,of_string(" of size "));
          \$18731\ := work.Int.print(clk,work.Int.add(eclat_resize(work.Int.lsr(
                                                                   \$18724_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
          \$18732\ := work.Print.print_string(clk,of_string(" from "));
          \$18733\ := work.Int.print(clk,eclat_resize(\$18701\(0 to 30),16));
          \$18734\ := work.Print.print_string(clk,of_string(" to "));
          \$18735\ := work.Int.print(clk,\$18686_copy_root_in_ram6635880_arg\(32 to 47));
          \$18736\ := work.Print.print_newline(clk,eclat_unit);
          \$v6024\ := \$ram_lock\;
          if \$v6024\(0) = '1' then
            state_var7464 := Q_WAIT6023;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(\$18686_copy_root_in_ram6635880_arg\(32 to 47)));
            \$ram_write\ <= \$18724_hd\; \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET6022;
          end if;
        when PAUSE_GET6029 =>
          \$18719_w\ := \$ram_value\;
          release(\$ram_lock\);
          \$v6028\ := eclat_if(work.Bool.lnot(""&\$18719_w\(31)) & eclat_if(
                                                                   work.Int.le(
                                                                   \$18686_copy_root_in_ram6635880_arg\(64 to 79), eclat_resize(\$18719_w\(0 to 30),16)) & 
                                                                   work.Int.lt(
                                                                   eclat_resize(\$18719_w\(0 to 30),16), 
                                                                   work.Int.add(
                                                                   \$18686_copy_root_in_ram6635880_arg\(64 to 79), X"1770")) & eclat_false) & eclat_false);
          if \$v6028\(0) = '1' then
            \$18705\ := \$18719_w\ & \$18686_copy_root_in_ram6635880_arg\(32 to 47);
            \$v6015\ := \$ram_lock\;
            if \$v6015\(0) = '1' then
              state_var7464 := Q_WAIT6014;
            else
              acquire(\$ram_lock\);
              \$ram_ptr_write\ <= to_integer(unsigned(\$18686_copy_root_in_ram6635880_arg\(0 to 15)));
              \$ram_write\ <= \$18705\(0 to 31); \$ram_write_request\ <= '1';
              state_var7464 := PAUSE_SET6013;
            end if;
          else
            \$v6027\ := \$ram_lock\;
            if \$v6027\(0) = '1' then
              state_var7464 := Q_WAIT6026;
            else
              acquire(\$ram_lock\);
              \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18701\(0 to 30),16)));
              state_var7464 := PAUSE_GET6025;
            end if;
          end if;
        when PAUSE_GET6033 =>
          \$18701\ := \$ram_value\;
          release(\$ram_lock\);
          \$v6032\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$18701\(31)) & 
                                     eclat_if(work.Int.le(\$18686_copy_root_in_ram6635880_arg\(48 to 63), eclat_resize(\$18701\(0 to 30),16)) & 
                                     work.Int.lt(eclat_resize(\$18701\(0 to 30),16), 
                                                 work.Int.add(\$18686_copy_root_in_ram6635880_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false));
          if \$v6032\(0) = '1' then
            \$18705\ := \$18701\ & \$18686_copy_root_in_ram6635880_arg\(32 to 47);
            \$v6015\ := \$ram_lock\;
            if \$v6015\(0) = '1' then
              state_var7464 := Q_WAIT6014;
            else
              acquire(\$ram_lock\);
              \$ram_ptr_write\ <= to_integer(unsigned(\$18686_copy_root_in_ram6635880_arg\(0 to 15)));
              \$ram_write\ <= \$18705\(0 to 31); \$ram_write_request\ <= '1';
              state_var7464 := PAUSE_SET6013;
            end if;
          else
            \$v6031\ := \$ram_lock\;
            if \$v6031\(0) = '1' then
              state_var7464 := Q_WAIT6030;
            else
              acquire(\$ram_lock\);
              \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18701\(0 to 30),16), X"000" & X"1")));
              state_var7464 := PAUSE_GET6029;
            end if;
          end if;
        when PAUSE_GET6037 =>
          \$18665\ := \$global_end_value\;
          release(\$global_end_lock\);
          \$18686_copy_root_in_ram6635880_id\ := "000000000111";
          \$18686_copy_root_in_ram6635880_arg\ := X"3e80" & \$18665\ & \$18664_next\ & \$18621\(96 to 111) & \$18621\(112 to 127);
          state_var7464 := \$18686_COPY_ROOT_IN_RAM6635880\;
        when PAUSE_GET6052 =>
          \$18831_hd\ := \$ram_value\;
          release(\$ram_lock\);
          \$18835\ := work.Print.print_string(clk,of_string("bloc "));
          \$18836\ := work.Int.print(clk,eclat_resize(\$18808\(0 to 30),16));
          \$18837\ := work.Print.print_string(clk,of_string(" of size "));
          \$18838\ := work.Int.print(clk,work.Int.add(eclat_resize(work.Int.lsr(
                                                                   \$18831_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
          \$18839\ := work.Print.print_string(clk,of_string(" from "));
          \$18840\ := work.Int.print(clk,eclat_resize(\$18808\(0 to 30),16));
          \$18841\ := work.Print.print_string(clk,of_string(" to "));
          \$18842\ := work.Int.print(clk,\$18793_copy_root_in_ram6635879_arg\(32 to 47));
          \$18843\ := work.Print.print_newline(clk,eclat_unit);
          \$v6051\ := \$ram_lock\;
          if \$v6051\(0) = '1' then
            state_var7464 := Q_WAIT6050;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(\$18793_copy_root_in_ram6635879_arg\(32 to 47)));
            \$ram_write\ <= \$18831_hd\; \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET6049;
          end if;
        when PAUSE_GET6056 =>
          \$18826_w\ := \$ram_value\;
          release(\$ram_lock\);
          \$v6055\ := eclat_if(work.Bool.lnot(""&\$18826_w\(31)) & eclat_if(
                                                                   work.Int.le(
                                                                   \$18793_copy_root_in_ram6635879_arg\(64 to 79), eclat_resize(\$18826_w\(0 to 30),16)) & 
                                                                   work.Int.lt(
                                                                   eclat_resize(\$18826_w\(0 to 30),16), 
                                                                   work.Int.add(
                                                                   \$18793_copy_root_in_ram6635879_arg\(64 to 79), X"1770")) & eclat_false) & eclat_false);
          if \$v6055\(0) = '1' then
            \$18812\ := \$18826_w\ & \$18793_copy_root_in_ram6635879_arg\(32 to 47);
            \$v6042\ := \$ram_lock\;
            if \$v6042\(0) = '1' then
              state_var7464 := Q_WAIT6041;
            else
              acquire(\$ram_lock\);
              \$ram_ptr_write\ <= to_integer(unsigned(\$18793_copy_root_in_ram6635879_arg\(0 to 15)));
              \$ram_write\ <= \$18812\(0 to 31); \$ram_write_request\ <= '1';
              state_var7464 := PAUSE_SET6040;
            end if;
          else
            \$v6054\ := \$ram_lock\;
            if \$v6054\(0) = '1' then
              state_var7464 := Q_WAIT6053;
            else
              acquire(\$ram_lock\);
              \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18808\(0 to 30),16)));
              state_var7464 := PAUSE_GET6052;
            end if;
          end if;
        when PAUSE_GET6060 =>
          \$18808\ := \$ram_value\;
          release(\$ram_lock\);
          \$v6059\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$18808\(31)) & 
                                     eclat_if(work.Int.le(\$18793_copy_root_in_ram6635879_arg\(48 to 63), eclat_resize(\$18808\(0 to 30),16)) & 
                                     work.Int.lt(eclat_resize(\$18808\(0 to 30),16), 
                                                 work.Int.add(\$18793_copy_root_in_ram6635879_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false));
          if \$v6059\(0) = '1' then
            \$18812\ := \$18808\ & \$18793_copy_root_in_ram6635879_arg\(32 to 47);
            \$v6042\ := \$ram_lock\;
            if \$v6042\(0) = '1' then
              state_var7464 := Q_WAIT6041;
            else
              acquire(\$ram_lock\);
              \$ram_ptr_write\ <= to_integer(unsigned(\$18793_copy_root_in_ram6635879_arg\(0 to 15)));
              \$ram_write\ <= \$18812\(0 to 31); \$ram_write_request\ <= '1';
              state_var7464 := PAUSE_SET6040;
            end if;
          else
            \$v6058\ := \$ram_lock\;
            if \$v6058\(0) = '1' then
              state_var7464 := Q_WAIT6057;
            else
              acquire(\$ram_lock\);
              \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18808\(0 to 30),16), X"000" & X"1")));
              state_var7464 := PAUSE_GET6056;
            end if;
          end if;
        when PAUSE_GET6073 =>
          \$18909_hd\ := \$ram_value\;
          release(\$ram_lock\);
          \$18913\ := work.Print.print_string(clk,of_string("bloc "));
          \$18914\ := work.Int.print(clk,eclat_resize(\$12522_wait662_arg\(33 to 63),16));
          \$18915\ := work.Print.print_string(clk,of_string(" of size "));
          \$18916\ := work.Int.print(clk,work.Int.add(eclat_resize(work.Int.lsr(
                                                                   \$18909_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
          \$18917\ := work.Print.print_string(clk,of_string(" from "));
          \$18918\ := work.Int.print(clk,eclat_resize(\$12522_wait662_arg\(33 to 63),16));
          \$18919\ := work.Print.print_string(clk,of_string(" to "));
          \$18920\ := work.Int.print(clk,\$18644\(32 to 47));
          \$18921\ := work.Print.print_newline(clk,eclat_unit);
          \$v6072\ := \$ram_lock\;
          if \$v6072\(0) = '1' then
            state_var7464 := Q_WAIT6071;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(\$18644\(32 to 47)));
            \$ram_write\ <= \$18909_hd\; \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET6070;
          end if;
        when PAUSE_GET6077 =>
          \$18904_w\ := \$ram_value\;
          release(\$ram_lock\);
          \$v6076\ := eclat_if(work.Bool.lnot(""&\$18904_w\(31)) & eclat_if(
                                                                   work.Int.le(
                                                                   \$18621\(112 to 127), eclat_resize(\$18904_w\(0 to 30),16)) & 
                                                                   work.Int.lt(
                                                                   eclat_resize(\$18904_w\(0 to 30),16), 
                                                                   work.Int.add(
                                                                   \$18621\(112 to 127), X"1770")) & eclat_false) & eclat_false);
          if \$v6076\(0) = '1' then
            \$18661\ := \$18904_w\ & \$18644\(32 to 47);
            \$18793_copy_root_in_ram6635879_id\ := "000000001001";
            \$18793_copy_root_in_ram6635879_arg\ := X"0" & X"3e8" & \$12522_wait662_arg\(65 to 80) & \$18661\(32 to 47) & \$18621\(96 to 111) & \$18621\(112 to 127);
            state_var7464 := \$18793_COPY_ROOT_IN_RAM6635879\;
          else
            \$v6075\ := \$ram_lock\;
            if \$v6075\(0) = '1' then
              state_var7464 := Q_WAIT6074;
            else
              acquire(\$ram_lock\);
              \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$12522_wait662_arg\(33 to 63),16)));
              state_var7464 := PAUSE_GET6073;
            end if;
          end if;
        when PAUSE_GET6090 =>
          \$18987_hd\ := \$ram_value\;
          release(\$ram_lock\);
          \$18991\ := work.Print.print_string(clk,of_string("bloc "));
          \$18992\ := work.Int.print(clk,eclat_resize(\$12522_wait662_arg\(1 to 31),16));
          \$18993\ := work.Print.print_string(clk,of_string(" of size "));
          \$18994\ := work.Int.print(clk,work.Int.add(eclat_resize(work.Int.lsr(
                                                                   \$18987_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
          \$18995\ := work.Print.print_string(clk,of_string(" from "));
          \$18996\ := work.Int.print(clk,eclat_resize(\$12522_wait662_arg\(1 to 31),16));
          \$18997\ := work.Print.print_string(clk,of_string(" to "));
          \$18998\ := work.Int.print(clk,\$18621\(112 to 127));
          \$18999\ := work.Print.print_newline(clk,eclat_unit);
          \$v6089\ := \$ram_lock\;
          if \$v6089\(0) = '1' then
            state_var7464 := Q_WAIT6088;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(\$18621\(112 to 127)));
            \$ram_write\ <= \$18987_hd\; \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET6087;
          end if;
        when PAUSE_GET6094 =>
          \$18982_w\ := \$ram_value\;
          release(\$ram_lock\);
          \$v6093\ := eclat_if(work.Bool.lnot(""&\$18982_w\(31)) & eclat_if(
                                                                   work.Int.le(
                                                                   \$18621\(112 to 127), eclat_resize(\$18982_w\(0 to 30),16)) & 
                                                                   work.Int.lt(
                                                                   eclat_resize(\$18982_w\(0 to 30),16), 
                                                                   work.Int.add(
                                                                   \$18621\(112 to 127), X"1770")) & eclat_false) & eclat_false);
          if \$v6093\(0) = '1' then
            \$18644\ := \$18982_w\ & \$18621\(112 to 127);
            \$v6080\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$12522_wait662_arg\(64)) & 
                                       eclat_if(work.Int.le(\$18621\(96 to 111), eclat_resize(\$12522_wait662_arg\(33 to 63),16)) & 
                                       work.Int.lt(eclat_resize(\$12522_wait662_arg\(33 to 63),16), 
                                                   work.Int.add(\$18621\(96 to 111), X"1770")) & eclat_false) & eclat_false));
            if \$v6080\(0) = '1' then
              \$18661\ := \$12522_wait662_arg\(33 to 64) & \$18644\(32 to 47);
              \$18793_copy_root_in_ram6635879_id\ := "000000001001";
              \$18793_copy_root_in_ram6635879_arg\ := X"0" & X"3e8" & \$12522_wait662_arg\(65 to 80) & \$18661\(32 to 47) & \$18621\(96 to 111) & \$18621\(112 to 127);
              state_var7464 := \$18793_COPY_ROOT_IN_RAM6635879\;
            else
              \$v6079\ := \$ram_lock\;
              if \$v6079\(0) = '1' then
                state_var7464 := Q_WAIT6078;
              else
                acquire(\$ram_lock\);
                \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$12522_wait662_arg\(33 to 63),16), X"000" & X"1")));
                state_var7464 := PAUSE_GET6077;
              end if;
            end if;
          else
            \$v6092\ := \$ram_lock\;
            if \$v6092\(0) = '1' then
              state_var7464 := Q_WAIT6091;
            else
              acquire(\$ram_lock\);
              \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$12522_wait662_arg\(1 to 31),16)));
              state_var7464 := PAUSE_GET6090;
            end if;
          end if;
        when PAUSE_SET5977 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$19214\ := eclat_unit;
          \$18632_loop666_arg\ := work.Int.add(\$18632_loop666_arg\(0 to 15), X"000" & X"1") & \$18632_loop666_arg\(16 to 31) & \$18632_loop666_arg\(32 to 47) & \$18632_loop666_arg\(48 to 63);
          state_var7464 := \$18632_LOOP666\;
        when PAUSE_SET5984 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$19118\ := eclat_unit;
          \$18633_loop665_arg\ := work.Int.add(\$18633_loop665_arg\(0 to 15), X"000" & X"1") & \$19115\(32 to 47) & \$18633_loop665_arg\(32 to 47) & \$18633_loop665_arg\(48 to 63) & \$18633_loop665_arg\(64 to 79) & \$18633_loop665_arg\(80 to 95);
          state_var7464 := \$18633_LOOP665\;
        when PAUSE_SET5987 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$19148\ := eclat_unit;
          \$19115\ := eclat_resize(\$18633_loop665_arg\(16 to 31),31) & eclat_false & 
          work.Int.add(\$18633_loop665_arg\(16 to 31), work.Int.add(eclat_resize(
                                                                    work.Int.lsr(
                                                                    \$19132_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
          \$v5986\ := \$ram_lock\;
          if \$v5986\(0) = '1' then
            state_var7464 := Q_WAIT5985;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(\$18633_loop665_arg\(64 to 79), \$18633_loop665_arg\(0 to 15))));
            \$ram_write\ <= \$19115\(0 to 31); \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET5984;
          end if;
        when PAUSE_SET5990 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$19147\ := eclat_unit;
          \$v5989\ := \$ram_lock\;
          if \$v5989\(0) = '1' then
            state_var7464 := Q_WAIT5988;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19111\(0 to 30),16), X"000" & X"1")));
            \$ram_write\ <= eclat_resize(\$18633_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET5987;
          end if;
        when PAUSE_SET5993 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$19145\ := eclat_unit;
          \$18632_loop666_id\ := "000000000010";
          \$18632_loop666_arg\ := X"000" & X"1" & \$18633_loop665_arg\(16 to 31) & eclat_resize(\$19111\(0 to 30),16) & eclat_resize(
          work.Int.lsr(\$19132_hd\(0 to 30), X"0000000" & X"2"),16);
          state_var7464 := \$18632_LOOP666\;
        when PAUSE_SET6013 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$18708\ := eclat_unit;
          \$18709\ := work.Print.print_string(clk,of_string(" next="));
          \$18710\ := work.Int.print(clk,\$18705\(32 to 47));
          \$18711\ := work.Print.print_newline(clk,eclat_unit);
          \$18686_copy_root_in_ram6635880_arg\ := work.Int.add(\$18686_copy_root_in_ram6635880_arg\(0 to 15), X"000" & X"1") & \$18686_copy_root_in_ram6635880_arg\(16 to 31) & \$18705\(32 to 47) & \$18686_copy_root_in_ram6635880_arg\(48 to 63) & \$18686_copy_root_in_ram6635880_arg\(64 to 79);
          state_var7464 := \$18686_COPY_ROOT_IN_RAM6635880\;
        when PAUSE_SET6016 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$18740\ := eclat_unit;
          \$18705\ := eclat_resize(\$18686_copy_root_in_ram6635880_arg\(32 to 47),31) & eclat_false & 
          work.Int.add(\$18686_copy_root_in_ram6635880_arg\(32 to 47), 
                       work.Int.add(eclat_resize(work.Int.lsr(\$18724_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
          \$v6015\ := \$ram_lock\;
          if \$v6015\(0) = '1' then
            state_var7464 := Q_WAIT6014;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(\$18686_copy_root_in_ram6635880_arg\(0 to 15)));
            \$ram_write\ <= \$18705\(0 to 31); \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET6013;
          end if;
        when PAUSE_SET6019 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$18739\ := eclat_unit;
          \$v6018\ := \$ram_lock\;
          if \$v6018\(0) = '1' then
            state_var7464 := Q_WAIT6017;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18701\(0 to 30),16), X"000" & X"1")));
            \$ram_write\ <= eclat_resize(\$18686_copy_root_in_ram6635880_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET6016;
          end if;
        when PAUSE_SET6022 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$18737\ := eclat_unit;
          \$18632_loop666_id\ := "000000000110";
          \$18632_loop666_arg\ := X"000" & X"1" & \$18686_copy_root_in_ram6635880_arg\(32 to 47) & eclat_resize(\$18701\(0 to 30),16) & eclat_resize(
          work.Int.lsr(\$18724_hd\(0 to 30), X"0000000" & X"2"),16);
          state_var7464 := \$18632_LOOP666\;
        when PAUSE_SET6040 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$18815\ := eclat_unit;
          \$18816\ := work.Print.print_string(clk,of_string(" next="));
          \$18817\ := work.Int.print(clk,\$18812\(32 to 47));
          \$18818\ := work.Print.print_newline(clk,eclat_unit);
          \$18793_copy_root_in_ram6635879_arg\ := work.Int.add(\$18793_copy_root_in_ram6635879_arg\(0 to 15), X"000" & X"1") & \$18793_copy_root_in_ram6635879_arg\(16 to 31) & \$18812\(32 to 47) & \$18793_copy_root_in_ram6635879_arg\(48 to 63) & \$18793_copy_root_in_ram6635879_arg\(64 to 79);
          state_var7464 := \$18793_COPY_ROOT_IN_RAM6635879\;
        when PAUSE_SET6043 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$18847\ := eclat_unit;
          \$18812\ := eclat_resize(\$18793_copy_root_in_ram6635879_arg\(32 to 47),31) & eclat_false & 
          work.Int.add(\$18793_copy_root_in_ram6635879_arg\(32 to 47), 
                       work.Int.add(eclat_resize(work.Int.lsr(\$18831_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
          \$v6042\ := \$ram_lock\;
          if \$v6042\(0) = '1' then
            state_var7464 := Q_WAIT6041;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(\$18793_copy_root_in_ram6635879_arg\(0 to 15)));
            \$ram_write\ <= \$18812\(0 to 31); \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET6040;
          end if;
        when PAUSE_SET6046 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$18846\ := eclat_unit;
          \$v6045\ := \$ram_lock\;
          if \$v6045\(0) = '1' then
            state_var7464 := Q_WAIT6044;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18808\(0 to 30),16), X"000" & X"1")));
            \$ram_write\ <= eclat_resize(\$18793_copy_root_in_ram6635879_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET6043;
          end if;
        when PAUSE_SET6049 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$18844\ := eclat_unit;
          \$18632_loop666_id\ := "000000001000";
          \$18632_loop666_arg\ := X"000" & X"1" & \$18793_copy_root_in_ram6635879_arg\(32 to 47) & eclat_resize(\$18808\(0 to 30),16) & eclat_resize(
          work.Int.lsr(\$18831_hd\(0 to 30), X"0000000" & X"2"),16);
          state_var7464 := \$18632_LOOP666\;
        when PAUSE_SET6064 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$18925\ := eclat_unit;
          \$18661\ := eclat_resize(\$18644\(32 to 47),31) & eclat_false & 
          work.Int.add(\$18644\(32 to 47), work.Int.add(eclat_resize(
                                                        work.Int.lsr(
                                                        \$18909_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
          \$18793_copy_root_in_ram6635879_id\ := "000000001001";
          \$18793_copy_root_in_ram6635879_arg\ := X"0" & X"3e8" & \$12522_wait662_arg\(65 to 80) & \$18661\(32 to 47) & \$18621\(96 to 111) & \$18621\(112 to 127);
          state_var7464 := \$18793_COPY_ROOT_IN_RAM6635879\;
        when PAUSE_SET6067 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$18924\ := eclat_unit;
          \$v6066\ := \$ram_lock\;
          if \$v6066\(0) = '1' then
            state_var7464 := Q_WAIT6065;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$12522_wait662_arg\(33 to 63),16), X"000" & X"1")));
            \$ram_write\ <= eclat_resize(\$18644\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET6064;
          end if;
        when PAUSE_SET6070 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$18922\ := eclat_unit;
          \$18632_loop666_id\ := "000000001010";
          \$18632_loop666_arg\ := X"000" & X"1" & \$18644\(32 to 47) & eclat_resize(\$12522_wait662_arg\(33 to 63),16) & eclat_resize(
          work.Int.lsr(\$18909_hd\(0 to 30), X"0000000" & X"2"),16);
          state_var7464 := \$18632_LOOP666\;
        when PAUSE_SET6081 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$19003\ := eclat_unit;
          \$18644\ := eclat_resize(\$18621\(112 to 127),31) & eclat_false & 
          work.Int.add(\$18621\(112 to 127), work.Int.add(eclat_resize(
                                                          work.Int.lsr(
                                                          \$18987_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
          \$v6080\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$12522_wait662_arg\(64)) & 
                                     eclat_if(work.Int.le(\$18621\(96 to 111), eclat_resize(\$12522_wait662_arg\(33 to 63),16)) & 
                                     work.Int.lt(eclat_resize(\$12522_wait662_arg\(33 to 63),16), 
                                                 work.Int.add(\$18621\(96 to 111), X"1770")) & eclat_false) & eclat_false));
          if \$v6080\(0) = '1' then
            \$18661\ := \$12522_wait662_arg\(33 to 64) & \$18644\(32 to 47);
            \$18793_copy_root_in_ram6635879_id\ := "000000001001";
            \$18793_copy_root_in_ram6635879_arg\ := X"0" & X"3e8" & \$12522_wait662_arg\(65 to 80) & \$18661\(32 to 47) & \$18621\(96 to 111) & \$18621\(112 to 127);
            state_var7464 := \$18793_COPY_ROOT_IN_RAM6635879\;
          else
            \$v6079\ := \$ram_lock\;
            if \$v6079\(0) = '1' then
              state_var7464 := Q_WAIT6078;
            else
              acquire(\$ram_lock\);
              \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$12522_wait662_arg\(33 to 63),16), X"000" & X"1")));
              state_var7464 := PAUSE_GET6077;
            end if;
          end if;
        when PAUSE_SET6084 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$19002\ := eclat_unit;
          \$v6083\ := \$ram_lock\;
          if \$v6083\(0) = '1' then
            state_var7464 := Q_WAIT6082;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$12522_wait662_arg\(1 to 31),16), X"000" & X"1")));
            \$ram_write\ <= eclat_resize(\$18621\(112 to 127),31) & eclat_false; \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET6081;
          end if;
        when PAUSE_SET6087 =>
          \$ram_write_request\ <= '0';
          release(\$ram_lock\);
          \$19000\ := eclat_unit;
          \$18632_loop666_id\ := "000000001011";
          \$18632_loop666_arg\ := X"000" & X"1" & \$18621\(112 to 127) & eclat_resize(\$12522_wait662_arg\(1 to 31),16) & eclat_resize(
          work.Int.lsr(\$18987_hd\(0 to 30), X"0000000" & X"2"),16);
          state_var7464 := \$18632_LOOP666\;
        when Q_WAIT5978 =>
          \$v5979\ := \$ram_lock\;
          if \$v5979\(0) = '1' then
            state_var7464 := Q_WAIT5978;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(\$18632_loop666_arg\(16 to 31), \$18632_loop666_arg\(0 to 15))));
            \$ram_write\ <= \$19213\; \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET5977;
          end if;
        when Q_WAIT5981 =>
          \$v5982\ := \$ram_lock\;
          if \$v5982\(0) = '1' then
            state_var7464 := Q_WAIT5981;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$18632_loop666_arg\(32 to 47), \$18632_loop666_arg\(0 to 15))));
            state_var7464 := PAUSE_GET5980;
          end if;
        when Q_WAIT5985 =>
          \$v5986\ := \$ram_lock\;
          if \$v5986\(0) = '1' then
            state_var7464 := Q_WAIT5985;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(\$18633_loop665_arg\(64 to 79), \$18633_loop665_arg\(0 to 15))));
            \$ram_write\ <= \$19115\(0 to 31); \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET5984;
          end if;
        when Q_WAIT5988 =>
          \$v5989\ := \$ram_lock\;
          if \$v5989\(0) = '1' then
            state_var7464 := Q_WAIT5988;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19111\(0 to 30),16), X"000" & X"1")));
            \$ram_write\ <= eclat_resize(\$18633_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET5987;
          end if;
        when Q_WAIT5991 =>
          \$v5992\ := \$ram_lock\;
          if \$v5992\(0) = '1' then
            state_var7464 := Q_WAIT5991;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$19111\(0 to 30),16)));
            \$ram_write\ <= eclat_resize(\$18633_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET5990;
          end if;
        when Q_WAIT5994 =>
          \$v5995\ := \$ram_lock\;
          if \$v5995\(0) = '1' then
            state_var7464 := Q_WAIT5994;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(\$18633_loop665_arg\(16 to 31)));
            \$ram_write\ <= \$19132_hd\; \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET5993;
          end if;
        when Q_WAIT5997 =>
          \$v5998\ := \$ram_lock\;
          if \$v5998\(0) = '1' then
            state_var7464 := Q_WAIT5997;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$19111\(0 to 30),16)));
            state_var7464 := PAUSE_GET5996;
          end if;
        when Q_WAIT6001 =>
          \$v6002\ := \$ram_lock\;
          if \$v6002\(0) = '1' then
            state_var7464 := Q_WAIT6001;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19111\(0 to 30),16), X"000" & X"1")));
            state_var7464 := PAUSE_GET6000;
          end if;
        when Q_WAIT6005 =>
          \$v6006\ := \$ram_lock\;
          if \$v6006\(0) = '1' then
            state_var7464 := Q_WAIT6005;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$18633_loop665_arg\(64 to 79), \$18633_loop665_arg\(0 to 15))));
            state_var7464 := PAUSE_GET6004;
          end if;
        when Q_WAIT6009 =>
          \$v6010\ := \$ram_lock\;
          if \$v6010\(0) = '1' then
            state_var7464 := Q_WAIT6009;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(\$18634_aux664_arg\(0 to 15)));
            state_var7464 := PAUSE_GET6008;
          end if;
        when Q_WAIT6014 =>
          \$v6015\ := \$ram_lock\;
          if \$v6015\(0) = '1' then
            state_var7464 := Q_WAIT6014;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(\$18686_copy_root_in_ram6635880_arg\(0 to 15)));
            \$ram_write\ <= \$18705\(0 to 31); \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET6013;
          end if;
        when Q_WAIT6017 =>
          \$v6018\ := \$ram_lock\;
          if \$v6018\(0) = '1' then
            state_var7464 := Q_WAIT6017;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18701\(0 to 30),16), X"000" & X"1")));
            \$ram_write\ <= eclat_resize(\$18686_copy_root_in_ram6635880_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET6016;
          end if;
        when Q_WAIT6020 =>
          \$v6021\ := \$ram_lock\;
          if \$v6021\(0) = '1' then
            state_var7464 := Q_WAIT6020;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18701\(0 to 30),16)));
            \$ram_write\ <= eclat_resize(\$18686_copy_root_in_ram6635880_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET6019;
          end if;
        when Q_WAIT6023 =>
          \$v6024\ := \$ram_lock\;
          if \$v6024\(0) = '1' then
            state_var7464 := Q_WAIT6023;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(\$18686_copy_root_in_ram6635880_arg\(32 to 47)));
            \$ram_write\ <= \$18724_hd\; \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET6022;
          end if;
        when Q_WAIT6026 =>
          \$v6027\ := \$ram_lock\;
          if \$v6027\(0) = '1' then
            state_var7464 := Q_WAIT6026;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18701\(0 to 30),16)));
            state_var7464 := PAUSE_GET6025;
          end if;
        when Q_WAIT6030 =>
          \$v6031\ := \$ram_lock\;
          if \$v6031\(0) = '1' then
            state_var7464 := Q_WAIT6030;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18701\(0 to 30),16), X"000" & X"1")));
            state_var7464 := PAUSE_GET6029;
          end if;
        when Q_WAIT6034 =>
          \$v6035\ := \$ram_lock\;
          if \$v6035\(0) = '1' then
            state_var7464 := Q_WAIT6034;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(\$18686_copy_root_in_ram6635880_arg\(0 to 15)));
            state_var7464 := PAUSE_GET6033;
          end if;
        when Q_WAIT6038 =>
          \$v6039\ := \$global_end_lock\;
          if \$v6039\(0) = '1' then
            state_var7464 := Q_WAIT6038;
          else
            acquire(\$global_end_lock\);
            \$global_end_ptr\ <= 0;
            state_var7464 := PAUSE_GET6037;
          end if;
        when Q_WAIT6041 =>
          \$v6042\ := \$ram_lock\;
          if \$v6042\(0) = '1' then
            state_var7464 := Q_WAIT6041;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(\$18793_copy_root_in_ram6635879_arg\(0 to 15)));
            \$ram_write\ <= \$18812\(0 to 31); \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET6040;
          end if;
        when Q_WAIT6044 =>
          \$v6045\ := \$ram_lock\;
          if \$v6045\(0) = '1' then
            state_var7464 := Q_WAIT6044;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18808\(0 to 30),16), X"000" & X"1")));
            \$ram_write\ <= eclat_resize(\$18793_copy_root_in_ram6635879_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET6043;
          end if;
        when Q_WAIT6047 =>
          \$v6048\ := \$ram_lock\;
          if \$v6048\(0) = '1' then
            state_var7464 := Q_WAIT6047;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18808\(0 to 30),16)));
            \$ram_write\ <= eclat_resize(\$18793_copy_root_in_ram6635879_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET6046;
          end if;
        when Q_WAIT6050 =>
          \$v6051\ := \$ram_lock\;
          if \$v6051\(0) = '1' then
            state_var7464 := Q_WAIT6050;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(\$18793_copy_root_in_ram6635879_arg\(32 to 47)));
            \$ram_write\ <= \$18831_hd\; \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET6049;
          end if;
        when Q_WAIT6053 =>
          \$v6054\ := \$ram_lock\;
          if \$v6054\(0) = '1' then
            state_var7464 := Q_WAIT6053;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18808\(0 to 30),16)));
            state_var7464 := PAUSE_GET6052;
          end if;
        when Q_WAIT6057 =>
          \$v6058\ := \$ram_lock\;
          if \$v6058\(0) = '1' then
            state_var7464 := Q_WAIT6057;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18808\(0 to 30),16), X"000" & X"1")));
            state_var7464 := PAUSE_GET6056;
          end if;
        when Q_WAIT6061 =>
          \$v6062\ := \$ram_lock\;
          if \$v6062\(0) = '1' then
            state_var7464 := Q_WAIT6061;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(\$18793_copy_root_in_ram6635879_arg\(0 to 15)));
            state_var7464 := PAUSE_GET6060;
          end if;
        when Q_WAIT6065 =>
          \$v6066\ := \$ram_lock\;
          if \$v6066\(0) = '1' then
            state_var7464 := Q_WAIT6065;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$12522_wait662_arg\(33 to 63),16), X"000" & X"1")));
            \$ram_write\ <= eclat_resize(\$18644\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET6064;
          end if;
        when Q_WAIT6068 =>
          \$v6069\ := \$ram_lock\;
          if \$v6069\(0) = '1' then
            state_var7464 := Q_WAIT6068;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$12522_wait662_arg\(33 to 63),16)));
            \$ram_write\ <= eclat_resize(\$18644\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET6067;
          end if;
        when Q_WAIT6071 =>
          \$v6072\ := \$ram_lock\;
          if \$v6072\(0) = '1' then
            state_var7464 := Q_WAIT6071;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(\$18644\(32 to 47)));
            \$ram_write\ <= \$18909_hd\; \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET6070;
          end if;
        when Q_WAIT6074 =>
          \$v6075\ := \$ram_lock\;
          if \$v6075\(0) = '1' then
            state_var7464 := Q_WAIT6074;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$12522_wait662_arg\(33 to 63),16)));
            state_var7464 := PAUSE_GET6073;
          end if;
        when Q_WAIT6078 =>
          \$v6079\ := \$ram_lock\;
          if \$v6079\(0) = '1' then
            state_var7464 := Q_WAIT6078;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$12522_wait662_arg\(33 to 63),16), X"000" & X"1")));
            state_var7464 := PAUSE_GET6077;
          end if;
        when Q_WAIT6082 =>
          \$v6083\ := \$ram_lock\;
          if \$v6083\(0) = '1' then
            state_var7464 := Q_WAIT6082;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$12522_wait662_arg\(1 to 31),16), X"000" & X"1")));
            \$ram_write\ <= eclat_resize(\$18621\(112 to 127),31) & eclat_false; \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET6081;
          end if;
        when Q_WAIT6085 =>
          \$v6086\ := \$ram_lock\;
          if \$v6086\(0) = '1' then
            state_var7464 := Q_WAIT6085;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$12522_wait662_arg\(1 to 31),16)));
            \$ram_write\ <= eclat_resize(\$18621\(112 to 127),31) & eclat_false; \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET6084;
          end if;
        when Q_WAIT6088 =>
          \$v6089\ := \$ram_lock\;
          if \$v6089\(0) = '1' then
            state_var7464 := Q_WAIT6088;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(\$18621\(112 to 127)));
            \$ram_write\ <= \$18987_hd\; \$ram_write_request\ <= '1';
            state_var7464 := PAUSE_SET6087;
          end if;
        when Q_WAIT6091 =>
          \$v6092\ := \$ram_lock\;
          if \$v6092\(0) = '1' then
            state_var7464 := Q_WAIT6091;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$12522_wait662_arg\(1 to 31),16)));
            state_var7464 := PAUSE_GET6090;
          end if;
        when Q_WAIT6095 =>
          \$v6096\ := \$ram_lock\;
          if \$v6096\(0) = '1' then
            state_var7464 := Q_WAIT6095;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$12522_wait662_arg\(1 to 31),16), X"000" & X"1")));
            state_var7464 := PAUSE_GET6094;
          end if;
        when IDLE5976 =>
          rdy5975 := eclat_false;
          \$v6098\ := work.Int.gt(work.Int.add(\$18621\(80 to 95), \$12522_wait662_arg\(81 to 96)), 
                                  work.Int.add(\$18621\(96 to 111), X"1770"));
          if \$v6098\(0) = '1' then
            \$18637\ := work.Print.print_newline(clk,eclat_unit);
            \$18638\ := work.Print.print_newline(clk,eclat_unit);
            \$18639\ := work.Print.print_string(clk,of_string("[================= GC START ======================]"));
            \$19056\ := work.Print.print_newline(clk,eclat_unit);
            \$18640\ := work.Print.print_newline(clk,eclat_unit);
            \$v6097\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$12522_wait662_arg\(32)) & 
                                       eclat_if(work.Int.le(\$18621\(96 to 111), eclat_resize(\$12522_wait662_arg\(1 to 31),16)) & 
                                       work.Int.lt(eclat_resize(\$12522_wait662_arg\(1 to 31),16), 
                                                   work.Int.add(\$18621\(96 to 111), X"1770")) & eclat_false) & eclat_false));
            if \$v6097\(0) = '1' then
              \$18644\ := \$12522_wait662_arg\(1 to 32) & \$18621\(112 to 127);
              \$v6080\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$12522_wait662_arg\(64)) & 
                                         eclat_if(work.Int.le(\$18621\(96 to 111), eclat_resize(\$12522_wait662_arg\(33 to 63),16)) & 
                                         work.Int.lt(eclat_resize(\$12522_wait662_arg\(33 to 63),16), 
                                                     work.Int.add(\$18621\(96 to 111), X"1770")) & eclat_false) & eclat_false));
              if \$v6080\(0) = '1' then
                \$18661\ := \$12522_wait662_arg\(33 to 64) & \$18644\(32 to 47);
                \$18793_copy_root_in_ram6635879_id\ := "000000001001";
                \$18793_copy_root_in_ram6635879_arg\ := X"0" & X"3e8" & \$12522_wait662_arg\(65 to 80) & \$18661\(32 to 47) & \$18621\(96 to 111) & \$18621\(112 to 127);
                state_var7464 := \$18793_COPY_ROOT_IN_RAM6635879\;
              else
                \$v6079\ := \$ram_lock\;
                if \$v6079\(0) = '1' then
                  state_var7464 := Q_WAIT6078;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$12522_wait662_arg\(33 to 63),16), X"000" & X"1")));
                  state_var7464 := PAUSE_GET6077;
                end if;
              end if;
            else
              \$v6096\ := \$ram_lock\;
              if \$v6096\(0) = '1' then
                state_var7464 := Q_WAIT6095;
              else
                acquire(\$ram_lock\);
                \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$12522_wait662_arg\(1 to 31),16), X"000" & X"1")));
                state_var7464 := PAUSE_GET6094;
              end if;
            end if;
          else
            result5974 := \$12522_wait662_arg\(1 to 32) & \$12522_wait662_arg\(33 to 64) & \$18621\(80 to 95) & 
            work.Int.add(\$18621\(80 to 95), \$12522_wait662_arg\(81 to 96)) & \$18621\(96 to 111) & \$18621\(112 to 127);
            rdy5975 := eclat_true;
            state_var7464 := IDLE5976;
          end if;
        end case;
        
        if rdy5975(0) = '1' then
          
        else
          result5974 := \$18621\(0 to 31) & \$18621\(32 to 63) & \$18621\(64 to 79) & \$18621\(80 to 95) & \$18621\(96 to 111) & \$18621\(112 to 127);
        end if;
        \$18621\ := result5974 & rdy5975;
        \$18611\ := \$18621\;
        \$v5973\ := ""&\$18611\(128);
        if \$v5973\(0) = '1' then
          \$12522_wait662_result\ := \$18611\(0 to 31) & \$18611\(32 to 63) & \$18611\(64 to 79);
          \$18566\ := \$12522_wait662_result\;
          \$18570\ := work.Print.print_string(clk,of_string("size:"));
          \$18571\ := work.Int.print(clk,eclat_if(work.Int.eq(\$12523_make_block579_arg\(112 to 127), X"000" & X"0") & X"000" & X"1" & \$12523_make_block579_arg\(112 to 127)));
          \$18572\ := work.Print.print_newline(clk,eclat_unit);
          \$v6102\ := \$ram_lock\;
          if \$v6102\(0) = '1' then
            state := Q_WAIT6101;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(\$18566\(64 to 79)));
            \$ram_write\ <= work.Int.lor(work.Int.lsl(eclat_resize(\$12523_make_block579_arg\(80 to 111),31), X"000000" & X"18"), 
                                         work.Int.lsl(eclat_resize(eclat_if(
                                                                   work.Int.eq(
                                                                   \$12523_make_block579_arg\(112 to 127), X"000" & X"0") & X"000" & X"1" & \$12523_make_block579_arg\(112 to 127)),31), X"0000000" & X"2")) & eclat_true; \$ram_write_request\ <= '1';
            state := PAUSE_SET6100;
          end if;
        else
          \$12522_wait662_arg\ := eclat_unit & \$12522_wait662_arg\(1 to 32) & \$12522_wait662_arg\(33 to 64) & \$12522_wait662_arg\(65 to 80) & \$12522_wait662_arg\(81 to 96);
          state := \$12522_WAIT662\;
        end if;
      when \$12523_MAKE_BLOCK579\ =>
        \$18563\ := work.Print.print_string(clk,of_string("GC-ALLOC:(size="));
        \$18564\ := work.Int.print(clk,work.Int.add(eclat_if(work.Int.eq(
                                                             \$12523_make_block579_arg\(112 to 127), X"000" & X"0") & X"000" & X"1" & \$12523_make_block579_arg\(112 to 127)), X"000" & X"1"));
        \$18565\ := work.Print.print_string(clk,of_string(")"));
        \$18589\ := work.Print.print_newline(clk,eclat_unit);
        \$12522_wait662_id\ := "000000001100";
        \$12522_wait662_arg\ := eclat_unit & \$12523_make_block579_arg\(16 to 47) & \$12523_make_block579_arg\(48 to 79) & \$12523_make_block579_arg\(0 to 15) & 
        work.Int.add(eclat_if(work.Int.eq(\$12523_make_block579_arg\(112 to 127), X"000" & X"0") & X"000" & X"1" & \$12523_make_block579_arg\(112 to 127)), X"000" & X"1");
        state := \$12522_WAIT662\;
      when PAUSE_GET5945 =>
        \$19337\ := \$ram_value\;
        release(\$ram_lock\);
        \$v5944\ := \$ram_lock\;
        if \$v5944\(0) = '1' then
          state := Q_WAIT5943;
        else
          acquire(\$ram_lock\);
          \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(\$12520_loop666_arg\(16 to 31), \$12520_loop666_arg\(0 to 15))));
          \$ram_write\ <= \$19337\; \$ram_write_request\ <= '1';
          state := PAUSE_SET5942;
        end if;
      when PAUSE_GET5961 =>
        \$19256_hd\ := \$ram_value\;
        release(\$ram_lock\);
        \$19260\ := work.Print.print_string(clk,of_string("bloc "));
        \$19261\ := work.Int.print(clk,eclat_resize(\$19235\(0 to 30),16));
        \$19262\ := work.Print.print_string(clk,of_string(" of size "));
        \$19263\ := work.Int.print(clk,work.Int.add(eclat_resize(work.Int.lsr(
                                                                 \$19256_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
        \$19264\ := work.Print.print_string(clk,of_string(" from "));
        \$19265\ := work.Int.print(clk,eclat_resize(\$19235\(0 to 30),16));
        \$19266\ := work.Print.print_string(clk,of_string(" to "));
        \$19267\ := work.Int.print(clk,\$12521_loop665_arg\(16 to 31));
        \$19268\ := work.Print.print_newline(clk,eclat_unit);
        \$v5960\ := \$ram_lock\;
        if \$v5960\(0) = '1' then
          state := Q_WAIT5959;
        else
          acquire(\$ram_lock\);
          \$ram_ptr_write\ <= to_integer(unsigned(\$12521_loop665_arg\(16 to 31)));
          \$ram_write\ <= \$19256_hd\; \$ram_write_request\ <= '1';
          state := PAUSE_SET5958;
        end if;
      when PAUSE_GET5965 =>
        \$19251_w\ := \$ram_value\;
        release(\$ram_lock\);
        \$v5964\ := eclat_if(work.Bool.lnot(""&\$19251_w\(31)) & eclat_if(
                                                                 work.Int.le(
                                                                 \$12521_loop665_arg\(48 to 63), eclat_resize(\$19251_w\(0 to 30),16)) & 
                                                                 work.Int.lt(
                                                                 eclat_resize(\$19251_w\(0 to 30),16), 
                                                                 work.Int.add(
                                                                 \$12521_loop665_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false);
        if \$v5964\(0) = '1' then
          \$19239\ := \$19251_w\ & \$12521_loop665_arg\(16 to 31);
          \$v5951\ := \$ram_lock\;
          if \$v5951\(0) = '1' then
            state := Q_WAIT5950;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(\$12521_loop665_arg\(64 to 79), \$12521_loop665_arg\(0 to 15))));
            \$ram_write\ <= \$19239\(0 to 31); \$ram_write_request\ <= '1';
            state := PAUSE_SET5949;
          end if;
        else
          \$v5963\ := \$ram_lock\;
          if \$v5963\(0) = '1' then
            state := Q_WAIT5962;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$19235\(0 to 30),16)));
            state := PAUSE_GET5961;
          end if;
        end if;
      when PAUSE_GET5969 =>
        \$19235\ := \$ram_value\;
        release(\$ram_lock\);
        \$v5968\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$19235\(31)) & 
                                   eclat_if(work.Int.le(\$12521_loop665_arg\(32 to 47), eclat_resize(\$19235\(0 to 30),16)) & 
                                   work.Int.lt(eclat_resize(\$19235\(0 to 30),16), 
                                               work.Int.add(\$12521_loop665_arg\(32 to 47), X"1770")) & eclat_false) & eclat_false));
        if \$v5968\(0) = '1' then
          \$19239\ := \$19235\ & \$12521_loop665_arg\(16 to 31);
          \$v5951\ := \$ram_lock\;
          if \$v5951\(0) = '1' then
            state := Q_WAIT5950;
          else
            acquire(\$ram_lock\);
            \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(\$12521_loop665_arg\(64 to 79), \$12521_loop665_arg\(0 to 15))));
            \$ram_write\ <= \$19239\(0 to 31); \$ram_write_request\ <= '1';
            state := PAUSE_SET5949;
          end if;
        else
          \$v5967\ := \$ram_lock\;
          if \$v5967\(0) = '1' then
            state := Q_WAIT5966;
          else
            acquire(\$ram_lock\);
            \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19235\(0 to 30),16), X"000" & X"1")));
            state := PAUSE_GET5965;
          end if;
        end if;
      when PAUSE_SET5942 =>
        \$ram_write_request\ <= '0';
        release(\$ram_lock\);
        \$19338\ := eclat_unit;
        \$12520_loop666_arg\ := work.Int.add(\$12520_loop666_arg\(0 to 15), X"000" & X"1") & \$12520_loop666_arg\(16 to 31) & \$12520_loop666_arg\(32 to 47) & \$12520_loop666_arg\(48 to 63);
        state := \$12520_LOOP666\;
      when PAUSE_SET5949 =>
        \$ram_write_request\ <= '0';
        release(\$ram_lock\);
        \$19242\ := eclat_unit;
        \$12521_loop665_arg\ := work.Int.add(\$12521_loop665_arg\(0 to 15), X"000" & X"1") & \$19239\(32 to 47) & \$12521_loop665_arg\(32 to 47) & \$12521_loop665_arg\(48 to 63) & \$12521_loop665_arg\(64 to 79) & \$12521_loop665_arg\(80 to 95);
        state := \$12521_LOOP665\;
      when PAUSE_SET5952 =>
        \$ram_write_request\ <= '0';
        release(\$ram_lock\);
        \$19272\ := eclat_unit;
        \$19239\ := eclat_resize(\$12521_loop665_arg\(16 to 31),31) & eclat_false & 
        work.Int.add(\$12521_loop665_arg\(16 to 31), work.Int.add(eclat_resize(
                                                                  work.Int.lsr(
                                                                  \$19256_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
        \$v5951\ := \$ram_lock\;
        if \$v5951\(0) = '1' then
          state := Q_WAIT5950;
        else
          acquire(\$ram_lock\);
          \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(\$12521_loop665_arg\(64 to 79), \$12521_loop665_arg\(0 to 15))));
          \$ram_write\ <= \$19239\(0 to 31); \$ram_write_request\ <= '1';
          state := PAUSE_SET5949;
        end if;
      when PAUSE_SET5955 =>
        \$ram_write_request\ <= '0';
        release(\$ram_lock\);
        \$19271\ := eclat_unit;
        \$v5954\ := \$ram_lock\;
        if \$v5954\(0) = '1' then
          state := Q_WAIT5953;
        else
          acquire(\$ram_lock\);
          \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19235\(0 to 30),16), X"000" & X"1")));
          \$ram_write\ <= eclat_resize(\$12521_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
          state := PAUSE_SET5952;
        end if;
      when PAUSE_SET5958 =>
        \$ram_write_request\ <= '0';
        release(\$ram_lock\);
        \$19269\ := eclat_unit;
        \$12520_loop666_id\ := "000000000001";
        \$12520_loop666_arg\ := X"000" & X"1" & \$12521_loop665_arg\(16 to 31) & eclat_resize(\$19235\(0 to 30),16) & eclat_resize(
        work.Int.lsr(\$19256_hd\(0 to 30), X"0000000" & X"2"),16);
        state := \$12520_LOOP666\;
      when PAUSE_SET6100 =>
        \$ram_write_request\ <= '0';
        release(\$ram_lock\);
        \$18573\ := eclat_unit;
        \$12523_make_block579_result\ := \$18566\(0 to 31) & \$18566\(32 to 63) & eclat_resize(\$18566\(64 to 79),31) & eclat_false;
        state := \$12523_MAKE_BLOCK579\;
      when Q_WAIT5943 =>
        \$v5944\ := \$ram_lock\;
        if \$v5944\(0) = '1' then
          state := Q_WAIT5943;
        else
          acquire(\$ram_lock\);
          \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(\$12520_loop666_arg\(16 to 31), \$12520_loop666_arg\(0 to 15))));
          \$ram_write\ <= \$19337\; \$ram_write_request\ <= '1';
          state := PAUSE_SET5942;
        end if;
      when Q_WAIT5946 =>
        \$v5947\ := \$ram_lock\;
        if \$v5947\(0) = '1' then
          state := Q_WAIT5946;
        else
          acquire(\$ram_lock\);
          \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$12520_loop666_arg\(32 to 47), \$12520_loop666_arg\(0 to 15))));
          state := PAUSE_GET5945;
        end if;
      when Q_WAIT5950 =>
        \$v5951\ := \$ram_lock\;
        if \$v5951\(0) = '1' then
          state := Q_WAIT5950;
        else
          acquire(\$ram_lock\);
          \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(\$12521_loop665_arg\(64 to 79), \$12521_loop665_arg\(0 to 15))));
          \$ram_write\ <= \$19239\(0 to 31); \$ram_write_request\ <= '1';
          state := PAUSE_SET5949;
        end if;
      when Q_WAIT5953 =>
        \$v5954\ := \$ram_lock\;
        if \$v5954\(0) = '1' then
          state := Q_WAIT5953;
        else
          acquire(\$ram_lock\);
          \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19235\(0 to 30),16), X"000" & X"1")));
          \$ram_write\ <= eclat_resize(\$12521_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
          state := PAUSE_SET5952;
        end if;
      when Q_WAIT5956 =>
        \$v5957\ := \$ram_lock\;
        if \$v5957\(0) = '1' then
          state := Q_WAIT5956;
        else
          acquire(\$ram_lock\);
          \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$19235\(0 to 30),16)));
          \$ram_write\ <= eclat_resize(\$12521_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
          state := PAUSE_SET5955;
        end if;
      when Q_WAIT5959 =>
        \$v5960\ := \$ram_lock\;
        if \$v5960\(0) = '1' then
          state := Q_WAIT5959;
        else
          acquire(\$ram_lock\);
          \$ram_ptr_write\ <= to_integer(unsigned(\$12521_loop665_arg\(16 to 31)));
          \$ram_write\ <= \$19256_hd\; \$ram_write_request\ <= '1';
          state := PAUSE_SET5958;
        end if;
      when Q_WAIT5962 =>
        \$v5963\ := \$ram_lock\;
        if \$v5963\(0) = '1' then
          state := Q_WAIT5962;
        else
          acquire(\$ram_lock\);
          \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$19235\(0 to 30),16)));
          state := PAUSE_GET5961;
        end if;
      when Q_WAIT5966 =>
        \$v5967\ := \$ram_lock\;
        if \$v5967\(0) = '1' then
          state := Q_WAIT5966;
        else
          acquire(\$ram_lock\);
          \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$19235\(0 to 30),16), X"000" & X"1")));
          state := PAUSE_GET5965;
        end if;
      when Q_WAIT5970 =>
        \$v5971\ := \$ram_lock\;
        if \$v5971\(0) = '1' then
          state := Q_WAIT5970;
        else
          acquire(\$ram_lock\);
          \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$12521_loop665_arg\(64 to 79), \$12521_loop665_arg\(0 to 15))));
          state := PAUSE_GET5969;
        end if;
      when Q_WAIT6101 =>
        \$v6102\ := \$ram_lock\;
        if \$v6102\(0) = '1' then
          state := Q_WAIT6101;
        else
          acquire(\$ram_lock\);
          \$ram_ptr_write\ <= to_integer(unsigned(\$18566\(64 to 79)));
          \$ram_write\ <= work.Int.lor(work.Int.lsl(eclat_resize(\$12523_make_block579_arg\(80 to 111),31), X"000000" & X"18"), 
                                       work.Int.lsl(eclat_resize(eclat_if(
                                                                 work.Int.eq(
                                                                 \$12523_make_block579_arg\(112 to 127), X"000" & X"0") & X"000" & X"1" & \$12523_make_block579_arg\(112 to 127)),31), X"0000000" & X"2")) & eclat_true; \$ram_write_request\ <= '1';
          state := PAUSE_SET6100;
        end if;
      when IDLE5941 =>
        rdy5940 := eclat_false;
        \$v7459\ := work.Bool.lnot(""&argument(10));
        if \$v7459\(0) = '1' then
          result5939 := ""&argument(11) & ""&argument(11) & ""&argument(11) & ""&argument(11) & ""&argument(11) & ""&argument(11) & ""&argument(11) & ""&argument(11) & ""&argument(11) & ""&argument(11) & "01100011" & "00000011" & "01110001" & "01110001" & "01100001" & "01100001";
          rdy5940 := eclat_true;
          state := IDLE5941;
        else
          if \$v5866\(0) = '1' then
            
          else
            \$v5866\ := eclat_true;
            \$18553\ := X"0000000" & X"0";
          end if;
          \$18553\ := eclat_if(""&argument(11) & X"0000000" & X"0" & 
                      work.Int.add(\$18553\, X"0000000" & X"1"));
          \$12538_cy\ := \$18553\;
          if \$v5867\(0) = '1' then
            
          else
            \$v5867\ := eclat_true;
            \$12662\ := eclat_false & eclat_false & eclat_false & eclat_false;
          end if;
          \$v7458\ := work.Bool.lnot(""&\$12662\(2));
          if \$v7458\(0) = '1' then
            case state_var7462 is
            when \$12679_LOOP666\ =>
              \$v6121\ := work.Int.ge(\$12679_loop666_arg\(0 to 15), 
                                      work.Int.add(\$12679_loop666_arg\(48 to 63), X"000" & X"1"));
              if \$v6121\(0) = '1' then
                \$12679_loop666_result\ := eclat_unit;
                \$13822\ := \$12679_loop666_result\;
                \$v6130\ := \$ram_lock\;
                if \$v6130\(0) = '1' then
                  state_var7462 := Q_WAIT6129;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$13787\(0 to 30),16)));
                  \$ram_write\ <= eclat_resize(\$12680_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var7462 := PAUSE_SET6128;
                end if;
              else
                \$v6120\ := \$ram_lock\;
                if \$v6120\(0) = '1' then
                  state_var7462 := Q_WAIT6119;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$12679_loop666_arg\(32 to 47), \$12679_loop666_arg\(0 to 15))));
                  state_var7462 := PAUSE_GET6118;
                end if;
              end if;
            when \$12680_LOOP665\ =>
              \$v6145\ := work.Int.ge(\$12680_loop665_arg\(0 to 15), 
                                      work.Int.add(\$12680_loop665_arg\(80 to 95), X"000" & X"1"));
              if \$v6145\(0) = '1' then
                \$12680_loop665_result\ := \$12680_loop665_arg\(16 to 31);
                state_var7462 := \$12680_LOOP665\;
              else
                \$v6144\ := \$ram_lock\;
                if \$v6144\(0) = '1' then
                  state_var7462 := Q_WAIT6143;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$12680_loop665_arg\(64 to 79), \$12680_loop665_arg\(0 to 15))));
                  state_var7462 := PAUSE_GET6142;
                end if;
              end if;
            when \$12681_WAIT662\ =>
              if \$v5869\(0) = '1' then
                
              else
                \$v5869\ := eclat_true;
                \$12792\ := \$12681_wait662_arg\(1 to 32) & \$12681_wait662_arg\(33 to 64) & X"0" & X"fa0" & X"0" & X"fa0" & X"0" & X"fa0" & 
                work.Int.add(X"0" & X"fa0", X"1770") & eclat_false;
              end if;
              case state_var7463 is
              when \$12803_LOOP666\ =>
                \$v6156\ := work.Int.ge(\$12803_loop666_arg\(0 to 15), 
                                        work.Int.add(\$12803_loop666_arg\(48 to 63), X"000" & X"1"));
                if \$v6156\(0) = '1' then
                  \$12803_loop666_result\ := eclat_unit;
                  \$13698\ := \$12803_loop666_result\;
                  \$v6165\ := \$ram_lock\;
                  if \$v6165\(0) = '1' then
                    state_var7463 := Q_WAIT6164;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$13663\(0 to 30),16)));
                    \$ram_write\ <= eclat_resize(\$12804_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var7463 := PAUSE_SET6163;
                  end if;
                else
                  \$v6155\ := \$ram_lock\;
                  if \$v6155\(0) = '1' then
                    state_var7463 := Q_WAIT6154;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$12803_loop666_arg\(32 to 47), \$12803_loop666_arg\(0 to 15))));
                    state_var7463 := PAUSE_GET6153;
                  end if;
                end if;
              when \$12804_LOOP665\ =>
                \$v6180\ := work.Int.ge(\$12804_loop665_arg\(0 to 15), 
                                        work.Int.add(\$12804_loop665_arg\(80 to 95), X"000" & X"1"));
                if \$v6180\(0) = '1' then
                  \$12804_loop665_result\ := \$12804_loop665_arg\(16 to 31);
                  \$13632_next\ := \$12804_loop665_result\;
                  \$12805_aux664_arg\ := work.Int.add(\$12805_aux664_arg\(0 to 15), 
                                                      work.Int.add(eclat_resize(
                                                                   work.Int.lsr(
                                                                   eclat_resize(eclat_resize(\$13628\(0 to 30),16),31), X"0000000" & X"2"),16), X"000" & X"1")) & \$13632_next\ & \$12805_aux664_arg\(32 to 47) & \$12805_aux664_arg\(48 to 63);
                  state_var7463 := \$12805_AUX664\;
                else
                  \$v6179\ := \$ram_lock\;
                  if \$v6179\(0) = '1' then
                    state_var7463 := Q_WAIT6178;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$12804_loop665_arg\(64 to 79), \$12804_loop665_arg\(0 to 15))));
                    state_var7463 := PAUSE_GET6177;
                  end if;
                end if;
              when \$12805_AUX664\ =>
                \$13622\ := work.Print.print_string(clk,of_string("     scan="));
                \$13623\ := work.Int.print(clk,\$12805_aux664_arg\(0 to 15));
                \$13624\ := work.Print.print_string(clk,of_string(" | next="));
                \$13625\ := work.Int.print(clk,\$12805_aux664_arg\(16 to 31));
                \$13626\ := work.Print.print_newline(clk,eclat_unit);
                \$v6184\ := work.Int.ge(\$12805_aux664_arg\(0 to 15), \$12805_aux664_arg\(16 to 31));
                if \$v6184\(0) = '1' then
                  \$12805_aux664_result\ := \$12805_aux664_arg\(16 to 31);
                  state_var7463 := \$12805_AUX664\;
                else
                  \$v6183\ := \$ram_lock\;
                  if \$v6183\(0) = '1' then
                    state_var7463 := Q_WAIT6182;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(\$12805_aux664_arg\(0 to 15)));
                    state_var7463 := PAUSE_GET6181;
                  end if;
                end if;
              when \$12806_LOOP666\ =>
                \$v6191\ := work.Int.ge(\$12806_loop666_arg\(0 to 15), 
                                        work.Int.add(\$12806_loop666_arg\(48 to 63), X"000" & X"1"));
                if \$v6191\(0) = '1' then
                  \$12806_loop666_result\ := eclat_unit;
                  case \$12806_loop666_id\ is
                  when "000000010000" =>
                    \$13538\ := \$12806_loop666_result\;
                    \$v6200\ := \$ram_lock\;
                    if \$v6200\(0) = '1' then
                      state_var7463 := Q_WAIT6199;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$13503\(0 to 30),16)));
                      \$ram_write\ <= eclat_resize(\$12807_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                      state_var7463 := PAUSE_SET6198;
                    end if;
                  when "000000010101" =>
                    \$12943\ := \$12806_loop666_result\;
                    \$v6229\ := \$ram_lock\;
                    if \$v6229\(0) = '1' then
                      state_var7463 := Q_WAIT6228;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$12906\(0 to 30),16)));
                      \$ram_write\ <= eclat_resize(\$12891_copy_root_in_ram6635884_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                      state_var7463 := PAUSE_SET6227;
                    end if;
                  when "000000010111" =>
                    \$13023\ := \$12806_loop666_result\;
                    \$v6253\ := \$ram_lock\;
                    if \$v6253\(0) = '1' then
                      state_var7463 := Q_WAIT6252;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$12879\(0 to 30),16)));
                      \$ram_write\ <= eclat_resize(\$12864_copy_root_in_ram6635886_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                      state_var7463 := PAUSE_SET6251;
                    end if;
                  when "000000011001" =>
                    \$13157\ := \$12806_loop666_result\;
                    \$v6280\ := \$ram_lock\;
                    if \$v6280\(0) = '1' then
                      state_var7463 := Q_WAIT6279;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$13120\(0 to 30),16)));
                      \$ram_write\ <= eclat_resize(\$13105_copy_root_in_ram6635884_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                      state_var7463 := PAUSE_SET6278;
                    end if;
                  when "000000011011" =>
                    \$13237\ := \$12806_loop666_result\;
                    \$v6304\ := \$ram_lock\;
                    if \$v6304\(0) = '1' then
                      state_var7463 := Q_WAIT6303;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$13093\(0 to 30),16)));
                      \$ram_write\ <= eclat_resize(\$13078_copy_root_in_ram6635885_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                      state_var7463 := PAUSE_SET6302;
                    end if;
                  when "000000011101" =>
                    \$13315\ := \$12806_loop666_result\;
                    \$v6325\ := \$ram_lock\;
                    if \$v6325\(0) = '1' then
                      state_var7463 := Q_WAIT6324;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$12681_wait662_arg\(33 to 63),16)));
                      \$ram_write\ <= eclat_resize(\$12818\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                      state_var7463 := PAUSE_SET6323;
                    end if;
                  when "000000011110" =>
                    \$13393\ := \$12806_loop666_result\;
                    \$v6342\ := \$ram_lock\;
                    if \$v6342\(0) = '1' then
                      state_var7463 := Q_WAIT6341;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$12681_wait662_arg\(1 to 31),16)));
                      \$ram_write\ <= eclat_resize(\$12792\(112 to 127),31) & eclat_false; \$ram_write_request\ <= '1';
                      state_var7463 := PAUSE_SET6340;
                    end if;
                  when others =>
                    
                  end case;
                else
                  \$v6190\ := \$ram_lock\;
                  if \$v6190\(0) = '1' then
                    state_var7463 := Q_WAIT6189;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$12806_loop666_arg\(32 to 47), \$12806_loop666_arg\(0 to 15))));
                    state_var7463 := PAUSE_GET6188;
                  end if;
                end if;
              when \$12807_LOOP665\ =>
                \$v6215\ := work.Int.ge(\$12807_loop665_arg\(0 to 15), 
                                        work.Int.add(\$12807_loop665_arg\(80 to 95), X"000" & X"1"));
                if \$v6215\(0) = '1' then
                  \$12807_loop665_result\ := \$12807_loop665_arg\(16 to 31);
                  \$13472_next\ := \$12807_loop665_result\;
                  \$12808_aux664_arg\ := work.Int.add(\$12808_aux664_arg\(0 to 15), 
                                                      work.Int.add(eclat_resize(
                                                                   work.Int.lsr(
                                                                   eclat_resize(eclat_resize(\$13468\(0 to 30),16),31), X"0000000" & X"2"),16), X"000" & X"1")) & \$13472_next\ & \$12808_aux664_arg\(32 to 47) & \$12808_aux664_arg\(48 to 63);
                  state_var7463 := \$12808_AUX664\;
                else
                  \$v6214\ := \$ram_lock\;
                  if \$v6214\(0) = '1' then
                    state_var7463 := Q_WAIT6213;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$12807_loop665_arg\(64 to 79), \$12807_loop665_arg\(0 to 15))));
                    state_var7463 := PAUSE_GET6212;
                  end if;
                end if;
              when \$12808_AUX664\ =>
                \$13462\ := work.Print.print_string(clk,of_string("     scan="));
                \$13463\ := work.Int.print(clk,\$12808_aux664_arg\(0 to 15));
                \$13464\ := work.Print.print_string(clk,of_string(" | next="));
                \$13465\ := work.Int.print(clk,\$12808_aux664_arg\(16 to 31));
                \$13466\ := work.Print.print_newline(clk,eclat_unit);
                \$v6219\ := work.Int.ge(\$12808_aux664_arg\(0 to 15), \$12808_aux664_arg\(16 to 31));
                if \$v6219\(0) = '1' then
                  \$12808_aux664_result\ := \$12808_aux664_arg\(16 to 31);
                  \$12844_next\ := \$12808_aux664_result\;
                  \$12845\ := work.Print.print_string(clk,of_string("memory copied in to_space : "));
                  \$12846\ := work.Int.print(clk,work.Int.sub(\$12844_next\, \$12792\(112 to 127)));
                  \$12847\ := work.Print.print_string(clk,of_string(" words"));
                  \$12848\ := work.Print.print_newline(clk,eclat_unit);
                  \$v6220\ := work.Int.gt(work.Int.sub(\$12844_next\, \$12792\(112 to 127)), X"1770");
                  if \$v6220\(0) = '1' then
                    \$12850\ := work.Print.print_string(clk,of_string("fatal error: "));
                    \$12851\ := work.Print.print_string(clk,of_string("Out of memory"));
                    \$12852\ := work.Print.print_newline(clk,eclat_unit);
                    \$12853_forever6705887_id\ := "000000010011";
                    \$12853_forever6705887_arg\ := eclat_unit;
                    state_var7463 := \$12853_FOREVER6705887\;
                  else
                    \$12824\ := \$12818\(0 to 31) & \$12835\(0 to 31) & \$12844_next\;
                    \$12829\ := work.Print.print_newline(clk,eclat_unit);
                    \$12830\ := work.Print.print_newline(clk,eclat_unit);
                    \$12831\ := work.Print.print_string(clk,of_string("[================= GC END ======================]"));
                    \$12834\ := work.Print.print_newline(clk,eclat_unit);
                    \$12832\ := work.Print.print_newline(clk,eclat_unit);
                    result6147 := \$12824\(0 to 31) & \$12824\(32 to 63) & \$12824\(64 to 79) & 
                    work.Int.add(\$12824\(64 to 79), \$12681_wait662_arg\(81 to 96)) & \$12792\(112 to 127) & \$12792\(96 to 111);
                    rdy6148 := eclat_true;
                    state_var7463 := IDLE6149;
                  end if;
                else
                  \$v6218\ := \$ram_lock\;
                  if \$v6218\(0) = '1' then
                    state_var7463 := Q_WAIT6217;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(\$12808_aux664_arg\(0 to 15)));
                    state_var7463 := PAUSE_GET6216;
                  end if;
                end if;
              when \$12853_FOREVER6705887\ =>
                \$12857_forever6705883_id\ := "000000010010";
                \$12857_forever6705883_arg\ := eclat_unit;
                state_var7463 := \$12857_FOREVER6705883\;
              when \$12857_FOREVER6705883\ =>
                \$12857_forever6705883_arg\ := eclat_unit;
                state_var7463 := \$12857_FOREVER6705883\;
              when \$12864_COPY_ROOT_IN_RAM6635886\ =>
                \$v6268\ := work.Int.ge(\$12864_copy_root_in_ram6635886_arg\(0 to 15), \$12864_copy_root_in_ram6635886_arg\(16 to 31));
                if \$v6268\(0) = '1' then
                  \$12864_copy_root_in_ram6635886_result\ := \$12864_copy_root_in_ram6635886_arg\(32 to 47);
                  \$12840_next\ := \$12864_copy_root_in_ram6635886_result\;
                  \$12842\ := work.Print.print_string(clk,of_string("======================================="));
                  \$12843\ := work.Print.print_newline(clk,eclat_unit);
                  \$12808_aux664_id\ := "000000010100";
                  \$12808_aux664_arg\ := \$12792\(112 to 127) & \$12840_next\ & \$12792\(96 to 111) & \$12792\(112 to 127);
                  state_var7463 := \$12808_AUX664\;
                else
                  \$12876\ := work.Print.print_string(clk,of_string("racine:"));
                  \$12877\ := work.Int.print(clk,\$12864_copy_root_in_ram6635886_arg\(0 to 15));
                  \$12878\ := work.Print.print_newline(clk,eclat_unit);
                  \$v6267\ := \$ram_lock\;
                  if \$v6267\(0) = '1' then
                    state_var7463 := Q_WAIT6266;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(\$12864_copy_root_in_ram6635886_arg\(0 to 15)));
                    state_var7463 := PAUSE_GET6265;
                  end if;
                end if;
              when \$12891_COPY_ROOT_IN_RAM6635884\ =>
                \$v6244\ := work.Int.ge(\$12891_copy_root_in_ram6635884_arg\(0 to 15), \$12891_copy_root_in_ram6635884_arg\(16 to 31));
                if \$v6244\(0) = '1' then
                  \$12891_copy_root_in_ram6635884_result\ := \$12891_copy_root_in_ram6635884_arg\(32 to 47);
                  \$12864_copy_root_in_ram6635886_result\ := \$12891_copy_root_in_ram6635884_result\;
                  \$12840_next\ := \$12864_copy_root_in_ram6635886_result\;
                  \$12842\ := work.Print.print_string(clk,of_string("======================================="));
                  \$12843\ := work.Print.print_newline(clk,eclat_unit);
                  \$12808_aux664_id\ := "000000010100";
                  \$12808_aux664_arg\ := \$12792\(112 to 127) & \$12840_next\ & \$12792\(96 to 111) & \$12792\(112 to 127);
                  state_var7463 := \$12808_AUX664\;
                else
                  \$12903\ := work.Print.print_string(clk,of_string("racine:"));
                  \$12904\ := work.Int.print(clk,\$12891_copy_root_in_ram6635884_arg\(0 to 15));
                  \$12905\ := work.Print.print_newline(clk,eclat_unit);
                  \$v6243\ := \$ram_lock\;
                  if \$v6243\(0) = '1' then
                    state_var7463 := Q_WAIT6242;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(\$12891_copy_root_in_ram6635884_arg\(0 to 15)));
                    state_var7463 := PAUSE_GET6241;
                  end if;
                end if;
              when \$13078_COPY_ROOT_IN_RAM6635885\ =>
                \$v6319\ := work.Int.ge(\$13078_copy_root_in_ram6635885_arg\(0 to 15), \$13078_copy_root_in_ram6635885_arg\(16 to 31));
                if \$v6319\(0) = '1' then
                  \$13078_copy_root_in_ram6635885_result\ := \$13078_copy_root_in_ram6635885_arg\(32 to 47);
                  \$12838_next\ := \$13078_copy_root_in_ram6635885_result\;
                  \$v6271\ := \$global_end_lock\;
                  if \$v6271\(0) = '1' then
                    state_var7463 := Q_WAIT6270;
                  else
                    acquire(\$global_end_lock\);
                    \$global_end_ptr\ <= 0;
                    state_var7463 := PAUSE_GET6269;
                  end if;
                else
                  \$13090\ := work.Print.print_string(clk,of_string("racine:"));
                  \$13091\ := work.Int.print(clk,\$13078_copy_root_in_ram6635885_arg\(0 to 15));
                  \$13092\ := work.Print.print_newline(clk,eclat_unit);
                  \$v6318\ := \$ram_lock\;
                  if \$v6318\(0) = '1' then
                    state_var7463 := Q_WAIT6317;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(\$13078_copy_root_in_ram6635885_arg\(0 to 15)));
                    state_var7463 := PAUSE_GET6316;
                  end if;
                end if;
              when \$13105_COPY_ROOT_IN_RAM6635884\ =>
                \$v6295\ := work.Int.ge(\$13105_copy_root_in_ram6635884_arg\(0 to 15), \$13105_copy_root_in_ram6635884_arg\(16 to 31));
                if \$v6295\(0) = '1' then
                  \$13105_copy_root_in_ram6635884_result\ := \$13105_copy_root_in_ram6635884_arg\(32 to 47);
                  \$13078_copy_root_in_ram6635885_result\ := \$13105_copy_root_in_ram6635884_result\;
                  \$12838_next\ := \$13078_copy_root_in_ram6635885_result\;
                  \$v6271\ := \$global_end_lock\;
                  if \$v6271\(0) = '1' then
                    state_var7463 := Q_WAIT6270;
                  else
                    acquire(\$global_end_lock\);
                    \$global_end_ptr\ <= 0;
                    state_var7463 := PAUSE_GET6269;
                  end if;
                else
                  \$13117\ := work.Print.print_string(clk,of_string("racine:"));
                  \$13118\ := work.Int.print(clk,\$13105_copy_root_in_ram6635884_arg\(0 to 15));
                  \$13119\ := work.Print.print_newline(clk,eclat_unit);
                  \$v6294\ := \$ram_lock\;
                  if \$v6294\(0) = '1' then
                    state_var7463 := Q_WAIT6293;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(\$13105_copy_root_in_ram6635884_arg\(0 to 15)));
                    state_var7463 := PAUSE_GET6292;
                  end if;
                end if;
              when PAUSE_GET6153 =>
                \$13765\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6152\ := \$ram_lock\;
                if \$v6152\(0) = '1' then
                  state_var7463 := Q_WAIT6151;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$12803_loop666_arg\(16 to 31), \$12803_loop666_arg\(0 to 15))));
                  \$ram_write\ <= \$13765\; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6150;
                end if;
              when PAUSE_GET6169 =>
                \$13684_hd\ := \$ram_value\;
                release(\$ram_lock\);
                \$13688\ := work.Print.print_string(clk,of_string("bloc "));
                \$13689\ := work.Int.print(clk,eclat_resize(\$13663\(0 to 30),16));
                \$13690\ := work.Print.print_string(clk,of_string(" of size "));
                \$13691\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                            work.Int.lsr(
                                                            \$13684_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$13692\ := work.Print.print_string(clk,of_string(" from "));
                \$13693\ := work.Int.print(clk,eclat_resize(\$13663\(0 to 30),16));
                \$13694\ := work.Print.print_string(clk,of_string(" to "));
                \$13695\ := work.Int.print(clk,\$12804_loop665_arg\(16 to 31));
                \$13696\ := work.Print.print_newline(clk,eclat_unit);
                \$v6168\ := \$ram_lock\;
                if \$v6168\(0) = '1' then
                  state_var7463 := Q_WAIT6167;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$12804_loop665_arg\(16 to 31)));
                  \$ram_write\ <= \$13684_hd\; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6166;
                end if;
              when PAUSE_GET6173 =>
                \$13679_w\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6172\ := eclat_if(work.Bool.lnot(""&\$13679_w\(31)) & 
                            eclat_if(work.Int.le(\$12804_loop665_arg\(48 to 63), eclat_resize(\$13679_w\(0 to 30),16)) & 
                            work.Int.lt(eclat_resize(\$13679_w\(0 to 30),16), 
                                        work.Int.add(\$12804_loop665_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false);
                if \$v6172\(0) = '1' then
                  \$13667\ := \$13679_w\ & \$12804_loop665_arg\(16 to 31);
                  \$v6159\ := \$ram_lock\;
                  if \$v6159\(0) = '1' then
                    state_var7463 := Q_WAIT6158;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            \$12804_loop665_arg\(64 to 79), \$12804_loop665_arg\(0 to 15))));
                    \$ram_write\ <= \$13667\(0 to 31); \$ram_write_request\ <= '1';
                    state_var7463 := PAUSE_SET6157;
                  end if;
                else
                  \$v6171\ := \$ram_lock\;
                  if \$v6171\(0) = '1' then
                    state_var7463 := Q_WAIT6170;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$13663\(0 to 30),16)));
                    state_var7463 := PAUSE_GET6169;
                  end if;
                end if;
              when PAUSE_GET6177 =>
                \$13663\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6176\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$13663\(31)) & 
                                           eclat_if(work.Int.le(\$12804_loop665_arg\(32 to 47), eclat_resize(\$13663\(0 to 30),16)) & 
                                           work.Int.lt(eclat_resize(\$13663\(0 to 30),16), 
                                                       work.Int.add(\$12804_loop665_arg\(32 to 47), X"1770")) & eclat_false) & eclat_false));
                if \$v6176\(0) = '1' then
                  \$13667\ := \$13663\ & \$12804_loop665_arg\(16 to 31);
                  \$v6159\ := \$ram_lock\;
                  if \$v6159\(0) = '1' then
                    state_var7463 := Q_WAIT6158;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            \$12804_loop665_arg\(64 to 79), \$12804_loop665_arg\(0 to 15))));
                    \$ram_write\ <= \$13667\(0 to 31); \$ram_write_request\ <= '1';
                    state_var7463 := PAUSE_SET6157;
                  end if;
                else
                  \$v6175\ := \$ram_lock\;
                  if \$v6175\(0) = '1' then
                    state_var7463 := Q_WAIT6174;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$13663\(0 to 30),16), X"000" & X"1")));
                    state_var7463 := PAUSE_GET6173;
                  end if;
                end if;
              when PAUSE_GET6181 =>
                \$13628\ := \$ram_value\;
                release(\$ram_lock\);
                \$12804_loop665_id\ := "000000001111";
                \$12804_loop665_arg\ := X"000" & X"1" & \$12805_aux664_arg\(16 to 31) & \$12805_aux664_arg\(32 to 47) & \$12805_aux664_arg\(48 to 63) & \$12805_aux664_arg\(0 to 15) & eclat_resize(
                work.Int.lsr(eclat_resize(eclat_resize(\$13628\(0 to 30),16),31), X"0000000" & X"2"),16);
                state_var7463 := \$12804_LOOP665\;
              when PAUSE_GET6188 =>
                \$13605\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6187\ := \$ram_lock\;
                if \$v6187\(0) = '1' then
                  state_var7463 := Q_WAIT6186;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$12806_loop666_arg\(16 to 31), \$12806_loop666_arg\(0 to 15))));
                  \$ram_write\ <= \$13605\; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6185;
                end if;
              when PAUSE_GET6204 =>
                \$13524_hd\ := \$ram_value\;
                release(\$ram_lock\);
                \$13528\ := work.Print.print_string(clk,of_string("bloc "));
                \$13529\ := work.Int.print(clk,eclat_resize(\$13503\(0 to 30),16));
                \$13530\ := work.Print.print_string(clk,of_string(" of size "));
                \$13531\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                            work.Int.lsr(
                                                            \$13524_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$13532\ := work.Print.print_string(clk,of_string(" from "));
                \$13533\ := work.Int.print(clk,eclat_resize(\$13503\(0 to 30),16));
                \$13534\ := work.Print.print_string(clk,of_string(" to "));
                \$13535\ := work.Int.print(clk,\$12807_loop665_arg\(16 to 31));
                \$13536\ := work.Print.print_newline(clk,eclat_unit);
                \$v6203\ := \$ram_lock\;
                if \$v6203\(0) = '1' then
                  state_var7463 := Q_WAIT6202;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$12807_loop665_arg\(16 to 31)));
                  \$ram_write\ <= \$13524_hd\; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6201;
                end if;
              when PAUSE_GET6208 =>
                \$13519_w\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6207\ := eclat_if(work.Bool.lnot(""&\$13519_w\(31)) & 
                            eclat_if(work.Int.le(\$12807_loop665_arg\(48 to 63), eclat_resize(\$13519_w\(0 to 30),16)) & 
                            work.Int.lt(eclat_resize(\$13519_w\(0 to 30),16), 
                                        work.Int.add(\$12807_loop665_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false);
                if \$v6207\(0) = '1' then
                  \$13507\ := \$13519_w\ & \$12807_loop665_arg\(16 to 31);
                  \$v6194\ := \$ram_lock\;
                  if \$v6194\(0) = '1' then
                    state_var7463 := Q_WAIT6193;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            \$12807_loop665_arg\(64 to 79), \$12807_loop665_arg\(0 to 15))));
                    \$ram_write\ <= \$13507\(0 to 31); \$ram_write_request\ <= '1';
                    state_var7463 := PAUSE_SET6192;
                  end if;
                else
                  \$v6206\ := \$ram_lock\;
                  if \$v6206\(0) = '1' then
                    state_var7463 := Q_WAIT6205;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$13503\(0 to 30),16)));
                    state_var7463 := PAUSE_GET6204;
                  end if;
                end if;
              when PAUSE_GET6212 =>
                \$13503\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6211\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$13503\(31)) & 
                                           eclat_if(work.Int.le(\$12807_loop665_arg\(32 to 47), eclat_resize(\$13503\(0 to 30),16)) & 
                                           work.Int.lt(eclat_resize(\$13503\(0 to 30),16), 
                                                       work.Int.add(\$12807_loop665_arg\(32 to 47), X"1770")) & eclat_false) & eclat_false));
                if \$v6211\(0) = '1' then
                  \$13507\ := \$13503\ & \$12807_loop665_arg\(16 to 31);
                  \$v6194\ := \$ram_lock\;
                  if \$v6194\(0) = '1' then
                    state_var7463 := Q_WAIT6193;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            \$12807_loop665_arg\(64 to 79), \$12807_loop665_arg\(0 to 15))));
                    \$ram_write\ <= \$13507\(0 to 31); \$ram_write_request\ <= '1';
                    state_var7463 := PAUSE_SET6192;
                  end if;
                else
                  \$v6210\ := \$ram_lock\;
                  if \$v6210\(0) = '1' then
                    state_var7463 := Q_WAIT6209;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$13503\(0 to 30),16), X"000" & X"1")));
                    state_var7463 := PAUSE_GET6208;
                  end if;
                end if;
              when PAUSE_GET6216 =>
                \$13468\ := \$ram_value\;
                release(\$ram_lock\);
                \$12807_loop665_id\ := "000000010001";
                \$12807_loop665_arg\ := X"000" & X"1" & \$12808_aux664_arg\(16 to 31) & \$12808_aux664_arg\(32 to 47) & \$12808_aux664_arg\(48 to 63) & \$12808_aux664_arg\(0 to 15) & eclat_resize(
                work.Int.lsr(eclat_resize(eclat_resize(\$13468\(0 to 30),16),31), X"0000000" & X"2"),16);
                state_var7463 := \$12807_LOOP665\;
              when PAUSE_GET6233 =>
                \$12929_hd\ := \$ram_value\;
                release(\$ram_lock\);
                \$12933\ := work.Print.print_string(clk,of_string("bloc "));
                \$12934\ := work.Int.print(clk,eclat_resize(\$12906\(0 to 30),16));
                \$12935\ := work.Print.print_string(clk,of_string(" of size "));
                \$12936\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                            work.Int.lsr(
                                                            \$12929_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$12937\ := work.Print.print_string(clk,of_string(" from "));
                \$12938\ := work.Int.print(clk,eclat_resize(\$12906\(0 to 30),16));
                \$12939\ := work.Print.print_string(clk,of_string(" to "));
                \$12940\ := work.Int.print(clk,\$12891_copy_root_in_ram6635884_arg\(32 to 47));
                \$12941\ := work.Print.print_newline(clk,eclat_unit);
                \$v6232\ := \$ram_lock\;
                if \$v6232\(0) = '1' then
                  state_var7463 := Q_WAIT6231;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$12891_copy_root_in_ram6635884_arg\(32 to 47)));
                  \$ram_write\ <= \$12929_hd\; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6230;
                end if;
              when PAUSE_GET6237 =>
                \$12924_w\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6236\ := eclat_if(work.Bool.lnot(""&\$12924_w\(31)) & 
                            eclat_if(work.Int.le(\$12891_copy_root_in_ram6635884_arg\(64 to 79), eclat_resize(\$12924_w\(0 to 30),16)) & 
                            work.Int.lt(eclat_resize(\$12924_w\(0 to 30),16), 
                                        work.Int.add(\$12891_copy_root_in_ram6635884_arg\(64 to 79), X"1770")) & eclat_false) & eclat_false);
                if \$v6236\(0) = '1' then
                  \$12910\ := \$12924_w\ & \$12891_copy_root_in_ram6635884_arg\(32 to 47);
                  \$v6223\ := \$ram_lock\;
                  if \$v6223\(0) = '1' then
                    state_var7463 := Q_WAIT6222;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$12891_copy_root_in_ram6635884_arg\(0 to 15)));
                    \$ram_write\ <= \$12910\(0 to 31); \$ram_write_request\ <= '1';
                    state_var7463 := PAUSE_SET6221;
                  end if;
                else
                  \$v6235\ := \$ram_lock\;
                  if \$v6235\(0) = '1' then
                    state_var7463 := Q_WAIT6234;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$12906\(0 to 30),16)));
                    state_var7463 := PAUSE_GET6233;
                  end if;
                end if;
              when PAUSE_GET6241 =>
                \$12906\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6240\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$12906\(31)) & 
                                           eclat_if(work.Int.le(\$12891_copy_root_in_ram6635884_arg\(48 to 63), eclat_resize(\$12906\(0 to 30),16)) & 
                                           work.Int.lt(eclat_resize(\$12906\(0 to 30),16), 
                                                       work.Int.add(\$12891_copy_root_in_ram6635884_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false));
                if \$v6240\(0) = '1' then
                  \$12910\ := \$12906\ & \$12891_copy_root_in_ram6635884_arg\(32 to 47);
                  \$v6223\ := \$ram_lock\;
                  if \$v6223\(0) = '1' then
                    state_var7463 := Q_WAIT6222;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$12891_copy_root_in_ram6635884_arg\(0 to 15)));
                    \$ram_write\ <= \$12910\(0 to 31); \$ram_write_request\ <= '1';
                    state_var7463 := PAUSE_SET6221;
                  end if;
                else
                  \$v6239\ := \$ram_lock\;
                  if \$v6239\(0) = '1' then
                    state_var7463 := Q_WAIT6238;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$12906\(0 to 30),16), X"000" & X"1")));
                    state_var7463 := PAUSE_GET6237;
                  end if;
                end if;
              when PAUSE_GET6257 =>
                \$13009_hd\ := \$ram_value\;
                release(\$ram_lock\);
                \$13013\ := work.Print.print_string(clk,of_string("bloc "));
                \$13014\ := work.Int.print(clk,eclat_resize(\$12879\(0 to 30),16));
                \$13015\ := work.Print.print_string(clk,of_string(" of size "));
                \$13016\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                            work.Int.lsr(
                                                            \$13009_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$13017\ := work.Print.print_string(clk,of_string(" from "));
                \$13018\ := work.Int.print(clk,eclat_resize(\$12879\(0 to 30),16));
                \$13019\ := work.Print.print_string(clk,of_string(" to "));
                \$13020\ := work.Int.print(clk,\$12864_copy_root_in_ram6635886_arg\(32 to 47));
                \$13021\ := work.Print.print_newline(clk,eclat_unit);
                \$v6256\ := \$ram_lock\;
                if \$v6256\(0) = '1' then
                  state_var7463 := Q_WAIT6255;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$12864_copy_root_in_ram6635886_arg\(32 to 47)));
                  \$ram_write\ <= \$13009_hd\; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6254;
                end if;
              when PAUSE_GET6261 =>
                \$13004_w\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6260\ := eclat_if(work.Bool.lnot(""&\$13004_w\(31)) & 
                            eclat_if(work.Int.le(\$12864_copy_root_in_ram6635886_arg\(64 to 79), eclat_resize(\$13004_w\(0 to 30),16)) & 
                            work.Int.lt(eclat_resize(\$13004_w\(0 to 30),16), 
                                        work.Int.add(\$12864_copy_root_in_ram6635886_arg\(64 to 79), X"1770")) & eclat_false) & eclat_false);
                if \$v6260\(0) = '1' then
                  \$12883\ := \$13004_w\ & \$12864_copy_root_in_ram6635886_arg\(32 to 47);
                  \$v6247\ := \$ram_lock\;
                  if \$v6247\(0) = '1' then
                    state_var7463 := Q_WAIT6246;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$12864_copy_root_in_ram6635886_arg\(0 to 15)));
                    \$ram_write\ <= \$12883\(0 to 31); \$ram_write_request\ <= '1';
                    state_var7463 := PAUSE_SET6245;
                  end if;
                else
                  \$v6259\ := \$ram_lock\;
                  if \$v6259\(0) = '1' then
                    state_var7463 := Q_WAIT6258;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$12879\(0 to 30),16)));
                    state_var7463 := PAUSE_GET6257;
                  end if;
                end if;
              when PAUSE_GET6265 =>
                \$12879\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6264\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$12879\(31)) & 
                                           eclat_if(work.Int.le(\$12864_copy_root_in_ram6635886_arg\(48 to 63), eclat_resize(\$12879\(0 to 30),16)) & 
                                           work.Int.lt(eclat_resize(\$12879\(0 to 30),16), 
                                                       work.Int.add(\$12864_copy_root_in_ram6635886_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false));
                if \$v6264\(0) = '1' then
                  \$12883\ := \$12879\ & \$12864_copy_root_in_ram6635886_arg\(32 to 47);
                  \$v6247\ := \$ram_lock\;
                  if \$v6247\(0) = '1' then
                    state_var7463 := Q_WAIT6246;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$12864_copy_root_in_ram6635886_arg\(0 to 15)));
                    \$ram_write\ <= \$12883\(0 to 31); \$ram_write_request\ <= '1';
                    state_var7463 := PAUSE_SET6245;
                  end if;
                else
                  \$v6263\ := \$ram_lock\;
                  if \$v6263\(0) = '1' then
                    state_var7463 := Q_WAIT6262;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$12879\(0 to 30),16), X"000" & X"1")));
                    state_var7463 := PAUSE_GET6261;
                  end if;
                end if;
              when PAUSE_GET6269 =>
                \$12839\ := \$global_end_value\;
                release(\$global_end_lock\);
                \$12864_copy_root_in_ram6635886_id\ := "000000011000";
                \$12864_copy_root_in_ram6635886_arg\ := X"3e80" & \$12839\ & \$12838_next\ & \$12792\(96 to 111) & \$12792\(112 to 127);
                state_var7463 := \$12864_COPY_ROOT_IN_RAM6635886\;
              when PAUSE_GET6284 =>
                \$13143_hd\ := \$ram_value\;
                release(\$ram_lock\);
                \$13147\ := work.Print.print_string(clk,of_string("bloc "));
                \$13148\ := work.Int.print(clk,eclat_resize(\$13120\(0 to 30),16));
                \$13149\ := work.Print.print_string(clk,of_string(" of size "));
                \$13150\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                            work.Int.lsr(
                                                            \$13143_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$13151\ := work.Print.print_string(clk,of_string(" from "));
                \$13152\ := work.Int.print(clk,eclat_resize(\$13120\(0 to 30),16));
                \$13153\ := work.Print.print_string(clk,of_string(" to "));
                \$13154\ := work.Int.print(clk,\$13105_copy_root_in_ram6635884_arg\(32 to 47));
                \$13155\ := work.Print.print_newline(clk,eclat_unit);
                \$v6283\ := \$ram_lock\;
                if \$v6283\(0) = '1' then
                  state_var7463 := Q_WAIT6282;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13105_copy_root_in_ram6635884_arg\(32 to 47)));
                  \$ram_write\ <= \$13143_hd\; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6281;
                end if;
              when PAUSE_GET6288 =>
                \$13138_w\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6287\ := eclat_if(work.Bool.lnot(""&\$13138_w\(31)) & 
                            eclat_if(work.Int.le(\$13105_copy_root_in_ram6635884_arg\(64 to 79), eclat_resize(\$13138_w\(0 to 30),16)) & 
                            work.Int.lt(eclat_resize(\$13138_w\(0 to 30),16), 
                                        work.Int.add(\$13105_copy_root_in_ram6635884_arg\(64 to 79), X"1770")) & eclat_false) & eclat_false);
                if \$v6287\(0) = '1' then
                  \$13124\ := \$13138_w\ & \$13105_copy_root_in_ram6635884_arg\(32 to 47);
                  \$v6274\ := \$ram_lock\;
                  if \$v6274\(0) = '1' then
                    state_var7463 := Q_WAIT6273;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13105_copy_root_in_ram6635884_arg\(0 to 15)));
                    \$ram_write\ <= \$13124\(0 to 31); \$ram_write_request\ <= '1';
                    state_var7463 := PAUSE_SET6272;
                  end if;
                else
                  \$v6286\ := \$ram_lock\;
                  if \$v6286\(0) = '1' then
                    state_var7463 := Q_WAIT6285;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$13120\(0 to 30),16)));
                    state_var7463 := PAUSE_GET6284;
                  end if;
                end if;
              when PAUSE_GET6292 =>
                \$13120\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6291\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$13120\(31)) & 
                                           eclat_if(work.Int.le(\$13105_copy_root_in_ram6635884_arg\(48 to 63), eclat_resize(\$13120\(0 to 30),16)) & 
                                           work.Int.lt(eclat_resize(\$13120\(0 to 30),16), 
                                                       work.Int.add(\$13105_copy_root_in_ram6635884_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false));
                if \$v6291\(0) = '1' then
                  \$13124\ := \$13120\ & \$13105_copy_root_in_ram6635884_arg\(32 to 47);
                  \$v6274\ := \$ram_lock\;
                  if \$v6274\(0) = '1' then
                    state_var7463 := Q_WAIT6273;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13105_copy_root_in_ram6635884_arg\(0 to 15)));
                    \$ram_write\ <= \$13124\(0 to 31); \$ram_write_request\ <= '1';
                    state_var7463 := PAUSE_SET6272;
                  end if;
                else
                  \$v6290\ := \$ram_lock\;
                  if \$v6290\(0) = '1' then
                    state_var7463 := Q_WAIT6289;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$13120\(0 to 30),16), X"000" & X"1")));
                    state_var7463 := PAUSE_GET6288;
                  end if;
                end if;
              when PAUSE_GET6308 =>
                \$13223_hd\ := \$ram_value\;
                release(\$ram_lock\);
                \$13227\ := work.Print.print_string(clk,of_string("bloc "));
                \$13228\ := work.Int.print(clk,eclat_resize(\$13093\(0 to 30),16));
                \$13229\ := work.Print.print_string(clk,of_string(" of size "));
                \$13230\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                            work.Int.lsr(
                                                            \$13223_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$13231\ := work.Print.print_string(clk,of_string(" from "));
                \$13232\ := work.Int.print(clk,eclat_resize(\$13093\(0 to 30),16));
                \$13233\ := work.Print.print_string(clk,of_string(" to "));
                \$13234\ := work.Int.print(clk,\$13078_copy_root_in_ram6635885_arg\(32 to 47));
                \$13235\ := work.Print.print_newline(clk,eclat_unit);
                \$v6307\ := \$ram_lock\;
                if \$v6307\(0) = '1' then
                  state_var7463 := Q_WAIT6306;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13078_copy_root_in_ram6635885_arg\(32 to 47)));
                  \$ram_write\ <= \$13223_hd\; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6305;
                end if;
              when PAUSE_GET6312 =>
                \$13218_w\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6311\ := eclat_if(work.Bool.lnot(""&\$13218_w\(31)) & 
                            eclat_if(work.Int.le(\$13078_copy_root_in_ram6635885_arg\(64 to 79), eclat_resize(\$13218_w\(0 to 30),16)) & 
                            work.Int.lt(eclat_resize(\$13218_w\(0 to 30),16), 
                                        work.Int.add(\$13078_copy_root_in_ram6635885_arg\(64 to 79), X"1770")) & eclat_false) & eclat_false);
                if \$v6311\(0) = '1' then
                  \$13097\ := \$13218_w\ & \$13078_copy_root_in_ram6635885_arg\(32 to 47);
                  \$v6298\ := \$ram_lock\;
                  if \$v6298\(0) = '1' then
                    state_var7463 := Q_WAIT6297;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13078_copy_root_in_ram6635885_arg\(0 to 15)));
                    \$ram_write\ <= \$13097\(0 to 31); \$ram_write_request\ <= '1';
                    state_var7463 := PAUSE_SET6296;
                  end if;
                else
                  \$v6310\ := \$ram_lock\;
                  if \$v6310\(0) = '1' then
                    state_var7463 := Q_WAIT6309;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$13093\(0 to 30),16)));
                    state_var7463 := PAUSE_GET6308;
                  end if;
                end if;
              when PAUSE_GET6316 =>
                \$13093\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6315\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$13093\(31)) & 
                                           eclat_if(work.Int.le(\$13078_copy_root_in_ram6635885_arg\(48 to 63), eclat_resize(\$13093\(0 to 30),16)) & 
                                           work.Int.lt(eclat_resize(\$13093\(0 to 30),16), 
                                                       work.Int.add(\$13078_copy_root_in_ram6635885_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false));
                if \$v6315\(0) = '1' then
                  \$13097\ := \$13093\ & \$13078_copy_root_in_ram6635885_arg\(32 to 47);
                  \$v6298\ := \$ram_lock\;
                  if \$v6298\(0) = '1' then
                    state_var7463 := Q_WAIT6297;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13078_copy_root_in_ram6635885_arg\(0 to 15)));
                    \$ram_write\ <= \$13097\(0 to 31); \$ram_write_request\ <= '1';
                    state_var7463 := PAUSE_SET6296;
                  end if;
                else
                  \$v6314\ := \$ram_lock\;
                  if \$v6314\(0) = '1' then
                    state_var7463 := Q_WAIT6313;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$13093\(0 to 30),16), X"000" & X"1")));
                    state_var7463 := PAUSE_GET6312;
                  end if;
                end if;
              when PAUSE_GET6329 =>
                \$13301_hd\ := \$ram_value\;
                release(\$ram_lock\);
                \$13305\ := work.Print.print_string(clk,of_string("bloc "));
                \$13306\ := work.Int.print(clk,eclat_resize(\$12681_wait662_arg\(33 to 63),16));
                \$13307\ := work.Print.print_string(clk,of_string(" of size "));
                \$13308\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                            work.Int.lsr(
                                                            \$13301_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$13309\ := work.Print.print_string(clk,of_string(" from "));
                \$13310\ := work.Int.print(clk,eclat_resize(\$12681_wait662_arg\(33 to 63),16));
                \$13311\ := work.Print.print_string(clk,of_string(" to "));
                \$13312\ := work.Int.print(clk,\$12818\(32 to 47));
                \$13313\ := work.Print.print_newline(clk,eclat_unit);
                \$v6328\ := \$ram_lock\;
                if \$v6328\(0) = '1' then
                  state_var7463 := Q_WAIT6327;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$12818\(32 to 47)));
                  \$ram_write\ <= \$13301_hd\; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6326;
                end if;
              when PAUSE_GET6333 =>
                \$13296_w\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6332\ := eclat_if(work.Bool.lnot(""&\$13296_w\(31)) & 
                            eclat_if(work.Int.le(\$12792\(112 to 127), eclat_resize(\$13296_w\(0 to 30),16)) & 
                            work.Int.lt(eclat_resize(\$13296_w\(0 to 30),16), 
                                        work.Int.add(\$12792\(112 to 127), X"1770")) & eclat_false) & eclat_false);
                if \$v6332\(0) = '1' then
                  \$12835\ := \$13296_w\ & \$12818\(32 to 47);
                  \$13078_copy_root_in_ram6635885_id\ := "000000011100";
                  \$13078_copy_root_in_ram6635885_arg\ := X"0" & X"3e8" & \$12681_wait662_arg\(65 to 80) & \$12835\(32 to 47) & \$12792\(96 to 111) & \$12792\(112 to 127);
                  state_var7463 := \$13078_COPY_ROOT_IN_RAM6635885\;
                else
                  \$v6331\ := \$ram_lock\;
                  if \$v6331\(0) = '1' then
                    state_var7463 := Q_WAIT6330;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$12681_wait662_arg\(33 to 63),16)));
                    state_var7463 := PAUSE_GET6329;
                  end if;
                end if;
              when PAUSE_GET6346 =>
                \$13379_hd\ := \$ram_value\;
                release(\$ram_lock\);
                \$13383\ := work.Print.print_string(clk,of_string("bloc "));
                \$13384\ := work.Int.print(clk,eclat_resize(\$12681_wait662_arg\(1 to 31),16));
                \$13385\ := work.Print.print_string(clk,of_string(" of size "));
                \$13386\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                            work.Int.lsr(
                                                            \$13379_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$13387\ := work.Print.print_string(clk,of_string(" from "));
                \$13388\ := work.Int.print(clk,eclat_resize(\$12681_wait662_arg\(1 to 31),16));
                \$13389\ := work.Print.print_string(clk,of_string(" to "));
                \$13390\ := work.Int.print(clk,\$12792\(112 to 127));
                \$13391\ := work.Print.print_newline(clk,eclat_unit);
                \$v6345\ := \$ram_lock\;
                if \$v6345\(0) = '1' then
                  state_var7463 := Q_WAIT6344;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$12792\(112 to 127)));
                  \$ram_write\ <= \$13379_hd\; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6343;
                end if;
              when PAUSE_GET6350 =>
                \$13374_w\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6349\ := eclat_if(work.Bool.lnot(""&\$13374_w\(31)) & 
                            eclat_if(work.Int.le(\$12792\(112 to 127), eclat_resize(\$13374_w\(0 to 30),16)) & 
                            work.Int.lt(eclat_resize(\$13374_w\(0 to 30),16), 
                                        work.Int.add(\$12792\(112 to 127), X"1770")) & eclat_false) & eclat_false);
                if \$v6349\(0) = '1' then
                  \$12818\ := \$13374_w\ & \$12792\(112 to 127);
                  \$v6336\ := work.Bool.lnot(eclat_if(work.Bool.lnot(
                                                      ""&\$12681_wait662_arg\(64)) & 
                                             eclat_if(work.Int.le(\$12792\(96 to 111), eclat_resize(\$12681_wait662_arg\(33 to 63),16)) & 
                                             work.Int.lt(eclat_resize(\$12681_wait662_arg\(33 to 63),16), 
                                                         work.Int.add(
                                                         \$12792\(96 to 111), X"1770")) & eclat_false) & eclat_false));
                  if \$v6336\(0) = '1' then
                    \$12835\ := \$12681_wait662_arg\(33 to 64) & \$12818\(32 to 47);
                    \$13078_copy_root_in_ram6635885_id\ := "000000011100";
                    \$13078_copy_root_in_ram6635885_arg\ := X"0" & X"3e8" & \$12681_wait662_arg\(65 to 80) & \$12835\(32 to 47) & \$12792\(96 to 111) & \$12792\(112 to 127);
                    state_var7463 := \$13078_COPY_ROOT_IN_RAM6635885\;
                  else
                    \$v6335\ := \$ram_lock\;
                    if \$v6335\(0) = '1' then
                      state_var7463 := Q_WAIT6334;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                        eclat_resize(\$12681_wait662_arg\(33 to 63),16), X"000" & X"1")));
                      state_var7463 := PAUSE_GET6333;
                    end if;
                  end if;
                else
                  \$v6348\ := \$ram_lock\;
                  if \$v6348\(0) = '1' then
                    state_var7463 := Q_WAIT6347;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$12681_wait662_arg\(1 to 31),16)));
                    state_var7463 := PAUSE_GET6346;
                  end if;
                end if;
              when PAUSE_SET6150 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$13766\ := eclat_unit;
                \$12803_loop666_arg\ := work.Int.add(\$12803_loop666_arg\(0 to 15), X"000" & X"1") & \$12803_loop666_arg\(16 to 31) & \$12803_loop666_arg\(32 to 47) & \$12803_loop666_arg\(48 to 63);
                state_var7463 := \$12803_LOOP666\;
              when PAUSE_SET6157 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$13670\ := eclat_unit;
                \$12804_loop665_arg\ := work.Int.add(\$12804_loop665_arg\(0 to 15), X"000" & X"1") & \$13667\(32 to 47) & \$12804_loop665_arg\(32 to 47) & \$12804_loop665_arg\(48 to 63) & \$12804_loop665_arg\(64 to 79) & \$12804_loop665_arg\(80 to 95);
                state_var7463 := \$12804_LOOP665\;
              when PAUSE_SET6160 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$13700\ := eclat_unit;
                \$13667\ := eclat_resize(\$12804_loop665_arg\(16 to 31),31) & eclat_false & 
                work.Int.add(\$12804_loop665_arg\(16 to 31), work.Int.add(
                                                             eclat_resize(
                                                             work.Int.lsr(
                                                             \$13684_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$v6159\ := \$ram_lock\;
                if \$v6159\(0) = '1' then
                  state_var7463 := Q_WAIT6158;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$12804_loop665_arg\(64 to 79), \$12804_loop665_arg\(0 to 15))));
                  \$ram_write\ <= \$13667\(0 to 31); \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6157;
                end if;
              when PAUSE_SET6163 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$13699\ := eclat_unit;
                \$v6162\ := \$ram_lock\;
                if \$v6162\(0) = '1' then
                  state_var7463 := Q_WAIT6161;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$13663\(0 to 30),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$12804_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6160;
                end if;
              when PAUSE_SET6166 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$13697\ := eclat_unit;
                \$12803_loop666_id\ := "000000001110";
                \$12803_loop666_arg\ := X"000" & X"1" & \$12804_loop665_arg\(16 to 31) & eclat_resize(\$13663\(0 to 30),16) & eclat_resize(
                work.Int.lsr(\$13684_hd\(0 to 30), X"0000000" & X"2"),16);
                state_var7463 := \$12803_LOOP666\;
              when PAUSE_SET6185 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$13606\ := eclat_unit;
                \$12806_loop666_arg\ := work.Int.add(\$12806_loop666_arg\(0 to 15), X"000" & X"1") & \$12806_loop666_arg\(16 to 31) & \$12806_loop666_arg\(32 to 47) & \$12806_loop666_arg\(48 to 63);
                state_var7463 := \$12806_LOOP666\;
              when PAUSE_SET6192 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$13510\ := eclat_unit;
                \$12807_loop665_arg\ := work.Int.add(\$12807_loop665_arg\(0 to 15), X"000" & X"1") & \$13507\(32 to 47) & \$12807_loop665_arg\(32 to 47) & \$12807_loop665_arg\(48 to 63) & \$12807_loop665_arg\(64 to 79) & \$12807_loop665_arg\(80 to 95);
                state_var7463 := \$12807_LOOP665\;
              when PAUSE_SET6195 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$13540\ := eclat_unit;
                \$13507\ := eclat_resize(\$12807_loop665_arg\(16 to 31),31) & eclat_false & 
                work.Int.add(\$12807_loop665_arg\(16 to 31), work.Int.add(
                                                             eclat_resize(
                                                             work.Int.lsr(
                                                             \$13524_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$v6194\ := \$ram_lock\;
                if \$v6194\(0) = '1' then
                  state_var7463 := Q_WAIT6193;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$12807_loop665_arg\(64 to 79), \$12807_loop665_arg\(0 to 15))));
                  \$ram_write\ <= \$13507\(0 to 31); \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6192;
                end if;
              when PAUSE_SET6198 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$13539\ := eclat_unit;
                \$v6197\ := \$ram_lock\;
                if \$v6197\(0) = '1' then
                  state_var7463 := Q_WAIT6196;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$13503\(0 to 30),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$12807_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6195;
                end if;
              when PAUSE_SET6201 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$13537\ := eclat_unit;
                \$12806_loop666_id\ := "000000010000";
                \$12806_loop666_arg\ := X"000" & X"1" & \$12807_loop665_arg\(16 to 31) & eclat_resize(\$13503\(0 to 30),16) & eclat_resize(
                work.Int.lsr(\$13524_hd\(0 to 30), X"0000000" & X"2"),16);
                state_var7463 := \$12806_LOOP666\;
              when PAUSE_SET6221 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$12913\ := eclat_unit;
                \$12914\ := work.Print.print_string(clk,of_string(" next="));
                \$12915\ := work.Int.print(clk,\$12910\(32 to 47));
                \$12916\ := work.Print.print_newline(clk,eclat_unit);
                \$12891_copy_root_in_ram6635884_arg\ := work.Int.add(
                                                        \$12891_copy_root_in_ram6635884_arg\(0 to 15), X"000" & X"1") & \$12891_copy_root_in_ram6635884_arg\(16 to 31) & \$12910\(32 to 47) & \$12891_copy_root_in_ram6635884_arg\(48 to 63) & \$12891_copy_root_in_ram6635884_arg\(64 to 79);
                state_var7463 := \$12891_COPY_ROOT_IN_RAM6635884\;
              when PAUSE_SET6224 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$12945\ := eclat_unit;
                \$12910\ := eclat_resize(\$12891_copy_root_in_ram6635884_arg\(32 to 47),31) & eclat_false & 
                work.Int.add(\$12891_copy_root_in_ram6635884_arg\(32 to 47), 
                             work.Int.add(eclat_resize(work.Int.lsr(\$12929_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$v6223\ := \$ram_lock\;
                if \$v6223\(0) = '1' then
                  state_var7463 := Q_WAIT6222;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$12891_copy_root_in_ram6635884_arg\(0 to 15)));
                  \$ram_write\ <= \$12910\(0 to 31); \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6221;
                end if;
              when PAUSE_SET6227 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$12944\ := eclat_unit;
                \$v6226\ := \$ram_lock\;
                if \$v6226\(0) = '1' then
                  state_var7463 := Q_WAIT6225;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$12906\(0 to 30),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$12891_copy_root_in_ram6635884_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6224;
                end if;
              when PAUSE_SET6230 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$12942\ := eclat_unit;
                \$12806_loop666_id\ := "000000010101";
                \$12806_loop666_arg\ := X"000" & X"1" & \$12891_copy_root_in_ram6635884_arg\(32 to 47) & eclat_resize(\$12906\(0 to 30),16) & eclat_resize(
                work.Int.lsr(\$12929_hd\(0 to 30), X"0000000" & X"2"),16);
                state_var7463 := \$12806_LOOP666\;
              when PAUSE_SET6245 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$12886\ := eclat_unit;
                \$12887\ := work.Print.print_string(clk,of_string(" next="));
                \$12888\ := work.Int.print(clk,\$12883\(32 to 47));
                \$12889\ := work.Print.print_newline(clk,eclat_unit);
                \$12891_copy_root_in_ram6635884_id\ := "000000010110";
                \$12891_copy_root_in_ram6635884_arg\ := work.Int.add(
                                                        \$12864_copy_root_in_ram6635886_arg\(0 to 15), X"000" & X"1") & \$12864_copy_root_in_ram6635886_arg\(16 to 31) & \$12883\(32 to 47) & \$12864_copy_root_in_ram6635886_arg\(48 to 63) & \$12864_copy_root_in_ram6635886_arg\(64 to 79);
                state_var7463 := \$12891_COPY_ROOT_IN_RAM6635884\;
              when PAUSE_SET6248 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$13025\ := eclat_unit;
                \$12883\ := eclat_resize(\$12864_copy_root_in_ram6635886_arg\(32 to 47),31) & eclat_false & 
                work.Int.add(\$12864_copy_root_in_ram6635886_arg\(32 to 47), 
                             work.Int.add(eclat_resize(work.Int.lsr(\$13009_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$v6247\ := \$ram_lock\;
                if \$v6247\(0) = '1' then
                  state_var7463 := Q_WAIT6246;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$12864_copy_root_in_ram6635886_arg\(0 to 15)));
                  \$ram_write\ <= \$12883\(0 to 31); \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6245;
                end if;
              when PAUSE_SET6251 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$13024\ := eclat_unit;
                \$v6250\ := \$ram_lock\;
                if \$v6250\(0) = '1' then
                  state_var7463 := Q_WAIT6249;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$12879\(0 to 30),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$12864_copy_root_in_ram6635886_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6248;
                end if;
              when PAUSE_SET6254 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$13022\ := eclat_unit;
                \$12806_loop666_id\ := "000000010111";
                \$12806_loop666_arg\ := X"000" & X"1" & \$12864_copy_root_in_ram6635886_arg\(32 to 47) & eclat_resize(\$12879\(0 to 30),16) & eclat_resize(
                work.Int.lsr(\$13009_hd\(0 to 30), X"0000000" & X"2"),16);
                state_var7463 := \$12806_LOOP666\;
              when PAUSE_SET6272 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$13127\ := eclat_unit;
                \$13128\ := work.Print.print_string(clk,of_string(" next="));
                \$13129\ := work.Int.print(clk,\$13124\(32 to 47));
                \$13130\ := work.Print.print_newline(clk,eclat_unit);
                \$13105_copy_root_in_ram6635884_arg\ := work.Int.add(
                                                        \$13105_copy_root_in_ram6635884_arg\(0 to 15), X"000" & X"1") & \$13105_copy_root_in_ram6635884_arg\(16 to 31) & \$13124\(32 to 47) & \$13105_copy_root_in_ram6635884_arg\(48 to 63) & \$13105_copy_root_in_ram6635884_arg\(64 to 79);
                state_var7463 := \$13105_COPY_ROOT_IN_RAM6635884\;
              when PAUSE_SET6275 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$13159\ := eclat_unit;
                \$13124\ := eclat_resize(\$13105_copy_root_in_ram6635884_arg\(32 to 47),31) & eclat_false & 
                work.Int.add(\$13105_copy_root_in_ram6635884_arg\(32 to 47), 
                             work.Int.add(eclat_resize(work.Int.lsr(\$13143_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$v6274\ := \$ram_lock\;
                if \$v6274\(0) = '1' then
                  state_var7463 := Q_WAIT6273;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13105_copy_root_in_ram6635884_arg\(0 to 15)));
                  \$ram_write\ <= \$13124\(0 to 31); \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6272;
                end if;
              when PAUSE_SET6278 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$13158\ := eclat_unit;
                \$v6277\ := \$ram_lock\;
                if \$v6277\(0) = '1' then
                  state_var7463 := Q_WAIT6276;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$13120\(0 to 30),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$13105_copy_root_in_ram6635884_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6275;
                end if;
              when PAUSE_SET6281 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$13156\ := eclat_unit;
                \$12806_loop666_id\ := "000000011001";
                \$12806_loop666_arg\ := X"000" & X"1" & \$13105_copy_root_in_ram6635884_arg\(32 to 47) & eclat_resize(\$13120\(0 to 30),16) & eclat_resize(
                work.Int.lsr(\$13143_hd\(0 to 30), X"0000000" & X"2"),16);
                state_var7463 := \$12806_LOOP666\;
              when PAUSE_SET6296 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$13100\ := eclat_unit;
                \$13101\ := work.Print.print_string(clk,of_string(" next="));
                \$13102\ := work.Int.print(clk,\$13097\(32 to 47));
                \$13103\ := work.Print.print_newline(clk,eclat_unit);
                \$13105_copy_root_in_ram6635884_id\ := "000000011010";
                \$13105_copy_root_in_ram6635884_arg\ := work.Int.add(
                                                        \$13078_copy_root_in_ram6635885_arg\(0 to 15), X"000" & X"1") & \$13078_copy_root_in_ram6635885_arg\(16 to 31) & \$13097\(32 to 47) & \$13078_copy_root_in_ram6635885_arg\(48 to 63) & \$13078_copy_root_in_ram6635885_arg\(64 to 79);
                state_var7463 := \$13105_COPY_ROOT_IN_RAM6635884\;
              when PAUSE_SET6299 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$13239\ := eclat_unit;
                \$13097\ := eclat_resize(\$13078_copy_root_in_ram6635885_arg\(32 to 47),31) & eclat_false & 
                work.Int.add(\$13078_copy_root_in_ram6635885_arg\(32 to 47), 
                             work.Int.add(eclat_resize(work.Int.lsr(\$13223_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$v6298\ := \$ram_lock\;
                if \$v6298\(0) = '1' then
                  state_var7463 := Q_WAIT6297;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13078_copy_root_in_ram6635885_arg\(0 to 15)));
                  \$ram_write\ <= \$13097\(0 to 31); \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6296;
                end if;
              when PAUSE_SET6302 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$13238\ := eclat_unit;
                \$v6301\ := \$ram_lock\;
                if \$v6301\(0) = '1' then
                  state_var7463 := Q_WAIT6300;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$13093\(0 to 30),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$13078_copy_root_in_ram6635885_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6299;
                end if;
              when PAUSE_SET6305 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$13236\ := eclat_unit;
                \$12806_loop666_id\ := "000000011011";
                \$12806_loop666_arg\ := X"000" & X"1" & \$13078_copy_root_in_ram6635885_arg\(32 to 47) & eclat_resize(\$13093\(0 to 30),16) & eclat_resize(
                work.Int.lsr(\$13223_hd\(0 to 30), X"0000000" & X"2"),16);
                state_var7463 := \$12806_LOOP666\;
              when PAUSE_SET6320 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$13317\ := eclat_unit;
                \$12835\ := eclat_resize(\$12818\(32 to 47),31) & eclat_false & 
                work.Int.add(\$12818\(32 to 47), work.Int.add(eclat_resize(
                                                              work.Int.lsr(
                                                              \$13301_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$13078_copy_root_in_ram6635885_id\ := "000000011100";
                \$13078_copy_root_in_ram6635885_arg\ := X"0" & X"3e8" & \$12681_wait662_arg\(65 to 80) & \$12835\(32 to 47) & \$12792\(96 to 111) & \$12792\(112 to 127);
                state_var7463 := \$13078_COPY_ROOT_IN_RAM6635885\;
              when PAUSE_SET6323 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$13316\ := eclat_unit;
                \$v6322\ := \$ram_lock\;
                if \$v6322\(0) = '1' then
                  state_var7463 := Q_WAIT6321;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$12681_wait662_arg\(33 to 63),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$12818\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6320;
                end if;
              when PAUSE_SET6326 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$13314\ := eclat_unit;
                \$12806_loop666_id\ := "000000011101";
                \$12806_loop666_arg\ := X"000" & X"1" & \$12818\(32 to 47) & eclat_resize(\$12681_wait662_arg\(33 to 63),16) & eclat_resize(
                work.Int.lsr(\$13301_hd\(0 to 30), X"0000000" & X"2"),16);
                state_var7463 := \$12806_LOOP666\;
              when PAUSE_SET6337 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$13395\ := eclat_unit;
                \$12818\ := eclat_resize(\$12792\(112 to 127),31) & eclat_false & 
                work.Int.add(\$12792\(112 to 127), work.Int.add(eclat_resize(
                                                                work.Int.lsr(
                                                                \$13379_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$v6336\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$12681_wait662_arg\(64)) & 
                                           eclat_if(work.Int.le(\$12792\(96 to 111), eclat_resize(\$12681_wait662_arg\(33 to 63),16)) & 
                                           work.Int.lt(eclat_resize(\$12681_wait662_arg\(33 to 63),16), 
                                                       work.Int.add(\$12792\(96 to 111), X"1770")) & eclat_false) & eclat_false));
                if \$v6336\(0) = '1' then
                  \$12835\ := \$12681_wait662_arg\(33 to 64) & \$12818\(32 to 47);
                  \$13078_copy_root_in_ram6635885_id\ := "000000011100";
                  \$13078_copy_root_in_ram6635885_arg\ := X"0" & X"3e8" & \$12681_wait662_arg\(65 to 80) & \$12835\(32 to 47) & \$12792\(96 to 111) & \$12792\(112 to 127);
                  state_var7463 := \$13078_COPY_ROOT_IN_RAM6635885\;
                else
                  \$v6335\ := \$ram_lock\;
                  if \$v6335\(0) = '1' then
                    state_var7463 := Q_WAIT6334;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$12681_wait662_arg\(33 to 63),16), X"000" & X"1")));
                    state_var7463 := PAUSE_GET6333;
                  end if;
                end if;
              when PAUSE_SET6340 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$13394\ := eclat_unit;
                \$v6339\ := \$ram_lock\;
                if \$v6339\(0) = '1' then
                  state_var7463 := Q_WAIT6338;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$12681_wait662_arg\(1 to 31),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$12792\(112 to 127),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6337;
                end if;
              when PAUSE_SET6343 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$13392\ := eclat_unit;
                \$12806_loop666_id\ := "000000011110";
                \$12806_loop666_arg\ := X"000" & X"1" & \$12792\(112 to 127) & eclat_resize(\$12681_wait662_arg\(1 to 31),16) & eclat_resize(
                work.Int.lsr(\$13379_hd\(0 to 30), X"0000000" & X"2"),16);
                state_var7463 := \$12806_LOOP666\;
              when Q_WAIT6151 =>
                \$v6152\ := \$ram_lock\;
                if \$v6152\(0) = '1' then
                  state_var7463 := Q_WAIT6151;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$12803_loop666_arg\(16 to 31), \$12803_loop666_arg\(0 to 15))));
                  \$ram_write\ <= \$13765\; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6150;
                end if;
              when Q_WAIT6154 =>
                \$v6155\ := \$ram_lock\;
                if \$v6155\(0) = '1' then
                  state_var7463 := Q_WAIT6154;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$12803_loop666_arg\(32 to 47), \$12803_loop666_arg\(0 to 15))));
                  state_var7463 := PAUSE_GET6153;
                end if;
              when Q_WAIT6158 =>
                \$v6159\ := \$ram_lock\;
                if \$v6159\(0) = '1' then
                  state_var7463 := Q_WAIT6158;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$12804_loop665_arg\(64 to 79), \$12804_loop665_arg\(0 to 15))));
                  \$ram_write\ <= \$13667\(0 to 31); \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6157;
                end if;
              when Q_WAIT6161 =>
                \$v6162\ := \$ram_lock\;
                if \$v6162\(0) = '1' then
                  state_var7463 := Q_WAIT6161;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$13663\(0 to 30),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$12804_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6160;
                end if;
              when Q_WAIT6164 =>
                \$v6165\ := \$ram_lock\;
                if \$v6165\(0) = '1' then
                  state_var7463 := Q_WAIT6164;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$13663\(0 to 30),16)));
                  \$ram_write\ <= eclat_resize(\$12804_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6163;
                end if;
              when Q_WAIT6167 =>
                \$v6168\ := \$ram_lock\;
                if \$v6168\(0) = '1' then
                  state_var7463 := Q_WAIT6167;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$12804_loop665_arg\(16 to 31)));
                  \$ram_write\ <= \$13684_hd\; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6166;
                end if;
              when Q_WAIT6170 =>
                \$v6171\ := \$ram_lock\;
                if \$v6171\(0) = '1' then
                  state_var7463 := Q_WAIT6170;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$13663\(0 to 30),16)));
                  state_var7463 := PAUSE_GET6169;
                end if;
              when Q_WAIT6174 =>
                \$v6175\ := \$ram_lock\;
                if \$v6175\(0) = '1' then
                  state_var7463 := Q_WAIT6174;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$13663\(0 to 30),16), X"000" & X"1")));
                  state_var7463 := PAUSE_GET6173;
                end if;
              when Q_WAIT6178 =>
                \$v6179\ := \$ram_lock\;
                if \$v6179\(0) = '1' then
                  state_var7463 := Q_WAIT6178;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$12804_loop665_arg\(64 to 79), \$12804_loop665_arg\(0 to 15))));
                  state_var7463 := PAUSE_GET6177;
                end if;
              when Q_WAIT6182 =>
                \$v6183\ := \$ram_lock\;
                if \$v6183\(0) = '1' then
                  state_var7463 := Q_WAIT6182;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(\$12805_aux664_arg\(0 to 15)));
                  state_var7463 := PAUSE_GET6181;
                end if;
              when Q_WAIT6186 =>
                \$v6187\ := \$ram_lock\;
                if \$v6187\(0) = '1' then
                  state_var7463 := Q_WAIT6186;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$12806_loop666_arg\(16 to 31), \$12806_loop666_arg\(0 to 15))));
                  \$ram_write\ <= \$13605\; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6185;
                end if;
              when Q_WAIT6189 =>
                \$v6190\ := \$ram_lock\;
                if \$v6190\(0) = '1' then
                  state_var7463 := Q_WAIT6189;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$12806_loop666_arg\(32 to 47), \$12806_loop666_arg\(0 to 15))));
                  state_var7463 := PAUSE_GET6188;
                end if;
              when Q_WAIT6193 =>
                \$v6194\ := \$ram_lock\;
                if \$v6194\(0) = '1' then
                  state_var7463 := Q_WAIT6193;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$12807_loop665_arg\(64 to 79), \$12807_loop665_arg\(0 to 15))));
                  \$ram_write\ <= \$13507\(0 to 31); \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6192;
                end if;
              when Q_WAIT6196 =>
                \$v6197\ := \$ram_lock\;
                if \$v6197\(0) = '1' then
                  state_var7463 := Q_WAIT6196;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$13503\(0 to 30),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$12807_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6195;
                end if;
              when Q_WAIT6199 =>
                \$v6200\ := \$ram_lock\;
                if \$v6200\(0) = '1' then
                  state_var7463 := Q_WAIT6199;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$13503\(0 to 30),16)));
                  \$ram_write\ <= eclat_resize(\$12807_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6198;
                end if;
              when Q_WAIT6202 =>
                \$v6203\ := \$ram_lock\;
                if \$v6203\(0) = '1' then
                  state_var7463 := Q_WAIT6202;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$12807_loop665_arg\(16 to 31)));
                  \$ram_write\ <= \$13524_hd\; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6201;
                end if;
              when Q_WAIT6205 =>
                \$v6206\ := \$ram_lock\;
                if \$v6206\(0) = '1' then
                  state_var7463 := Q_WAIT6205;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$13503\(0 to 30),16)));
                  state_var7463 := PAUSE_GET6204;
                end if;
              when Q_WAIT6209 =>
                \$v6210\ := \$ram_lock\;
                if \$v6210\(0) = '1' then
                  state_var7463 := Q_WAIT6209;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$13503\(0 to 30),16), X"000" & X"1")));
                  state_var7463 := PAUSE_GET6208;
                end if;
              when Q_WAIT6213 =>
                \$v6214\ := \$ram_lock\;
                if \$v6214\(0) = '1' then
                  state_var7463 := Q_WAIT6213;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$12807_loop665_arg\(64 to 79), \$12807_loop665_arg\(0 to 15))));
                  state_var7463 := PAUSE_GET6212;
                end if;
              when Q_WAIT6217 =>
                \$v6218\ := \$ram_lock\;
                if \$v6218\(0) = '1' then
                  state_var7463 := Q_WAIT6217;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(\$12808_aux664_arg\(0 to 15)));
                  state_var7463 := PAUSE_GET6216;
                end if;
              when Q_WAIT6222 =>
                \$v6223\ := \$ram_lock\;
                if \$v6223\(0) = '1' then
                  state_var7463 := Q_WAIT6222;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$12891_copy_root_in_ram6635884_arg\(0 to 15)));
                  \$ram_write\ <= \$12910\(0 to 31); \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6221;
                end if;
              when Q_WAIT6225 =>
                \$v6226\ := \$ram_lock\;
                if \$v6226\(0) = '1' then
                  state_var7463 := Q_WAIT6225;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$12906\(0 to 30),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$12891_copy_root_in_ram6635884_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6224;
                end if;
              when Q_WAIT6228 =>
                \$v6229\ := \$ram_lock\;
                if \$v6229\(0) = '1' then
                  state_var7463 := Q_WAIT6228;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$12906\(0 to 30),16)));
                  \$ram_write\ <= eclat_resize(\$12891_copy_root_in_ram6635884_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6227;
                end if;
              when Q_WAIT6231 =>
                \$v6232\ := \$ram_lock\;
                if \$v6232\(0) = '1' then
                  state_var7463 := Q_WAIT6231;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$12891_copy_root_in_ram6635884_arg\(32 to 47)));
                  \$ram_write\ <= \$12929_hd\; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6230;
                end if;
              when Q_WAIT6234 =>
                \$v6235\ := \$ram_lock\;
                if \$v6235\(0) = '1' then
                  state_var7463 := Q_WAIT6234;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$12906\(0 to 30),16)));
                  state_var7463 := PAUSE_GET6233;
                end if;
              when Q_WAIT6238 =>
                \$v6239\ := \$ram_lock\;
                if \$v6239\(0) = '1' then
                  state_var7463 := Q_WAIT6238;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$12906\(0 to 30),16), X"000" & X"1")));
                  state_var7463 := PAUSE_GET6237;
                end if;
              when Q_WAIT6242 =>
                \$v6243\ := \$ram_lock\;
                if \$v6243\(0) = '1' then
                  state_var7463 := Q_WAIT6242;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(\$12891_copy_root_in_ram6635884_arg\(0 to 15)));
                  state_var7463 := PAUSE_GET6241;
                end if;
              when Q_WAIT6246 =>
                \$v6247\ := \$ram_lock\;
                if \$v6247\(0) = '1' then
                  state_var7463 := Q_WAIT6246;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$12864_copy_root_in_ram6635886_arg\(0 to 15)));
                  \$ram_write\ <= \$12883\(0 to 31); \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6245;
                end if;
              when Q_WAIT6249 =>
                \$v6250\ := \$ram_lock\;
                if \$v6250\(0) = '1' then
                  state_var7463 := Q_WAIT6249;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$12879\(0 to 30),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$12864_copy_root_in_ram6635886_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6248;
                end if;
              when Q_WAIT6252 =>
                \$v6253\ := \$ram_lock\;
                if \$v6253\(0) = '1' then
                  state_var7463 := Q_WAIT6252;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$12879\(0 to 30),16)));
                  \$ram_write\ <= eclat_resize(\$12864_copy_root_in_ram6635886_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6251;
                end if;
              when Q_WAIT6255 =>
                \$v6256\ := \$ram_lock\;
                if \$v6256\(0) = '1' then
                  state_var7463 := Q_WAIT6255;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$12864_copy_root_in_ram6635886_arg\(32 to 47)));
                  \$ram_write\ <= \$13009_hd\; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6254;
                end if;
              when Q_WAIT6258 =>
                \$v6259\ := \$ram_lock\;
                if \$v6259\(0) = '1' then
                  state_var7463 := Q_WAIT6258;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$12879\(0 to 30),16)));
                  state_var7463 := PAUSE_GET6257;
                end if;
              when Q_WAIT6262 =>
                \$v6263\ := \$ram_lock\;
                if \$v6263\(0) = '1' then
                  state_var7463 := Q_WAIT6262;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$12879\(0 to 30),16), X"000" & X"1")));
                  state_var7463 := PAUSE_GET6261;
                end if;
              when Q_WAIT6266 =>
                \$v6267\ := \$ram_lock\;
                if \$v6267\(0) = '1' then
                  state_var7463 := Q_WAIT6266;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(\$12864_copy_root_in_ram6635886_arg\(0 to 15)));
                  state_var7463 := PAUSE_GET6265;
                end if;
              when Q_WAIT6270 =>
                \$v6271\ := \$global_end_lock\;
                if \$v6271\(0) = '1' then
                  state_var7463 := Q_WAIT6270;
                else
                  acquire(\$global_end_lock\);
                  \$global_end_ptr\ <= 0;
                  state_var7463 := PAUSE_GET6269;
                end if;
              when Q_WAIT6273 =>
                \$v6274\ := \$ram_lock\;
                if \$v6274\(0) = '1' then
                  state_var7463 := Q_WAIT6273;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13105_copy_root_in_ram6635884_arg\(0 to 15)));
                  \$ram_write\ <= \$13124\(0 to 31); \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6272;
                end if;
              when Q_WAIT6276 =>
                \$v6277\ := \$ram_lock\;
                if \$v6277\(0) = '1' then
                  state_var7463 := Q_WAIT6276;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$13120\(0 to 30),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$13105_copy_root_in_ram6635884_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6275;
                end if;
              when Q_WAIT6279 =>
                \$v6280\ := \$ram_lock\;
                if \$v6280\(0) = '1' then
                  state_var7463 := Q_WAIT6279;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$13120\(0 to 30),16)));
                  \$ram_write\ <= eclat_resize(\$13105_copy_root_in_ram6635884_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6278;
                end if;
              when Q_WAIT6282 =>
                \$v6283\ := \$ram_lock\;
                if \$v6283\(0) = '1' then
                  state_var7463 := Q_WAIT6282;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13105_copy_root_in_ram6635884_arg\(32 to 47)));
                  \$ram_write\ <= \$13143_hd\; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6281;
                end if;
              when Q_WAIT6285 =>
                \$v6286\ := \$ram_lock\;
                if \$v6286\(0) = '1' then
                  state_var7463 := Q_WAIT6285;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$13120\(0 to 30),16)));
                  state_var7463 := PAUSE_GET6284;
                end if;
              when Q_WAIT6289 =>
                \$v6290\ := \$ram_lock\;
                if \$v6290\(0) = '1' then
                  state_var7463 := Q_WAIT6289;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$13120\(0 to 30),16), X"000" & X"1")));
                  state_var7463 := PAUSE_GET6288;
                end if;
              when Q_WAIT6293 =>
                \$v6294\ := \$ram_lock\;
                if \$v6294\(0) = '1' then
                  state_var7463 := Q_WAIT6293;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(\$13105_copy_root_in_ram6635884_arg\(0 to 15)));
                  state_var7463 := PAUSE_GET6292;
                end if;
              when Q_WAIT6297 =>
                \$v6298\ := \$ram_lock\;
                if \$v6298\(0) = '1' then
                  state_var7463 := Q_WAIT6297;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13078_copy_root_in_ram6635885_arg\(0 to 15)));
                  \$ram_write\ <= \$13097\(0 to 31); \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6296;
                end if;
              when Q_WAIT6300 =>
                \$v6301\ := \$ram_lock\;
                if \$v6301\(0) = '1' then
                  state_var7463 := Q_WAIT6300;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$13093\(0 to 30),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$13078_copy_root_in_ram6635885_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6299;
                end if;
              when Q_WAIT6303 =>
                \$v6304\ := \$ram_lock\;
                if \$v6304\(0) = '1' then
                  state_var7463 := Q_WAIT6303;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$13093\(0 to 30),16)));
                  \$ram_write\ <= eclat_resize(\$13078_copy_root_in_ram6635885_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6302;
                end if;
              when Q_WAIT6306 =>
                \$v6307\ := \$ram_lock\;
                if \$v6307\(0) = '1' then
                  state_var7463 := Q_WAIT6306;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13078_copy_root_in_ram6635885_arg\(32 to 47)));
                  \$ram_write\ <= \$13223_hd\; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6305;
                end if;
              when Q_WAIT6309 =>
                \$v6310\ := \$ram_lock\;
                if \$v6310\(0) = '1' then
                  state_var7463 := Q_WAIT6309;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$13093\(0 to 30),16)));
                  state_var7463 := PAUSE_GET6308;
                end if;
              when Q_WAIT6313 =>
                \$v6314\ := \$ram_lock\;
                if \$v6314\(0) = '1' then
                  state_var7463 := Q_WAIT6313;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$13093\(0 to 30),16), X"000" & X"1")));
                  state_var7463 := PAUSE_GET6312;
                end if;
              when Q_WAIT6317 =>
                \$v6318\ := \$ram_lock\;
                if \$v6318\(0) = '1' then
                  state_var7463 := Q_WAIT6317;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(\$13078_copy_root_in_ram6635885_arg\(0 to 15)));
                  state_var7463 := PAUSE_GET6316;
                end if;
              when Q_WAIT6321 =>
                \$v6322\ := \$ram_lock\;
                if \$v6322\(0) = '1' then
                  state_var7463 := Q_WAIT6321;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$12681_wait662_arg\(33 to 63),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$12818\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6320;
                end if;
              when Q_WAIT6324 =>
                \$v6325\ := \$ram_lock\;
                if \$v6325\(0) = '1' then
                  state_var7463 := Q_WAIT6324;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$12681_wait662_arg\(33 to 63),16)));
                  \$ram_write\ <= eclat_resize(\$12818\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6323;
                end if;
              when Q_WAIT6327 =>
                \$v6328\ := \$ram_lock\;
                if \$v6328\(0) = '1' then
                  state_var7463 := Q_WAIT6327;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$12818\(32 to 47)));
                  \$ram_write\ <= \$13301_hd\; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6326;
                end if;
              when Q_WAIT6330 =>
                \$v6331\ := \$ram_lock\;
                if \$v6331\(0) = '1' then
                  state_var7463 := Q_WAIT6330;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$12681_wait662_arg\(33 to 63),16)));
                  state_var7463 := PAUSE_GET6329;
                end if;
              when Q_WAIT6334 =>
                \$v6335\ := \$ram_lock\;
                if \$v6335\(0) = '1' then
                  state_var7463 := Q_WAIT6334;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$12681_wait662_arg\(33 to 63),16), X"000" & X"1")));
                  state_var7463 := PAUSE_GET6333;
                end if;
              when Q_WAIT6338 =>
                \$v6339\ := \$ram_lock\;
                if \$v6339\(0) = '1' then
                  state_var7463 := Q_WAIT6338;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$12681_wait662_arg\(1 to 31),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$12792\(112 to 127),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6337;
                end if;
              when Q_WAIT6341 =>
                \$v6342\ := \$ram_lock\;
                if \$v6342\(0) = '1' then
                  state_var7463 := Q_WAIT6341;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$12681_wait662_arg\(1 to 31),16)));
                  \$ram_write\ <= eclat_resize(\$12792\(112 to 127),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6340;
                end if;
              when Q_WAIT6344 =>
                \$v6345\ := \$ram_lock\;
                if \$v6345\(0) = '1' then
                  state_var7463 := Q_WAIT6344;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$12792\(112 to 127)));
                  \$ram_write\ <= \$13379_hd\; \$ram_write_request\ <= '1';
                  state_var7463 := PAUSE_SET6343;
                end if;
              when Q_WAIT6347 =>
                \$v6348\ := \$ram_lock\;
                if \$v6348\(0) = '1' then
                  state_var7463 := Q_WAIT6347;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$12681_wait662_arg\(1 to 31),16)));
                  state_var7463 := PAUSE_GET6346;
                end if;
              when Q_WAIT6351 =>
                \$v6352\ := \$ram_lock\;
                if \$v6352\(0) = '1' then
                  state_var7463 := Q_WAIT6351;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$12681_wait662_arg\(1 to 31),16), X"000" & X"1")));
                  state_var7463 := PAUSE_GET6350;
                end if;
              when IDLE6149 =>
                rdy6148 := eclat_false;
                \$v6354\ := work.Int.gt(work.Int.add(\$12792\(80 to 95), \$12681_wait662_arg\(81 to 96)), 
                                        work.Int.add(\$12792\(96 to 111), X"1770"));
                if \$v6354\(0) = '1' then
                  \$12811\ := work.Print.print_newline(clk,eclat_unit);
                  \$12812\ := work.Print.print_newline(clk,eclat_unit);
                  \$12813\ := work.Print.print_string(clk,of_string("[================= GC START ======================]"));
                  \$13448\ := work.Print.print_newline(clk,eclat_unit);
                  \$12814\ := work.Print.print_newline(clk,eclat_unit);
                  \$v6353\ := work.Bool.lnot(eclat_if(work.Bool.lnot(
                                                      ""&\$12681_wait662_arg\(32)) & 
                                             eclat_if(work.Int.le(\$12792\(96 to 111), eclat_resize(\$12681_wait662_arg\(1 to 31),16)) & 
                                             work.Int.lt(eclat_resize(\$12681_wait662_arg\(1 to 31),16), 
                                                         work.Int.add(
                                                         \$12792\(96 to 111), X"1770")) & eclat_false) & eclat_false));
                  if \$v6353\(0) = '1' then
                    \$12818\ := \$12681_wait662_arg\(1 to 32) & \$12792\(112 to 127);
                    \$v6336\ := work.Bool.lnot(eclat_if(work.Bool.lnot(
                                                        ""&\$12681_wait662_arg\(64)) & 
                                               eclat_if(work.Int.le(\$12792\(96 to 111), eclat_resize(\$12681_wait662_arg\(33 to 63),16)) & 
                                               work.Int.lt(eclat_resize(\$12681_wait662_arg\(33 to 63),16), 
                                                           work.Int.add(
                                                           \$12792\(96 to 111), X"1770")) & eclat_false) & eclat_false));
                    if \$v6336\(0) = '1' then
                      \$12835\ := \$12681_wait662_arg\(33 to 64) & \$12818\(32 to 47);
                      \$13078_copy_root_in_ram6635885_id\ := "000000011100";
                      \$13078_copy_root_in_ram6635885_arg\ := X"0" & X"3e8" & \$12681_wait662_arg\(65 to 80) & \$12835\(32 to 47) & \$12792\(96 to 111) & \$12792\(112 to 127);
                      state_var7463 := \$13078_COPY_ROOT_IN_RAM6635885\;
                    else
                      \$v6335\ := \$ram_lock\;
                      if \$v6335\(0) = '1' then
                        state_var7463 := Q_WAIT6334;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$12681_wait662_arg\(33 to 63),16), X"000" & X"1")));
                        state_var7463 := PAUSE_GET6333;
                      end if;
                    end if;
                  else
                    \$v6352\ := \$ram_lock\;
                    if \$v6352\(0) = '1' then
                      state_var7463 := Q_WAIT6351;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                        eclat_resize(\$12681_wait662_arg\(1 to 31),16), X"000" & X"1")));
                      state_var7463 := PAUSE_GET6350;
                    end if;
                  end if;
                else
                  result6147 := \$12681_wait662_arg\(1 to 32) & \$12681_wait662_arg\(33 to 64) & \$12792\(80 to 95) & 
                  work.Int.add(\$12792\(80 to 95), \$12681_wait662_arg\(81 to 96)) & \$12792\(96 to 111) & \$12792\(112 to 127);
                  rdy6148 := eclat_true;
                  state_var7463 := IDLE6149;
                end if;
              end case;
              
              if rdy6148(0) = '1' then
                
              else
                result6147 := \$12792\(0 to 31) & \$12792\(32 to 63) & \$12792\(64 to 79) & \$12792\(80 to 95) & \$12792\(96 to 111) & \$12792\(112 to 127);
              end if;
              \$12792\ := result6147 & rdy6148;
              \$12782\ := \$12792\;
              \$v6146\ := ""&\$12782\(128);
              if \$v6146\(0) = '1' then
                \$12681_wait662_result\ := \$12782\(0 to 31) & \$12782\(32 to 63) & \$12782\(64 to 79);
                \$12737\ := \$12681_wait662_result\;
                \$12741\ := work.Print.print_string(clk,of_string("size:"));
                \$12742\ := work.Int.print(clk,eclat_if(work.Int.eq(\$12682_make_block579_arg\(112 to 127), X"000" & X"0") & X"000" & X"1" & \$12682_make_block579_arg\(112 to 127)));
                \$12743\ := work.Print.print_newline(clk,eclat_unit);
                \$v6358\ := \$ram_lock\;
                if \$v6358\(0) = '1' then
                  state_var7462 := Q_WAIT6357;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$12737\(64 to 79)));
                  \$ram_write\ <= work.Int.lor(work.Int.lsl(eclat_resize(\$12682_make_block579_arg\(80 to 111),31), X"000000" & X"18"), 
                                               work.Int.lsl(eclat_resize(
                                                            eclat_if(
                                                            work.Int.eq(
                                                            \$12682_make_block579_arg\(112 to 127), X"000" & X"0") & X"000" & X"1" & \$12682_make_block579_arg\(112 to 127)),31), X"0000000" & X"2")) & eclat_true; \$ram_write_request\ <= '1';
                  state_var7462 := PAUSE_SET6356;
                end if;
              else
                \$12681_wait662_arg\ := eclat_unit & \$12681_wait662_arg\(1 to 32) & \$12681_wait662_arg\(33 to 64) & \$12681_wait662_arg\(65 to 80) & \$12681_wait662_arg\(81 to 96);
                state_var7462 := \$12681_WAIT662\;
              end if;
            when \$12682_MAKE_BLOCK579\ =>
              \$12734\ := work.Print.print_string(clk,of_string("GC-ALLOC:(size="));
              \$12735\ := work.Int.print(clk,work.Int.add(eclat_if(work.Int.eq(
                                                                   \$12682_make_block579_arg\(112 to 127), X"000" & X"0") & X"000" & X"1" & \$12682_make_block579_arg\(112 to 127)), X"000" & X"1"));
              \$12736\ := work.Print.print_string(clk,of_string(")"));
              \$12760\ := work.Print.print_newline(clk,eclat_unit);
              \$12681_wait662_id\ := "000000011111";
              \$12681_wait662_arg\ := eclat_unit & \$12682_make_block579_arg\(16 to 47) & \$12682_make_block579_arg\(48 to 79) & \$12682_make_block579_arg\(0 to 15) & 
              work.Int.add(eclat_if(work.Int.eq(\$12682_make_block579_arg\(112 to 127), X"000" & X"0") & X"000" & X"1" & \$12682_make_block579_arg\(112 to 127)), X"000" & X"1");
              state_var7462 := \$12681_WAIT662\;
            when PAUSE_GET6118 =>
              \$13889\ := \$ram_value\;
              release(\$ram_lock\);
              \$v6117\ := \$ram_lock\;
              if \$v6117\(0) = '1' then
                state_var7462 := Q_WAIT6116;
              else
                acquire(\$ram_lock\);
                \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                        \$12679_loop666_arg\(16 to 31), \$12679_loop666_arg\(0 to 15))));
                \$ram_write\ <= \$13889\; \$ram_write_request\ <= '1';
                state_var7462 := PAUSE_SET6115;
              end if;
            when PAUSE_GET6134 =>
              \$13808_hd\ := \$ram_value\;
              release(\$ram_lock\);
              \$13812\ := work.Print.print_string(clk,of_string("bloc "));
              \$13813\ := work.Int.print(clk,eclat_resize(\$13787\(0 to 30),16));
              \$13814\ := work.Print.print_string(clk,of_string(" of size "));
              \$13815\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                          work.Int.lsr(
                                                          \$13808_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
              \$13816\ := work.Print.print_string(clk,of_string(" from "));
              \$13817\ := work.Int.print(clk,eclat_resize(\$13787\(0 to 30),16));
              \$13818\ := work.Print.print_string(clk,of_string(" to "));
              \$13819\ := work.Int.print(clk,\$12680_loop665_arg\(16 to 31));
              \$13820\ := work.Print.print_newline(clk,eclat_unit);
              \$v6133\ := \$ram_lock\;
              if \$v6133\(0) = '1' then
                state_var7462 := Q_WAIT6132;
              else
                acquire(\$ram_lock\);
                \$ram_ptr_write\ <= to_integer(unsigned(\$12680_loop665_arg\(16 to 31)));
                \$ram_write\ <= \$13808_hd\; \$ram_write_request\ <= '1';
                state_var7462 := PAUSE_SET6131;
              end if;
            when PAUSE_GET6138 =>
              \$13803_w\ := \$ram_value\;
              release(\$ram_lock\);
              \$v6137\ := eclat_if(work.Bool.lnot(""&\$13803_w\(31)) & 
                          eclat_if(work.Int.le(\$12680_loop665_arg\(48 to 63), eclat_resize(\$13803_w\(0 to 30),16)) & 
                          work.Int.lt(eclat_resize(\$13803_w\(0 to 30),16), 
                                      work.Int.add(\$12680_loop665_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false);
              if \$v6137\(0) = '1' then
                \$13791\ := \$13803_w\ & \$12680_loop665_arg\(16 to 31);
                \$v6124\ := \$ram_lock\;
                if \$v6124\(0) = '1' then
                  state_var7462 := Q_WAIT6123;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$12680_loop665_arg\(64 to 79), \$12680_loop665_arg\(0 to 15))));
                  \$ram_write\ <= \$13791\(0 to 31); \$ram_write_request\ <= '1';
                  state_var7462 := PAUSE_SET6122;
                end if;
              else
                \$v6136\ := \$ram_lock\;
                if \$v6136\(0) = '1' then
                  state_var7462 := Q_WAIT6135;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$13787\(0 to 30),16)));
                  state_var7462 := PAUSE_GET6134;
                end if;
              end if;
            when PAUSE_GET6142 =>
              \$13787\ := \$ram_value\;
              release(\$ram_lock\);
              \$v6141\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$13787\(31)) & 
                                         eclat_if(work.Int.le(\$12680_loop665_arg\(32 to 47), eclat_resize(\$13787\(0 to 30),16)) & 
                                         work.Int.lt(eclat_resize(\$13787\(0 to 30),16), 
                                                     work.Int.add(\$12680_loop665_arg\(32 to 47), X"1770")) & eclat_false) & eclat_false));
              if \$v6141\(0) = '1' then
                \$13791\ := \$13787\ & \$12680_loop665_arg\(16 to 31);
                \$v6124\ := \$ram_lock\;
                if \$v6124\(0) = '1' then
                  state_var7462 := Q_WAIT6123;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$12680_loop665_arg\(64 to 79), \$12680_loop665_arg\(0 to 15))));
                  \$ram_write\ <= \$13791\(0 to 31); \$ram_write_request\ <= '1';
                  state_var7462 := PAUSE_SET6122;
                end if;
              else
                \$v6140\ := \$ram_lock\;
                if \$v6140\(0) = '1' then
                  state_var7462 := Q_WAIT6139;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$13787\(0 to 30),16), X"000" & X"1")));
                  state_var7462 := PAUSE_GET6138;
                end if;
              end if;
            when PAUSE_SET6115 =>
              \$ram_write_request\ <= '0';
              release(\$ram_lock\);
              \$13890\ := eclat_unit;
              \$12679_loop666_arg\ := work.Int.add(\$12679_loop666_arg\(0 to 15), X"000" & X"1") & \$12679_loop666_arg\(16 to 31) & \$12679_loop666_arg\(32 to 47) & \$12679_loop666_arg\(48 to 63);
              state_var7462 := \$12679_LOOP666\;
            when PAUSE_SET6122 =>
              \$ram_write_request\ <= '0';
              release(\$ram_lock\);
              \$13794\ := eclat_unit;
              \$12680_loop665_arg\ := work.Int.add(\$12680_loop665_arg\(0 to 15), X"000" & X"1") & \$13791\(32 to 47) & \$12680_loop665_arg\(32 to 47) & \$12680_loop665_arg\(48 to 63) & \$12680_loop665_arg\(64 to 79) & \$12680_loop665_arg\(80 to 95);
              state_var7462 := \$12680_LOOP665\;
            when PAUSE_SET6125 =>
              \$ram_write_request\ <= '0';
              release(\$ram_lock\);
              \$13824\ := eclat_unit;
              \$13791\ := eclat_resize(\$12680_loop665_arg\(16 to 31),31) & eclat_false & 
              work.Int.add(\$12680_loop665_arg\(16 to 31), work.Int.add(
                                                           eclat_resize(
                                                           work.Int.lsr(
                                                           \$13808_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
              \$v6124\ := \$ram_lock\;
              if \$v6124\(0) = '1' then
                state_var7462 := Q_WAIT6123;
              else
                acquire(\$ram_lock\);
                \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                        \$12680_loop665_arg\(64 to 79), \$12680_loop665_arg\(0 to 15))));
                \$ram_write\ <= \$13791\(0 to 31); \$ram_write_request\ <= '1';
                state_var7462 := PAUSE_SET6122;
              end if;
            when PAUSE_SET6128 =>
              \$ram_write_request\ <= '0';
              release(\$ram_lock\);
              \$13823\ := eclat_unit;
              \$v6127\ := \$ram_lock\;
              if \$v6127\(0) = '1' then
                state_var7462 := Q_WAIT6126;
              else
                acquire(\$ram_lock\);
                \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                        eclat_resize(\$13787\(0 to 30),16), X"000" & X"1")));
                \$ram_write\ <= eclat_resize(\$12680_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                state_var7462 := PAUSE_SET6125;
              end if;
            when PAUSE_SET6131 =>
              \$ram_write_request\ <= '0';
              release(\$ram_lock\);
              \$13821\ := eclat_unit;
              \$12679_loop666_id\ := "000000001101";
              \$12679_loop666_arg\ := X"000" & X"1" & \$12680_loop665_arg\(16 to 31) & eclat_resize(\$13787\(0 to 30),16) & eclat_resize(
              work.Int.lsr(\$13808_hd\(0 to 30), X"0000000" & X"2"),16);
              state_var7462 := \$12679_LOOP666\;
            when PAUSE_SET6356 =>
              \$ram_write_request\ <= '0';
              release(\$ram_lock\);
              \$12744\ := eclat_unit;
              \$12682_make_block579_result\ := \$12737\(0 to 31) & \$12737\(32 to 63) & eclat_resize(\$12737\(64 to 79),31) & eclat_false;
              state_var7462 := \$12682_MAKE_BLOCK579\;
            when PAUSE_SET6359 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12721\ := eclat_unit;
              result6112 := eclat_unit;
              rdy6113 := eclat_true;
              state_var7462 := IDLE6114;
            when PAUSE_SET6362 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12720\ := eclat_unit;
              \$v6361\ := \$code_lock\;
              if \$v6361\(0) = '1' then
                state_var7462 := Q_WAIT6360;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 34;\$code_write\ <= "000"& X"00000" & X"8f"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6359;
              end if;
            when PAUSE_SET6365 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12719\ := eclat_unit;
              \$v6364\ := \$code_lock\;
              if \$v6364\(0) = '1' then
                state_var7462 := Q_WAIT6363;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 33;\$code_write\ <= "000"& X"000000" & X"1"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6362;
              end if;
            when PAUSE_SET6368 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12718\ := eclat_unit;
              \$v6367\ := \$code_lock\;
              if \$v6367\(0) = '1' then
                state_var7462 := Q_WAIT6366;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 32;\$code_write\ <= "000"& X"00000" & X"13"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6365;
              end if;
            when PAUSE_SET6371 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12717\ := eclat_unit;
              \$v6370\ := \$code_lock\;
              if \$v6370\(0) = '1' then
                state_var7462 := Q_WAIT6369;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 31;\$code_write\ <= "000"& X"000000" & X"0"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6368;
              end if;
            when PAUSE_SET6374 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12716\ := eclat_unit;
              \$v6373\ := \$code_lock\;
              if \$v6373\(0) = '1' then
                state_var7462 := Q_WAIT6372;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 30;\$code_write\ <= "000"& X"00000" & X"5d"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6371;
              end if;
            when PAUSE_SET6377 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12715\ := eclat_unit;
              \$v6376\ := \$code_lock\;
              if \$v6376\(0) = '1' then
                state_var7462 := Q_WAIT6375;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 29;\$code_write\ <= "000"& X"00000" & X"21"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6374;
              end if;
            when PAUSE_SET6380 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12714\ := eclat_unit;
              \$v6379\ := \$code_lock\;
              if \$v6379\(0) = '1' then
                state_var7462 := Q_WAIT6378;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 28;\$code_write\ <= "000"& X"000000" & X"b"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6377;
              end if;
            when PAUSE_SET6383 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12713\ := eclat_unit;
              \$v6382\ := \$code_lock\;
              if \$v6382\(0) = '1' then
                state_var7462 := Q_WAIT6381;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 27;\$code_write\ <= "000"& X"000000" & X"b"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6380;
              end if;
            when PAUSE_SET6386 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12712\ := eclat_unit;
              \$v6385\ := \$code_lock\;
              if \$v6385\(0) = '1' then
                state_var7462 := Q_WAIT6384;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 26;\$code_write\ <= "000"& X"00000" & X"67"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6383;
              end if;
            when PAUSE_SET6389 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12711\ := eclat_unit;
              \$v6388\ := \$code_lock\;
              if \$v6388\(0) = '1' then
                state_var7462 := Q_WAIT6387;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 25;\$code_write\ <= work.Int.neg(
                                                         "000"& X"00000" & X"17"); \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6386;
              end if;
            when PAUSE_SET6392 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12710\ := eclat_unit;
              \$v6391\ := \$code_lock\;
              if \$v6391\(0) = '1' then
                state_var7462 := Q_WAIT6390;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 24;\$code_write\ <= "000"& X"000000" & X"0"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6389;
              end if;
            when PAUSE_SET6395 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12709\ := eclat_unit;
              \$v6394\ := \$code_lock\;
              if \$v6394\(0) = '1' then
                state_var7462 := Q_WAIT6393;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 23;\$code_write\ <= "000"& X"000000" & X"1"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6392;
              end if;
            when PAUSE_SET6398 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12708\ := eclat_unit;
              \$v6397\ := \$code_lock\;
              if \$v6397\(0) = '1' then
                state_var7462 := Q_WAIT6396;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 22;\$code_write\ <= "000"& X"00000" & X"2c"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6395;
              end if;
            when PAUSE_SET6401 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12707\ := eclat_unit;
              \$v6400\ := \$code_lock\;
              if \$v6400\(0) = '1' then
                state_var7462 := Q_WAIT6399;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 21;\$code_write\ <= "000"& X"000000" & X"1"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6398;
              end if;
            when PAUSE_SET6404 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12706\ := eclat_unit;
              \$v6403\ := \$code_lock\;
              if \$v6403\(0) = '1' then
                state_var7462 := Q_WAIT6402;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 20;\$code_write\ <= "000"& X"00000" & X"28"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6401;
              end if;
            when PAUSE_SET6407 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12705\ := eclat_unit;
              \$v6406\ := \$code_lock\;
              if \$v6406\(0) = '1' then
                state_var7462 := Q_WAIT6405;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 19;\$code_write\ <= "000"& X"00000" & X"6e"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6404;
              end if;
            when PAUSE_SET6410 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12704\ := eclat_unit;
              \$v6409\ := \$code_lock\;
              if \$v6409\(0) = '1' then
                state_var7462 := Q_WAIT6408;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 18;\$code_write\ <= "000"& X"00000" & X"21"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6407;
              end if;
            when PAUSE_SET6413 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12703\ := eclat_unit;
              \$v6412\ := \$code_lock\;
              if \$v6412\(0) = '1' then
                state_var7462 := Q_WAIT6411;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 17;\$code_write\ <= "000"& X"00000" & X"32"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6410;
              end if;
            when PAUSE_SET6416 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12702\ := eclat_unit;
              \$v6415\ := \$code_lock\;
              if \$v6415\(0) = '1' then
                state_var7462 := Q_WAIT6414;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 16;\$code_write\ <= work.Int.neg(
                                                         "000"& X"000000" & X"1"); \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6413;
              end if;
            when PAUSE_SET6419 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12701\ := eclat_unit;
              \$v6418\ := \$code_lock\;
              if \$v6418\(0) = '1' then
                state_var7462 := Q_WAIT6417;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 15;\$code_write\ <= "000"& X"00000" & X"7f"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6416;
              end if;
            when PAUSE_SET6422 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12700\ := eclat_unit;
              \$v6421\ := \$code_lock\;
              if \$v6421\(0) = '1' then
                state_var7462 := Q_WAIT6420;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 14;\$code_write\ <= "000"& X"000000" & X"b"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6419;
              end if;
            when PAUSE_SET6425 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12699\ := eclat_unit;
              \$v6424\ := \$code_lock\;
              if \$v6424\(0) = '1' then
                state_var7462 := Q_WAIT6423;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 13;\$code_write\ <= "000"& X"00000" & X"21"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6422;
              end if;
            when PAUSE_SET6428 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12698\ := eclat_unit;
              \$v6427\ := \$code_lock\;
              if \$v6427\(0) = '1' then
                state_var7462 := Q_WAIT6426;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 12;\$code_write\ <= "000"& X"00000" & X"32"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6425;
              end if;
            when PAUSE_SET6431 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12697\ := eclat_unit;
              \$v6430\ := \$code_lock\;
              if \$v6430\(0) = '1' then
                state_var7462 := Q_WAIT6429;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 11;\$code_write\ <= work.Int.neg(
                                                         "000"& X"000000" & X"2"); \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6428;
              end if;
            when PAUSE_SET6434 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12696\ := eclat_unit;
              \$v6433\ := \$code_lock\;
              if \$v6433\(0) = '1' then
                state_var7462 := Q_WAIT6432;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 10;\$code_write\ <= "000"& X"00000" & X"7f"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6431;
              end if;
            when PAUSE_SET6437 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12695\ := eclat_unit;
              \$v6436\ := \$code_lock\;
              if \$v6436\(0) = '1' then
                state_var7462 := Q_WAIT6435;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 9;\$code_write\ <= "000"& X"000000" & X"0"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6434;
              end if;
            when PAUSE_SET6440 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12694\ := eclat_unit;
              \$v6439\ := \$code_lock\;
              if \$v6439\(0) = '1' then
                state_var7462 := Q_WAIT6438;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 8;\$code_write\ <= "000"& X"000000" & X"1"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6437;
              end if;
            when PAUSE_SET6443 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12693\ := eclat_unit;
              \$v6442\ := \$code_lock\;
              if \$v6442\(0) = '1' then
                state_var7462 := Q_WAIT6441;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 7;\$code_write\ <= "000"& X"00000" & X"28"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6440;
              end if;
            when PAUSE_SET6446 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12692\ := eclat_unit;
              \$v6445\ := \$code_lock\;
              if \$v6445\(0) = '1' then
                state_var7462 := Q_WAIT6444;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 6;\$code_write\ <= "000"& X"00000" & X"64"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6443;
              end if;
            when PAUSE_SET6449 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12691\ := eclat_unit;
              \$v6448\ := \$code_lock\;
              if \$v6448\(0) = '1' then
                state_var7462 := Q_WAIT6447;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 5;\$code_write\ <= "000"& X"000000" & X"4"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6446;
              end if;
            when PAUSE_SET6452 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12690\ := eclat_unit;
              \$v6451\ := \$code_lock\;
              if \$v6451\(0) = '1' then
                state_var7462 := Q_WAIT6450;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 4;\$code_write\ <= "000"& X"000000" & X"2"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6449;
              end if;
            when PAUSE_SET6455 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12689\ := eclat_unit;
              \$v6454\ := \$code_lock\;
              if \$v6454\(0) = '1' then
                state_var7462 := Q_WAIT6453;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 3;\$code_write\ <= "000"& X"00000" & X"86"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6452;
              end if;
            when PAUSE_SET6458 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12688\ := eclat_unit;
              \$v6457\ := \$code_lock\;
              if \$v6457\(0) = '1' then
                state_var7462 := Q_WAIT6456;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 2;\$code_write\ <= "000"& X"000000" & X"0"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6455;
              end if;
            when PAUSE_SET6461 =>
              \$code_write_request\ <= '0';
              release(\$code_lock\);
              \$12687\ := eclat_unit;
              \$v6460\ := \$code_lock\;
              if \$v6460\(0) = '1' then
                state_var7462 := Q_WAIT6459;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 1;\$code_write\ <= "000"& X"00000" & X"15"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6458;
              end if;
            when PAUSE_SET6464 =>
              \$global_end_write_request\ <= '0';
              release(\$global_end_lock\);
              \$12685\ := eclat_unit;
              \$v6463\ := \$code_lock\;
              if \$v6463\(0) = '1' then
                state_var7462 := Q_WAIT6462;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 0;\$code_write\ <= "000"& X"00000" & X"54"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6461;
              end if;
            when Q_WAIT6116 =>
              \$v6117\ := \$ram_lock\;
              if \$v6117\(0) = '1' then
                state_var7462 := Q_WAIT6116;
              else
                acquire(\$ram_lock\);
                \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                        \$12679_loop666_arg\(16 to 31), \$12679_loop666_arg\(0 to 15))));
                \$ram_write\ <= \$13889\; \$ram_write_request\ <= '1';
                state_var7462 := PAUSE_SET6115;
              end if;
            when Q_WAIT6119 =>
              \$v6120\ := \$ram_lock\;
              if \$v6120\(0) = '1' then
                state_var7462 := Q_WAIT6119;
              else
                acquire(\$ram_lock\);
                \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$12679_loop666_arg\(32 to 47), \$12679_loop666_arg\(0 to 15))));
                state_var7462 := PAUSE_GET6118;
              end if;
            when Q_WAIT6123 =>
              \$v6124\ := \$ram_lock\;
              if \$v6124\(0) = '1' then
                state_var7462 := Q_WAIT6123;
              else
                acquire(\$ram_lock\);
                \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                        \$12680_loop665_arg\(64 to 79), \$12680_loop665_arg\(0 to 15))));
                \$ram_write\ <= \$13791\(0 to 31); \$ram_write_request\ <= '1';
                state_var7462 := PAUSE_SET6122;
              end if;
            when Q_WAIT6126 =>
              \$v6127\ := \$ram_lock\;
              if \$v6127\(0) = '1' then
                state_var7462 := Q_WAIT6126;
              else
                acquire(\$ram_lock\);
                \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                        eclat_resize(\$13787\(0 to 30),16), X"000" & X"1")));
                \$ram_write\ <= eclat_resize(\$12680_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                state_var7462 := PAUSE_SET6125;
              end if;
            when Q_WAIT6129 =>
              \$v6130\ := \$ram_lock\;
              if \$v6130\(0) = '1' then
                state_var7462 := Q_WAIT6129;
              else
                acquire(\$ram_lock\);
                \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$13787\(0 to 30),16)));
                \$ram_write\ <= eclat_resize(\$12680_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                state_var7462 := PAUSE_SET6128;
              end if;
            when Q_WAIT6132 =>
              \$v6133\ := \$ram_lock\;
              if \$v6133\(0) = '1' then
                state_var7462 := Q_WAIT6132;
              else
                acquire(\$ram_lock\);
                \$ram_ptr_write\ <= to_integer(unsigned(\$12680_loop665_arg\(16 to 31)));
                \$ram_write\ <= \$13808_hd\; \$ram_write_request\ <= '1';
                state_var7462 := PAUSE_SET6131;
              end if;
            when Q_WAIT6135 =>
              \$v6136\ := \$ram_lock\;
              if \$v6136\(0) = '1' then
                state_var7462 := Q_WAIT6135;
              else
                acquire(\$ram_lock\);
                \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$13787\(0 to 30),16)));
                state_var7462 := PAUSE_GET6134;
              end if;
            when Q_WAIT6139 =>
              \$v6140\ := \$ram_lock\;
              if \$v6140\(0) = '1' then
                state_var7462 := Q_WAIT6139;
              else
                acquire(\$ram_lock\);
                \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$13787\(0 to 30),16), X"000" & X"1")));
                state_var7462 := PAUSE_GET6138;
              end if;
            when Q_WAIT6143 =>
              \$v6144\ := \$ram_lock\;
              if \$v6144\(0) = '1' then
                state_var7462 := Q_WAIT6143;
              else
                acquire(\$ram_lock\);
                \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$12680_loop665_arg\(64 to 79), \$12680_loop665_arg\(0 to 15))));
                state_var7462 := PAUSE_GET6142;
              end if;
            when Q_WAIT6357 =>
              \$v6358\ := \$ram_lock\;
              if \$v6358\(0) = '1' then
                state_var7462 := Q_WAIT6357;
              else
                acquire(\$ram_lock\);
                \$ram_ptr_write\ <= to_integer(unsigned(\$12737\(64 to 79)));
                \$ram_write\ <= work.Int.lor(work.Int.lsl(eclat_resize(\$12682_make_block579_arg\(80 to 111),31), X"000000" & X"18"), 
                                             work.Int.lsl(eclat_resize(
                                                          eclat_if(work.Int.eq(
                                                                   \$12682_make_block579_arg\(112 to 127), X"000" & X"0") & X"000" & X"1" & \$12682_make_block579_arg\(112 to 127)),31), X"0000000" & X"2")) & eclat_true; \$ram_write_request\ <= '1';
                state_var7462 := PAUSE_SET6356;
              end if;
            when Q_WAIT6360 =>
              \$v6361\ := \$code_lock\;
              if \$v6361\(0) = '1' then
                state_var7462 := Q_WAIT6360;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 34;\$code_write\ <= "000"& X"00000" & X"8f"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6359;
              end if;
            when Q_WAIT6363 =>
              \$v6364\ := \$code_lock\;
              if \$v6364\(0) = '1' then
                state_var7462 := Q_WAIT6363;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 33;\$code_write\ <= "000"& X"000000" & X"1"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6362;
              end if;
            when Q_WAIT6366 =>
              \$v6367\ := \$code_lock\;
              if \$v6367\(0) = '1' then
                state_var7462 := Q_WAIT6366;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 32;\$code_write\ <= "000"& X"00000" & X"13"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6365;
              end if;
            when Q_WAIT6369 =>
              \$v6370\ := \$code_lock\;
              if \$v6370\(0) = '1' then
                state_var7462 := Q_WAIT6369;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 31;\$code_write\ <= "000"& X"000000" & X"0"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6368;
              end if;
            when Q_WAIT6372 =>
              \$v6373\ := \$code_lock\;
              if \$v6373\(0) = '1' then
                state_var7462 := Q_WAIT6372;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 30;\$code_write\ <= "000"& X"00000" & X"5d"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6371;
              end if;
            when Q_WAIT6375 =>
              \$v6376\ := \$code_lock\;
              if \$v6376\(0) = '1' then
                state_var7462 := Q_WAIT6375;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 29;\$code_write\ <= "000"& X"00000" & X"21"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6374;
              end if;
            when Q_WAIT6378 =>
              \$v6379\ := \$code_lock\;
              if \$v6379\(0) = '1' then
                state_var7462 := Q_WAIT6378;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 28;\$code_write\ <= "000"& X"000000" & X"b"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6377;
              end if;
            when Q_WAIT6381 =>
              \$v6382\ := \$code_lock\;
              if \$v6382\(0) = '1' then
                state_var7462 := Q_WAIT6381;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 27;\$code_write\ <= "000"& X"000000" & X"b"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6380;
              end if;
            when Q_WAIT6384 =>
              \$v6385\ := \$code_lock\;
              if \$v6385\(0) = '1' then
                state_var7462 := Q_WAIT6384;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 26;\$code_write\ <= "000"& X"00000" & X"67"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6383;
              end if;
            when Q_WAIT6387 =>
              \$v6388\ := \$code_lock\;
              if \$v6388\(0) = '1' then
                state_var7462 := Q_WAIT6387;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 25;\$code_write\ <= work.Int.neg(
                                                         "000"& X"00000" & X"17"); \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6386;
              end if;
            when Q_WAIT6390 =>
              \$v6391\ := \$code_lock\;
              if \$v6391\(0) = '1' then
                state_var7462 := Q_WAIT6390;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 24;\$code_write\ <= "000"& X"000000" & X"0"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6389;
              end if;
            when Q_WAIT6393 =>
              \$v6394\ := \$code_lock\;
              if \$v6394\(0) = '1' then
                state_var7462 := Q_WAIT6393;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 23;\$code_write\ <= "000"& X"000000" & X"1"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6392;
              end if;
            when Q_WAIT6396 =>
              \$v6397\ := \$code_lock\;
              if \$v6397\(0) = '1' then
                state_var7462 := Q_WAIT6396;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 22;\$code_write\ <= "000"& X"00000" & X"2c"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6395;
              end if;
            when Q_WAIT6399 =>
              \$v6400\ := \$code_lock\;
              if \$v6400\(0) = '1' then
                state_var7462 := Q_WAIT6399;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 21;\$code_write\ <= "000"& X"000000" & X"1"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6398;
              end if;
            when Q_WAIT6402 =>
              \$v6403\ := \$code_lock\;
              if \$v6403\(0) = '1' then
                state_var7462 := Q_WAIT6402;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 20;\$code_write\ <= "000"& X"00000" & X"28"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6401;
              end if;
            when Q_WAIT6405 =>
              \$v6406\ := \$code_lock\;
              if \$v6406\(0) = '1' then
                state_var7462 := Q_WAIT6405;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 19;\$code_write\ <= "000"& X"00000" & X"6e"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6404;
              end if;
            when Q_WAIT6408 =>
              \$v6409\ := \$code_lock\;
              if \$v6409\(0) = '1' then
                state_var7462 := Q_WAIT6408;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 18;\$code_write\ <= "000"& X"00000" & X"21"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6407;
              end if;
            when Q_WAIT6411 =>
              \$v6412\ := \$code_lock\;
              if \$v6412\(0) = '1' then
                state_var7462 := Q_WAIT6411;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 17;\$code_write\ <= "000"& X"00000" & X"32"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6410;
              end if;
            when Q_WAIT6414 =>
              \$v6415\ := \$code_lock\;
              if \$v6415\(0) = '1' then
                state_var7462 := Q_WAIT6414;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 16;\$code_write\ <= work.Int.neg(
                                                         "000"& X"000000" & X"1"); \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6413;
              end if;
            when Q_WAIT6417 =>
              \$v6418\ := \$code_lock\;
              if \$v6418\(0) = '1' then
                state_var7462 := Q_WAIT6417;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 15;\$code_write\ <= "000"& X"00000" & X"7f"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6416;
              end if;
            when Q_WAIT6420 =>
              \$v6421\ := \$code_lock\;
              if \$v6421\(0) = '1' then
                state_var7462 := Q_WAIT6420;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 14;\$code_write\ <= "000"& X"000000" & X"b"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6419;
              end if;
            when Q_WAIT6423 =>
              \$v6424\ := \$code_lock\;
              if \$v6424\(0) = '1' then
                state_var7462 := Q_WAIT6423;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 13;\$code_write\ <= "000"& X"00000" & X"21"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6422;
              end if;
            when Q_WAIT6426 =>
              \$v6427\ := \$code_lock\;
              if \$v6427\(0) = '1' then
                state_var7462 := Q_WAIT6426;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 12;\$code_write\ <= "000"& X"00000" & X"32"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6425;
              end if;
            when Q_WAIT6429 =>
              \$v6430\ := \$code_lock\;
              if \$v6430\(0) = '1' then
                state_var7462 := Q_WAIT6429;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 11;\$code_write\ <= work.Int.neg(
                                                         "000"& X"000000" & X"2"); \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6428;
              end if;
            when Q_WAIT6432 =>
              \$v6433\ := \$code_lock\;
              if \$v6433\(0) = '1' then
                state_var7462 := Q_WAIT6432;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 10;\$code_write\ <= "000"& X"00000" & X"7f"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6431;
              end if;
            when Q_WAIT6435 =>
              \$v6436\ := \$code_lock\;
              if \$v6436\(0) = '1' then
                state_var7462 := Q_WAIT6435;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 9;\$code_write\ <= "000"& X"000000" & X"0"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6434;
              end if;
            when Q_WAIT6438 =>
              \$v6439\ := \$code_lock\;
              if \$v6439\(0) = '1' then
                state_var7462 := Q_WAIT6438;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 8;\$code_write\ <= "000"& X"000000" & X"1"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6437;
              end if;
            when Q_WAIT6441 =>
              \$v6442\ := \$code_lock\;
              if \$v6442\(0) = '1' then
                state_var7462 := Q_WAIT6441;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 7;\$code_write\ <= "000"& X"00000" & X"28"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6440;
              end if;
            when Q_WAIT6444 =>
              \$v6445\ := \$code_lock\;
              if \$v6445\(0) = '1' then
                state_var7462 := Q_WAIT6444;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 6;\$code_write\ <= "000"& X"00000" & X"64"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6443;
              end if;
            when Q_WAIT6447 =>
              \$v6448\ := \$code_lock\;
              if \$v6448\(0) = '1' then
                state_var7462 := Q_WAIT6447;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 5;\$code_write\ <= "000"& X"000000" & X"4"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6446;
              end if;
            when Q_WAIT6450 =>
              \$v6451\ := \$code_lock\;
              if \$v6451\(0) = '1' then
                state_var7462 := Q_WAIT6450;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 4;\$code_write\ <= "000"& X"000000" & X"2"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6449;
              end if;
            when Q_WAIT6453 =>
              \$v6454\ := \$code_lock\;
              if \$v6454\(0) = '1' then
                state_var7462 := Q_WAIT6453;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 3;\$code_write\ <= "000"& X"00000" & X"86"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6452;
              end if;
            when Q_WAIT6456 =>
              \$v6457\ := \$code_lock\;
              if \$v6457\(0) = '1' then
                state_var7462 := Q_WAIT6456;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 2;\$code_write\ <= "000"& X"000000" & X"0"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6455;
              end if;
            when Q_WAIT6459 =>
              \$v6460\ := \$code_lock\;
              if \$v6460\(0) = '1' then
                state_var7462 := Q_WAIT6459;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 1;\$code_write\ <= "000"& X"00000" & X"15"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6458;
              end if;
            when Q_WAIT6462 =>
              \$v6463\ := \$code_lock\;
              if \$v6463\(0) = '1' then
                state_var7462 := Q_WAIT6462;
              else
                acquire(\$code_lock\);
                \$code_ptr_write\ <= 0;\$code_write\ <= "000"& X"00000" & X"54"; \$code_write_request\ <= '1';
                state_var7462 := PAUSE_SET6461;
              end if;
            when Q_WAIT6465 =>
              \$v6466\ := \$global_end_lock\;
              if \$v6466\(0) = '1' then
                state_var7462 := Q_WAIT6465;
              else
                acquire(\$global_end_lock\);
                \$global_end_ptr_write\ <= 0;\$global_end_write\ <= work.Int.add(
                                                                    X"3e80", X"000" & X"c"); \$global_end_write_request\ <= '1';
                state_var7462 := PAUSE_SET6464;
              end if;
            when IDLE6114 =>
              rdy6113 := eclat_false;
              \$v6466\ := \$global_end_lock\;
              if \$v6466\(0) = '1' then
                state_var7462 := Q_WAIT6465;
              else
                acquire(\$global_end_lock\);
                \$global_end_ptr_write\ <= 0;\$global_end_write\ <= work.Int.add(
                                                                    X"3e80", X"000" & X"c"); \$global_end_write_request\ <= '1';
                state_var7462 := PAUSE_SET6464;
              end if;
            end case;
            
            if rdy6113(0) = '1' then
              
            else
              result6112 := eclat_unit;
            end if;
            \$12670\ := result6112 & rdy6113;
            if \$v5871\(0) = '1' then
              
            else
              \$v5871\ := eclat_true;
              \$12674\ := eclat_false;
            end if;
            \$12674\ := work.Bool.land(eclat_if(\$12674\ & eclat_true & ""&\$12670\(1)), 
                                       work.Bool.lnot(eclat_false));
            \$12673_rdy\ := \$12674\;
            \$12662\ := eclat_false & eclat_true & \$12673_rdy\ & ""&\$12662\(3);
          else
            if \$v5872\(0) = '1' then
              
            else
              \$v5872\ := eclat_true;
              \$13911\ := X"000" & X"0" & "000"& X"000000" & X"1" & eclat_true & X"0" & X"3e8" & "000"& X"000000" & X"1" & eclat_true & "00000000" & X"000" & X"0" & eclat_false & eclat_false & eclat_true;
            end if;
            \$v7457\ := work.Bool.lnot(""&\$12662\(2));
            if \$v7457\(0) = '1' then
              \$13911\ := \$13911\(0 to 121) & eclat_true;
            else
              case state_var7460 is
              when \$13920_LOOP666\ =>
                \$v6477\ := work.Int.ge(\$13920_loop666_arg\(0 to 15), 
                                        work.Int.add(\$13920_loop666_arg\(48 to 63), X"000" & X"1"));
                if \$v6477\(0) = '1' then
                  \$13920_loop666_result\ := eclat_unit;
                  \$18478\ := \$13920_loop666_result\;
                  \$v6486\ := \$ram_lock\;
                  if \$v6486\(0) = '1' then
                    state_var7460 := Q_WAIT6485;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18443\(0 to 30),16)));
                    \$ram_write\ <= eclat_resize(\$13921_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET6484;
                  end if;
                else
                  \$v6476\ := \$ram_lock\;
                  if \$v6476\(0) = '1' then
                    state_var7460 := Q_WAIT6475;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$13920_loop666_arg\(32 to 47), \$13920_loop666_arg\(0 to 15))));
                    state_var7460 := PAUSE_GET6474;
                  end if;
                end if;
              when \$13921_LOOP665\ =>
                \$v6501\ := work.Int.ge(\$13921_loop665_arg\(0 to 15), 
                                        work.Int.add(\$13921_loop665_arg\(80 to 95), X"000" & X"1"));
                if \$v6501\(0) = '1' then
                  \$13921_loop665_result\ := \$13921_loop665_arg\(16 to 31);
                  state_var7460 := \$13921_LOOP665\;
                else
                  \$v6500\ := \$ram_lock\;
                  if \$v6500\(0) = '1' then
                    state_var7460 := Q_WAIT6499;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$13921_loop665_arg\(64 to 79), \$13921_loop665_arg\(0 to 15))));
                    state_var7460 := PAUSE_GET6498;
                  end if;
                end if;
              when \$13922_WAIT662\ =>
                if \$v5874\(0) = '1' then
                  
                else
                  \$v5874\ := eclat_true;
                  \$17444\ := \$13922_wait662_arg\(1 to 32) & \$13922_wait662_arg\(33 to 64) & X"0" & X"fa0" & X"0" & X"fa0" & X"0" & X"fa0" & 
                  work.Int.add(X"0" & X"fa0", X"1770") & eclat_false;
                end if;
                case state_var7461 is
                when \$17455_LOOP666\ =>
                  \$v6512\ := work.Int.ge(\$17455_loop666_arg\(0 to 15), 
                                          work.Int.add(\$17455_loop666_arg\(48 to 63), X"000" & X"1"));
                  if \$v6512\(0) = '1' then
                    \$17455_loop666_result\ := eclat_unit;
                    \$18354\ := \$17455_loop666_result\;
                    \$v6521\ := \$ram_lock\;
                    if \$v6521\(0) = '1' then
                      state_var7461 := Q_WAIT6520;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18319\(0 to 30),16)));
                      \$ram_write\ <= eclat_resize(\$17456_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                      state_var7461 := PAUSE_SET6519;
                    end if;
                  else
                    \$v6511\ := \$ram_lock\;
                    if \$v6511\(0) = '1' then
                      state_var7461 := Q_WAIT6510;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                        \$17455_loop666_arg\(32 to 47), \$17455_loop666_arg\(0 to 15))));
                      state_var7461 := PAUSE_GET6509;
                    end if;
                  end if;
                when \$17456_LOOP665\ =>
                  \$v6536\ := work.Int.ge(\$17456_loop665_arg\(0 to 15), 
                                          work.Int.add(\$17456_loop665_arg\(80 to 95), X"000" & X"1"));
                  if \$v6536\(0) = '1' then
                    \$17456_loop665_result\ := \$17456_loop665_arg\(16 to 31);
                    \$18288_next\ := \$17456_loop665_result\;
                    \$17457_aux664_arg\ := work.Int.add(\$17457_aux664_arg\(0 to 15), 
                                                        work.Int.add(
                                                        eclat_resize(
                                                        work.Int.lsr(
                                                        eclat_resize(eclat_resize(\$18284\(0 to 30),16),31), X"0000000" & X"2"),16), X"000" & X"1")) & \$18288_next\ & \$17457_aux664_arg\(32 to 47) & \$17457_aux664_arg\(48 to 63);
                    state_var7461 := \$17457_AUX664\;
                  else
                    \$v6535\ := \$ram_lock\;
                    if \$v6535\(0) = '1' then
                      state_var7461 := Q_WAIT6534;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                        \$17456_loop665_arg\(64 to 79), \$17456_loop665_arg\(0 to 15))));
                      state_var7461 := PAUSE_GET6533;
                    end if;
                  end if;
                when \$17457_AUX664\ =>
                  \$18278\ := work.Print.print_string(clk,of_string("     scan="));
                  \$18279\ := work.Int.print(clk,\$17457_aux664_arg\(0 to 15));
                  \$18280\ := work.Print.print_string(clk,of_string(" | next="));
                  \$18281\ := work.Int.print(clk,\$17457_aux664_arg\(16 to 31));
                  \$18282\ := work.Print.print_newline(clk,eclat_unit);
                  \$v6540\ := work.Int.ge(\$17457_aux664_arg\(0 to 15), \$17457_aux664_arg\(16 to 31));
                  if \$v6540\(0) = '1' then
                    \$17457_aux664_result\ := \$17457_aux664_arg\(16 to 31);
                    state_var7461 := \$17457_AUX664\;
                  else
                    \$v6539\ := \$ram_lock\;
                    if \$v6539\(0) = '1' then
                      state_var7461 := Q_WAIT6538;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(\$17457_aux664_arg\(0 to 15)));
                      state_var7461 := PAUSE_GET6537;
                    end if;
                  end if;
                when \$17458_LOOP666\ =>
                  \$v6547\ := work.Int.ge(\$17458_loop666_arg\(0 to 15), 
                                          work.Int.add(\$17458_loop666_arg\(48 to 63), X"000" & X"1"));
                  if \$v6547\(0) = '1' then
                    \$17458_loop666_result\ := eclat_unit;
                    case \$17458_loop666_id\ is
                    when "000000100011" =>
                      \$18194\ := \$17458_loop666_result\;
                      \$v6556\ := \$ram_lock\;
                      if \$v6556\(0) = '1' then
                        state_var7461 := Q_WAIT6555;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18159\(0 to 30),16)));
                        \$ram_write\ <= eclat_resize(\$17459_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                        state_var7461 := PAUSE_SET6554;
                      end if;
                    when "000000101001" =>
                      \$17599\ := \$17458_loop666_result\;
                      \$v6585\ := \$ram_lock\;
                      if \$v6585\(0) = '1' then
                        state_var7461 := Q_WAIT6584;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$17562\(0 to 30),16)));
                        \$ram_write\ <= eclat_resize(\$17547_copy_root_in_ram6635891_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                        state_var7461 := PAUSE_SET6583;
                      end if;
                    when "000000101011" =>
                      \$17679\ := \$17458_loop666_result\;
                      \$v6609\ := \$ram_lock\;
                      if \$v6609\(0) = '1' then
                        state_var7461 := Q_WAIT6608;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$17535\(0 to 30),16)));
                        \$ram_write\ <= eclat_resize(\$17520_copy_root_in_ram6635893_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                        state_var7461 := PAUSE_SET6607;
                      end if;
                    when "000000101101" =>
                      \$17813\ := \$17458_loop666_result\;
                      \$v6636\ := \$ram_lock\;
                      if \$v6636\(0) = '1' then
                        state_var7461 := Q_WAIT6635;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$17776\(0 to 30),16)));
                        \$ram_write\ <= eclat_resize(\$17761_copy_root_in_ram6635891_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                        state_var7461 := PAUSE_SET6634;
                      end if;
                    when "000000101111" =>
                      \$17893\ := \$17458_loop666_result\;
                      \$v6660\ := \$ram_lock\;
                      if \$v6660\(0) = '1' then
                        state_var7461 := Q_WAIT6659;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$17749\(0 to 30),16)));
                        \$ram_write\ <= eclat_resize(\$17734_copy_root_in_ram6635892_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                        state_var7461 := PAUSE_SET6658;
                      end if;
                    when "000000110001" =>
                      \$17971\ := \$17458_loop666_result\;
                      \$v6681\ := \$ram_lock\;
                      if \$v6681\(0) = '1' then
                        state_var7461 := Q_WAIT6680;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$13922_wait662_arg\(33 to 63),16)));
                        \$ram_write\ <= eclat_resize(\$17470\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                        state_var7461 := PAUSE_SET6679;
                      end if;
                    when "000000110010" =>
                      \$18049\ := \$17458_loop666_result\;
                      \$v6698\ := \$ram_lock\;
                      if \$v6698\(0) = '1' then
                        state_var7461 := Q_WAIT6697;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$13922_wait662_arg\(1 to 31),16)));
                        \$ram_write\ <= eclat_resize(\$17444\(112 to 127),31) & eclat_false; \$ram_write_request\ <= '1';
                        state_var7461 := PAUSE_SET6696;
                      end if;
                    when others =>
                      
                    end case;
                  else
                    \$v6546\ := \$ram_lock\;
                    if \$v6546\(0) = '1' then
                      state_var7461 := Q_WAIT6545;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                        \$17458_loop666_arg\(32 to 47), \$17458_loop666_arg\(0 to 15))));
                      state_var7461 := PAUSE_GET6544;
                    end if;
                  end if;
                when \$17459_LOOP665\ =>
                  \$v6571\ := work.Int.ge(\$17459_loop665_arg\(0 to 15), 
                                          work.Int.add(\$17459_loop665_arg\(80 to 95), X"000" & X"1"));
                  if \$v6571\(0) = '1' then
                    \$17459_loop665_result\ := \$17459_loop665_arg\(16 to 31);
                    \$18128_next\ := \$17459_loop665_result\;
                    \$17460_aux664_arg\ := work.Int.add(\$17460_aux664_arg\(0 to 15), 
                                                        work.Int.add(
                                                        eclat_resize(
                                                        work.Int.lsr(
                                                        eclat_resize(eclat_resize(\$18124\(0 to 30),16),31), X"0000000" & X"2"),16), X"000" & X"1")) & \$18128_next\ & \$17460_aux664_arg\(32 to 47) & \$17460_aux664_arg\(48 to 63);
                    state_var7461 := \$17460_AUX664\;
                  else
                    \$v6570\ := \$ram_lock\;
                    if \$v6570\(0) = '1' then
                      state_var7461 := Q_WAIT6569;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                        \$17459_loop665_arg\(64 to 79), \$17459_loop665_arg\(0 to 15))));
                      state_var7461 := PAUSE_GET6568;
                    end if;
                  end if;
                when \$17460_AUX664\ =>
                  \$18118\ := work.Print.print_string(clk,of_string("     scan="));
                  \$18119\ := work.Int.print(clk,\$17460_aux664_arg\(0 to 15));
                  \$18120\ := work.Print.print_string(clk,of_string(" | next="));
                  \$18121\ := work.Int.print(clk,\$17460_aux664_arg\(16 to 31));
                  \$18122\ := work.Print.print_newline(clk,eclat_unit);
                  \$v6575\ := work.Int.ge(\$17460_aux664_arg\(0 to 15), \$17460_aux664_arg\(16 to 31));
                  if \$v6575\(0) = '1' then
                    \$17460_aux664_result\ := \$17460_aux664_arg\(16 to 31);
                    \$17496_next\ := \$17460_aux664_result\;
                    \$17497\ := work.Print.print_string(clk,of_string("memory copied in to_space : "));
                    \$17498\ := work.Int.print(clk,work.Int.sub(\$17496_next\, \$17444\(112 to 127)));
                    \$17499\ := work.Print.print_string(clk,of_string(" words"));
                    \$17500\ := work.Print.print_newline(clk,eclat_unit);
                    \$v6576\ := work.Int.gt(work.Int.sub(\$17496_next\, \$17444\(112 to 127)), X"1770");
                    if \$v6576\(0) = '1' then
                      \$17502\ := work.Print.print_string(clk,of_string("fatal error: "));
                      \$17503\ := work.Print.print_string(clk,of_string("Out of memory"));
                      \$17504\ := work.Print.print_newline(clk,eclat_unit);
                      \$17505_forever6705894_id\ := "000000100111";
                      \$17505_forever6705894_arg\ := eclat_unit;
                      state_var7461 := \$17505_FOREVER6705894\;
                    else
                      \$17476\ := \$17470\(0 to 31) & \$17487\(0 to 31) & \$17496_next\;
                      \$17481\ := work.Print.print_newline(clk,eclat_unit);
                      \$17482\ := work.Print.print_newline(clk,eclat_unit);
                      \$17483\ := work.Print.print_string(clk,of_string("[================= GC END ======================]"));
                      \$17486\ := work.Print.print_newline(clk,eclat_unit);
                      \$17484\ := work.Print.print_newline(clk,eclat_unit);
                      result6503 := \$17476\(0 to 31) & \$17476\(32 to 63) & \$17476\(64 to 79) & 
                      work.Int.add(\$17476\(64 to 79), \$13922_wait662_arg\(81 to 96)) & \$17444\(112 to 127) & \$17444\(96 to 111);
                      rdy6504 := eclat_true;
                      state_var7461 := IDLE6505;
                    end if;
                  else
                    \$v6574\ := \$ram_lock\;
                    if \$v6574\(0) = '1' then
                      state_var7461 := Q_WAIT6573;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(\$17460_aux664_arg\(0 to 15)));
                      state_var7461 := PAUSE_GET6572;
                    end if;
                  end if;
                when \$17505_FOREVER6705894\ =>
                  \$17509_forever6705890_id\ := "000000100110";
                  \$17509_forever6705890_arg\ := eclat_unit;
                  state_var7461 := \$17509_FOREVER6705890\;
                when \$17509_FOREVER6705890\ =>
                  \$17513_forever6705889_id\ := "000000100101";
                  \$17513_forever6705889_arg\ := eclat_unit;
                  state_var7461 := \$17513_FOREVER6705889\;
                when \$17513_FOREVER6705889\ =>
                  \$17513_forever6705889_arg\ := eclat_unit;
                  state_var7461 := \$17513_FOREVER6705889\;
                when \$17520_COPY_ROOT_IN_RAM6635893\ =>
                  \$v6624\ := work.Int.ge(\$17520_copy_root_in_ram6635893_arg\(0 to 15), \$17520_copy_root_in_ram6635893_arg\(16 to 31));
                  if \$v6624\(0) = '1' then
                    \$17520_copy_root_in_ram6635893_result\ := \$17520_copy_root_in_ram6635893_arg\(32 to 47);
                    \$17492_next\ := \$17520_copy_root_in_ram6635893_result\;
                    \$17494\ := work.Print.print_string(clk,of_string("======================================="));
                    \$17495\ := work.Print.print_newline(clk,eclat_unit);
                    \$17460_aux664_id\ := "000000101000";
                    \$17460_aux664_arg\ := \$17444\(112 to 127) & \$17492_next\ & \$17444\(96 to 111) & \$17444\(112 to 127);
                    state_var7461 := \$17460_AUX664\;
                  else
                    \$17532\ := work.Print.print_string(clk,of_string("racine:"));
                    \$17533\ := work.Int.print(clk,\$17520_copy_root_in_ram6635893_arg\(0 to 15));
                    \$17534\ := work.Print.print_newline(clk,eclat_unit);
                    \$v6623\ := \$ram_lock\;
                    if \$v6623\(0) = '1' then
                      state_var7461 := Q_WAIT6622;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(\$17520_copy_root_in_ram6635893_arg\(0 to 15)));
                      state_var7461 := PAUSE_GET6621;
                    end if;
                  end if;
                when \$17547_COPY_ROOT_IN_RAM6635891\ =>
                  \$v6600\ := work.Int.ge(\$17547_copy_root_in_ram6635891_arg\(0 to 15), \$17547_copy_root_in_ram6635891_arg\(16 to 31));
                  if \$v6600\(0) = '1' then
                    \$17547_copy_root_in_ram6635891_result\ := \$17547_copy_root_in_ram6635891_arg\(32 to 47);
                    \$17520_copy_root_in_ram6635893_result\ := \$17547_copy_root_in_ram6635891_result\;
                    \$17492_next\ := \$17520_copy_root_in_ram6635893_result\;
                    \$17494\ := work.Print.print_string(clk,of_string("======================================="));
                    \$17495\ := work.Print.print_newline(clk,eclat_unit);
                    \$17460_aux664_id\ := "000000101000";
                    \$17460_aux664_arg\ := \$17444\(112 to 127) & \$17492_next\ & \$17444\(96 to 111) & \$17444\(112 to 127);
                    state_var7461 := \$17460_AUX664\;
                  else
                    \$17559\ := work.Print.print_string(clk,of_string("racine:"));
                    \$17560\ := work.Int.print(clk,\$17547_copy_root_in_ram6635891_arg\(0 to 15));
                    \$17561\ := work.Print.print_newline(clk,eclat_unit);
                    \$v6599\ := \$ram_lock\;
                    if \$v6599\(0) = '1' then
                      state_var7461 := Q_WAIT6598;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(\$17547_copy_root_in_ram6635891_arg\(0 to 15)));
                      state_var7461 := PAUSE_GET6597;
                    end if;
                  end if;
                when \$17734_COPY_ROOT_IN_RAM6635892\ =>
                  \$v6675\ := work.Int.ge(\$17734_copy_root_in_ram6635892_arg\(0 to 15), \$17734_copy_root_in_ram6635892_arg\(16 to 31));
                  if \$v6675\(0) = '1' then
                    \$17734_copy_root_in_ram6635892_result\ := \$17734_copy_root_in_ram6635892_arg\(32 to 47);
                    \$17490_next\ := \$17734_copy_root_in_ram6635892_result\;
                    \$v6627\ := \$global_end_lock\;
                    if \$v6627\(0) = '1' then
                      state_var7461 := Q_WAIT6626;
                    else
                      acquire(\$global_end_lock\);
                      \$global_end_ptr\ <= 0;
                      state_var7461 := PAUSE_GET6625;
                    end if;
                  else
                    \$17746\ := work.Print.print_string(clk,of_string("racine:"));
                    \$17747\ := work.Int.print(clk,\$17734_copy_root_in_ram6635892_arg\(0 to 15));
                    \$17748\ := work.Print.print_newline(clk,eclat_unit);
                    \$v6674\ := \$ram_lock\;
                    if \$v6674\(0) = '1' then
                      state_var7461 := Q_WAIT6673;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(\$17734_copy_root_in_ram6635892_arg\(0 to 15)));
                      state_var7461 := PAUSE_GET6672;
                    end if;
                  end if;
                when \$17761_COPY_ROOT_IN_RAM6635891\ =>
                  \$v6651\ := work.Int.ge(\$17761_copy_root_in_ram6635891_arg\(0 to 15), \$17761_copy_root_in_ram6635891_arg\(16 to 31));
                  if \$v6651\(0) = '1' then
                    \$17761_copy_root_in_ram6635891_result\ := \$17761_copy_root_in_ram6635891_arg\(32 to 47);
                    \$17734_copy_root_in_ram6635892_result\ := \$17761_copy_root_in_ram6635891_result\;
                    \$17490_next\ := \$17734_copy_root_in_ram6635892_result\;
                    \$v6627\ := \$global_end_lock\;
                    if \$v6627\(0) = '1' then
                      state_var7461 := Q_WAIT6626;
                    else
                      acquire(\$global_end_lock\);
                      \$global_end_ptr\ <= 0;
                      state_var7461 := PAUSE_GET6625;
                    end if;
                  else
                    \$17773\ := work.Print.print_string(clk,of_string("racine:"));
                    \$17774\ := work.Int.print(clk,\$17761_copy_root_in_ram6635891_arg\(0 to 15));
                    \$17775\ := work.Print.print_newline(clk,eclat_unit);
                    \$v6650\ := \$ram_lock\;
                    if \$v6650\(0) = '1' then
                      state_var7461 := Q_WAIT6649;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(\$17761_copy_root_in_ram6635891_arg\(0 to 15)));
                      state_var7461 := PAUSE_GET6648;
                    end if;
                  end if;
                when PAUSE_GET6509 =>
                  \$18421\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v6508\ := \$ram_lock\;
                  if \$v6508\(0) = '1' then
                    state_var7461 := Q_WAIT6507;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            \$17455_loop666_arg\(16 to 31), \$17455_loop666_arg\(0 to 15))));
                    \$ram_write\ <= \$18421\; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6506;
                  end if;
                when PAUSE_GET6525 =>
                  \$18340_hd\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$18344\ := work.Print.print_string(clk,of_string("bloc "));
                  \$18345\ := work.Int.print(clk,eclat_resize(\$18319\(0 to 30),16));
                  \$18346\ := work.Print.print_string(clk,of_string(" of size "));
                  \$18347\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                              work.Int.lsr(
                                                              \$18340_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$18348\ := work.Print.print_string(clk,of_string(" from "));
                  \$18349\ := work.Int.print(clk,eclat_resize(\$18319\(0 to 30),16));
                  \$18350\ := work.Print.print_string(clk,of_string(" to "));
                  \$18351\ := work.Int.print(clk,\$17456_loop665_arg\(16 to 31));
                  \$18352\ := work.Print.print_newline(clk,eclat_unit);
                  \$v6524\ := \$ram_lock\;
                  if \$v6524\(0) = '1' then
                    state_var7461 := Q_WAIT6523;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17456_loop665_arg\(16 to 31)));
                    \$ram_write\ <= \$18340_hd\; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6522;
                  end if;
                when PAUSE_GET6529 =>
                  \$18335_w\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v6528\ := eclat_if(work.Bool.lnot(""&\$18335_w\(31)) & 
                              eclat_if(work.Int.le(\$17456_loop665_arg\(48 to 63), eclat_resize(\$18335_w\(0 to 30),16)) & 
                              work.Int.lt(eclat_resize(\$18335_w\(0 to 30),16), 
                                          work.Int.add(\$17456_loop665_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false);
                  if \$v6528\(0) = '1' then
                    \$18323\ := \$18335_w\ & \$17456_loop665_arg\(16 to 31);
                    \$v6515\ := \$ram_lock\;
                    if \$v6515\(0) = '1' then
                      state_var7461 := Q_WAIT6514;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                              \$17456_loop665_arg\(64 to 79), \$17456_loop665_arg\(0 to 15))));
                      \$ram_write\ <= \$18323\(0 to 31); \$ram_write_request\ <= '1';
                      state_var7461 := PAUSE_SET6513;
                    end if;
                  else
                    \$v6527\ := \$ram_lock\;
                    if \$v6527\(0) = '1' then
                      state_var7461 := Q_WAIT6526;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18319\(0 to 30),16)));
                      state_var7461 := PAUSE_GET6525;
                    end if;
                  end if;
                when PAUSE_GET6533 =>
                  \$18319\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v6532\ := work.Bool.lnot(eclat_if(work.Bool.lnot(
                                                      ""&\$18319\(31)) & 
                                             eclat_if(work.Int.le(\$17456_loop665_arg\(32 to 47), eclat_resize(\$18319\(0 to 30),16)) & 
                                             work.Int.lt(eclat_resize(\$18319\(0 to 30),16), 
                                                         work.Int.add(
                                                         \$17456_loop665_arg\(32 to 47), X"1770")) & eclat_false) & eclat_false));
                  if \$v6532\(0) = '1' then
                    \$18323\ := \$18319\ & \$17456_loop665_arg\(16 to 31);
                    \$v6515\ := \$ram_lock\;
                    if \$v6515\(0) = '1' then
                      state_var7461 := Q_WAIT6514;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                              \$17456_loop665_arg\(64 to 79), \$17456_loop665_arg\(0 to 15))));
                      \$ram_write\ <= \$18323\(0 to 31); \$ram_write_request\ <= '1';
                      state_var7461 := PAUSE_SET6513;
                    end if;
                  else
                    \$v6531\ := \$ram_lock\;
                    if \$v6531\(0) = '1' then
                      state_var7461 := Q_WAIT6530;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                        eclat_resize(\$18319\(0 to 30),16), X"000" & X"1")));
                      state_var7461 := PAUSE_GET6529;
                    end if;
                  end if;
                when PAUSE_GET6537 =>
                  \$18284\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$17456_loop665_id\ := "000000100010";
                  \$17456_loop665_arg\ := X"000" & X"1" & \$17457_aux664_arg\(16 to 31) & \$17457_aux664_arg\(32 to 47) & \$17457_aux664_arg\(48 to 63) & \$17457_aux664_arg\(0 to 15) & eclat_resize(
                  work.Int.lsr(eclat_resize(eclat_resize(\$18284\(0 to 30),16),31), X"0000000" & X"2"),16);
                  state_var7461 := \$17456_LOOP665\;
                when PAUSE_GET6544 =>
                  \$18261\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v6543\ := \$ram_lock\;
                  if \$v6543\(0) = '1' then
                    state_var7461 := Q_WAIT6542;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            \$17458_loop666_arg\(16 to 31), \$17458_loop666_arg\(0 to 15))));
                    \$ram_write\ <= \$18261\; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6541;
                  end if;
                when PAUSE_GET6560 =>
                  \$18180_hd\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$18184\ := work.Print.print_string(clk,of_string("bloc "));
                  \$18185\ := work.Int.print(clk,eclat_resize(\$18159\(0 to 30),16));
                  \$18186\ := work.Print.print_string(clk,of_string(" of size "));
                  \$18187\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                              work.Int.lsr(
                                                              \$18180_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$18188\ := work.Print.print_string(clk,of_string(" from "));
                  \$18189\ := work.Int.print(clk,eclat_resize(\$18159\(0 to 30),16));
                  \$18190\ := work.Print.print_string(clk,of_string(" to "));
                  \$18191\ := work.Int.print(clk,\$17459_loop665_arg\(16 to 31));
                  \$18192\ := work.Print.print_newline(clk,eclat_unit);
                  \$v6559\ := \$ram_lock\;
                  if \$v6559\(0) = '1' then
                    state_var7461 := Q_WAIT6558;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17459_loop665_arg\(16 to 31)));
                    \$ram_write\ <= \$18180_hd\; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6557;
                  end if;
                when PAUSE_GET6564 =>
                  \$18175_w\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v6563\ := eclat_if(work.Bool.lnot(""&\$18175_w\(31)) & 
                              eclat_if(work.Int.le(\$17459_loop665_arg\(48 to 63), eclat_resize(\$18175_w\(0 to 30),16)) & 
                              work.Int.lt(eclat_resize(\$18175_w\(0 to 30),16), 
                                          work.Int.add(\$17459_loop665_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false);
                  if \$v6563\(0) = '1' then
                    \$18163\ := \$18175_w\ & \$17459_loop665_arg\(16 to 31);
                    \$v6550\ := \$ram_lock\;
                    if \$v6550\(0) = '1' then
                      state_var7461 := Q_WAIT6549;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                              \$17459_loop665_arg\(64 to 79), \$17459_loop665_arg\(0 to 15))));
                      \$ram_write\ <= \$18163\(0 to 31); \$ram_write_request\ <= '1';
                      state_var7461 := PAUSE_SET6548;
                    end if;
                  else
                    \$v6562\ := \$ram_lock\;
                    if \$v6562\(0) = '1' then
                      state_var7461 := Q_WAIT6561;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18159\(0 to 30),16)));
                      state_var7461 := PAUSE_GET6560;
                    end if;
                  end if;
                when PAUSE_GET6568 =>
                  \$18159\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v6567\ := work.Bool.lnot(eclat_if(work.Bool.lnot(
                                                      ""&\$18159\(31)) & 
                                             eclat_if(work.Int.le(\$17459_loop665_arg\(32 to 47), eclat_resize(\$18159\(0 to 30),16)) & 
                                             work.Int.lt(eclat_resize(\$18159\(0 to 30),16), 
                                                         work.Int.add(
                                                         \$17459_loop665_arg\(32 to 47), X"1770")) & eclat_false) & eclat_false));
                  if \$v6567\(0) = '1' then
                    \$18163\ := \$18159\ & \$17459_loop665_arg\(16 to 31);
                    \$v6550\ := \$ram_lock\;
                    if \$v6550\(0) = '1' then
                      state_var7461 := Q_WAIT6549;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                              \$17459_loop665_arg\(64 to 79), \$17459_loop665_arg\(0 to 15))));
                      \$ram_write\ <= \$18163\(0 to 31); \$ram_write_request\ <= '1';
                      state_var7461 := PAUSE_SET6548;
                    end if;
                  else
                    \$v6566\ := \$ram_lock\;
                    if \$v6566\(0) = '1' then
                      state_var7461 := Q_WAIT6565;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                        eclat_resize(\$18159\(0 to 30),16), X"000" & X"1")));
                      state_var7461 := PAUSE_GET6564;
                    end if;
                  end if;
                when PAUSE_GET6572 =>
                  \$18124\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$17459_loop665_id\ := "000000100100";
                  \$17459_loop665_arg\ := X"000" & X"1" & \$17460_aux664_arg\(16 to 31) & \$17460_aux664_arg\(32 to 47) & \$17460_aux664_arg\(48 to 63) & \$17460_aux664_arg\(0 to 15) & eclat_resize(
                  work.Int.lsr(eclat_resize(eclat_resize(\$18124\(0 to 30),16),31), X"0000000" & X"2"),16);
                  state_var7461 := \$17459_LOOP665\;
                when PAUSE_GET6589 =>
                  \$17585_hd\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$17589\ := work.Print.print_string(clk,of_string("bloc "));
                  \$17590\ := work.Int.print(clk,eclat_resize(\$17562\(0 to 30),16));
                  \$17591\ := work.Print.print_string(clk,of_string(" of size "));
                  \$17592\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                              work.Int.lsr(
                                                              \$17585_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$17593\ := work.Print.print_string(clk,of_string(" from "));
                  \$17594\ := work.Int.print(clk,eclat_resize(\$17562\(0 to 30),16));
                  \$17595\ := work.Print.print_string(clk,of_string(" to "));
                  \$17596\ := work.Int.print(clk,\$17547_copy_root_in_ram6635891_arg\(32 to 47));
                  \$17597\ := work.Print.print_newline(clk,eclat_unit);
                  \$v6588\ := \$ram_lock\;
                  if \$v6588\(0) = '1' then
                    state_var7461 := Q_WAIT6587;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17547_copy_root_in_ram6635891_arg\(32 to 47)));
                    \$ram_write\ <= \$17585_hd\; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6586;
                  end if;
                when PAUSE_GET6593 =>
                  \$17580_w\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v6592\ := eclat_if(work.Bool.lnot(""&\$17580_w\(31)) & 
                              eclat_if(work.Int.le(\$17547_copy_root_in_ram6635891_arg\(64 to 79), eclat_resize(\$17580_w\(0 to 30),16)) & 
                              work.Int.lt(eclat_resize(\$17580_w\(0 to 30),16), 
                                          work.Int.add(\$17547_copy_root_in_ram6635891_arg\(64 to 79), X"1770")) & eclat_false) & eclat_false);
                  if \$v6592\(0) = '1' then
                    \$17566\ := \$17580_w\ & \$17547_copy_root_in_ram6635891_arg\(32 to 47);
                    \$v6579\ := \$ram_lock\;
                    if \$v6579\(0) = '1' then
                      state_var7461 := Q_WAIT6578;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(\$17547_copy_root_in_ram6635891_arg\(0 to 15)));
                      \$ram_write\ <= \$17566\(0 to 31); \$ram_write_request\ <= '1';
                      state_var7461 := PAUSE_SET6577;
                    end if;
                  else
                    \$v6591\ := \$ram_lock\;
                    if \$v6591\(0) = '1' then
                      state_var7461 := Q_WAIT6590;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$17562\(0 to 30),16)));
                      state_var7461 := PAUSE_GET6589;
                    end if;
                  end if;
                when PAUSE_GET6597 =>
                  \$17562\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v6596\ := work.Bool.lnot(eclat_if(work.Bool.lnot(
                                                      ""&\$17562\(31)) & 
                                             eclat_if(work.Int.le(\$17547_copy_root_in_ram6635891_arg\(48 to 63), eclat_resize(\$17562\(0 to 30),16)) & 
                                             work.Int.lt(eclat_resize(\$17562\(0 to 30),16), 
                                                         work.Int.add(
                                                         \$17547_copy_root_in_ram6635891_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false));
                  if \$v6596\(0) = '1' then
                    \$17566\ := \$17562\ & \$17547_copy_root_in_ram6635891_arg\(32 to 47);
                    \$v6579\ := \$ram_lock\;
                    if \$v6579\(0) = '1' then
                      state_var7461 := Q_WAIT6578;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(\$17547_copy_root_in_ram6635891_arg\(0 to 15)));
                      \$ram_write\ <= \$17566\(0 to 31); \$ram_write_request\ <= '1';
                      state_var7461 := PAUSE_SET6577;
                    end if;
                  else
                    \$v6595\ := \$ram_lock\;
                    if \$v6595\(0) = '1' then
                      state_var7461 := Q_WAIT6594;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                        eclat_resize(\$17562\(0 to 30),16), X"000" & X"1")));
                      state_var7461 := PAUSE_GET6593;
                    end if;
                  end if;
                when PAUSE_GET6613 =>
                  \$17665_hd\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$17669\ := work.Print.print_string(clk,of_string("bloc "));
                  \$17670\ := work.Int.print(clk,eclat_resize(\$17535\(0 to 30),16));
                  \$17671\ := work.Print.print_string(clk,of_string(" of size "));
                  \$17672\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                              work.Int.lsr(
                                                              \$17665_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$17673\ := work.Print.print_string(clk,of_string(" from "));
                  \$17674\ := work.Int.print(clk,eclat_resize(\$17535\(0 to 30),16));
                  \$17675\ := work.Print.print_string(clk,of_string(" to "));
                  \$17676\ := work.Int.print(clk,\$17520_copy_root_in_ram6635893_arg\(32 to 47));
                  \$17677\ := work.Print.print_newline(clk,eclat_unit);
                  \$v6612\ := \$ram_lock\;
                  if \$v6612\(0) = '1' then
                    state_var7461 := Q_WAIT6611;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17520_copy_root_in_ram6635893_arg\(32 to 47)));
                    \$ram_write\ <= \$17665_hd\; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6610;
                  end if;
                when PAUSE_GET6617 =>
                  \$17660_w\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v6616\ := eclat_if(work.Bool.lnot(""&\$17660_w\(31)) & 
                              eclat_if(work.Int.le(\$17520_copy_root_in_ram6635893_arg\(64 to 79), eclat_resize(\$17660_w\(0 to 30),16)) & 
                              work.Int.lt(eclat_resize(\$17660_w\(0 to 30),16), 
                                          work.Int.add(\$17520_copy_root_in_ram6635893_arg\(64 to 79), X"1770")) & eclat_false) & eclat_false);
                  if \$v6616\(0) = '1' then
                    \$17539\ := \$17660_w\ & \$17520_copy_root_in_ram6635893_arg\(32 to 47);
                    \$v6603\ := \$ram_lock\;
                    if \$v6603\(0) = '1' then
                      state_var7461 := Q_WAIT6602;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(\$17520_copy_root_in_ram6635893_arg\(0 to 15)));
                      \$ram_write\ <= \$17539\(0 to 31); \$ram_write_request\ <= '1';
                      state_var7461 := PAUSE_SET6601;
                    end if;
                  else
                    \$v6615\ := \$ram_lock\;
                    if \$v6615\(0) = '1' then
                      state_var7461 := Q_WAIT6614;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$17535\(0 to 30),16)));
                      state_var7461 := PAUSE_GET6613;
                    end if;
                  end if;
                when PAUSE_GET6621 =>
                  \$17535\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v6620\ := work.Bool.lnot(eclat_if(work.Bool.lnot(
                                                      ""&\$17535\(31)) & 
                                             eclat_if(work.Int.le(\$17520_copy_root_in_ram6635893_arg\(48 to 63), eclat_resize(\$17535\(0 to 30),16)) & 
                                             work.Int.lt(eclat_resize(\$17535\(0 to 30),16), 
                                                         work.Int.add(
                                                         \$17520_copy_root_in_ram6635893_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false));
                  if \$v6620\(0) = '1' then
                    \$17539\ := \$17535\ & \$17520_copy_root_in_ram6635893_arg\(32 to 47);
                    \$v6603\ := \$ram_lock\;
                    if \$v6603\(0) = '1' then
                      state_var7461 := Q_WAIT6602;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(\$17520_copy_root_in_ram6635893_arg\(0 to 15)));
                      \$ram_write\ <= \$17539\(0 to 31); \$ram_write_request\ <= '1';
                      state_var7461 := PAUSE_SET6601;
                    end if;
                  else
                    \$v6619\ := \$ram_lock\;
                    if \$v6619\(0) = '1' then
                      state_var7461 := Q_WAIT6618;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                        eclat_resize(\$17535\(0 to 30),16), X"000" & X"1")));
                      state_var7461 := PAUSE_GET6617;
                    end if;
                  end if;
                when PAUSE_GET6625 =>
                  \$17491\ := \$global_end_value\;
                  release(\$global_end_lock\);
                  \$17520_copy_root_in_ram6635893_id\ := "000000101100";
                  \$17520_copy_root_in_ram6635893_arg\ := X"3e80" & \$17491\ & \$17490_next\ & \$17444\(96 to 111) & \$17444\(112 to 127);
                  state_var7461 := \$17520_COPY_ROOT_IN_RAM6635893\;
                when PAUSE_GET6640 =>
                  \$17799_hd\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$17803\ := work.Print.print_string(clk,of_string("bloc "));
                  \$17804\ := work.Int.print(clk,eclat_resize(\$17776\(0 to 30),16));
                  \$17805\ := work.Print.print_string(clk,of_string(" of size "));
                  \$17806\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                              work.Int.lsr(
                                                              \$17799_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$17807\ := work.Print.print_string(clk,of_string(" from "));
                  \$17808\ := work.Int.print(clk,eclat_resize(\$17776\(0 to 30),16));
                  \$17809\ := work.Print.print_string(clk,of_string(" to "));
                  \$17810\ := work.Int.print(clk,\$17761_copy_root_in_ram6635891_arg\(32 to 47));
                  \$17811\ := work.Print.print_newline(clk,eclat_unit);
                  \$v6639\ := \$ram_lock\;
                  if \$v6639\(0) = '1' then
                    state_var7461 := Q_WAIT6638;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17761_copy_root_in_ram6635891_arg\(32 to 47)));
                    \$ram_write\ <= \$17799_hd\; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6637;
                  end if;
                when PAUSE_GET6644 =>
                  \$17794_w\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v6643\ := eclat_if(work.Bool.lnot(""&\$17794_w\(31)) & 
                              eclat_if(work.Int.le(\$17761_copy_root_in_ram6635891_arg\(64 to 79), eclat_resize(\$17794_w\(0 to 30),16)) & 
                              work.Int.lt(eclat_resize(\$17794_w\(0 to 30),16), 
                                          work.Int.add(\$17761_copy_root_in_ram6635891_arg\(64 to 79), X"1770")) & eclat_false) & eclat_false);
                  if \$v6643\(0) = '1' then
                    \$17780\ := \$17794_w\ & \$17761_copy_root_in_ram6635891_arg\(32 to 47);
                    \$v6630\ := \$ram_lock\;
                    if \$v6630\(0) = '1' then
                      state_var7461 := Q_WAIT6629;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(\$17761_copy_root_in_ram6635891_arg\(0 to 15)));
                      \$ram_write\ <= \$17780\(0 to 31); \$ram_write_request\ <= '1';
                      state_var7461 := PAUSE_SET6628;
                    end if;
                  else
                    \$v6642\ := \$ram_lock\;
                    if \$v6642\(0) = '1' then
                      state_var7461 := Q_WAIT6641;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$17776\(0 to 30),16)));
                      state_var7461 := PAUSE_GET6640;
                    end if;
                  end if;
                when PAUSE_GET6648 =>
                  \$17776\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v6647\ := work.Bool.lnot(eclat_if(work.Bool.lnot(
                                                      ""&\$17776\(31)) & 
                                             eclat_if(work.Int.le(\$17761_copy_root_in_ram6635891_arg\(48 to 63), eclat_resize(\$17776\(0 to 30),16)) & 
                                             work.Int.lt(eclat_resize(\$17776\(0 to 30),16), 
                                                         work.Int.add(
                                                         \$17761_copy_root_in_ram6635891_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false));
                  if \$v6647\(0) = '1' then
                    \$17780\ := \$17776\ & \$17761_copy_root_in_ram6635891_arg\(32 to 47);
                    \$v6630\ := \$ram_lock\;
                    if \$v6630\(0) = '1' then
                      state_var7461 := Q_WAIT6629;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(\$17761_copy_root_in_ram6635891_arg\(0 to 15)));
                      \$ram_write\ <= \$17780\(0 to 31); \$ram_write_request\ <= '1';
                      state_var7461 := PAUSE_SET6628;
                    end if;
                  else
                    \$v6646\ := \$ram_lock\;
                    if \$v6646\(0) = '1' then
                      state_var7461 := Q_WAIT6645;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                        eclat_resize(\$17776\(0 to 30),16), X"000" & X"1")));
                      state_var7461 := PAUSE_GET6644;
                    end if;
                  end if;
                when PAUSE_GET6664 =>
                  \$17879_hd\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$17883\ := work.Print.print_string(clk,of_string("bloc "));
                  \$17884\ := work.Int.print(clk,eclat_resize(\$17749\(0 to 30),16));
                  \$17885\ := work.Print.print_string(clk,of_string(" of size "));
                  \$17886\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                              work.Int.lsr(
                                                              \$17879_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$17887\ := work.Print.print_string(clk,of_string(" from "));
                  \$17888\ := work.Int.print(clk,eclat_resize(\$17749\(0 to 30),16));
                  \$17889\ := work.Print.print_string(clk,of_string(" to "));
                  \$17890\ := work.Int.print(clk,\$17734_copy_root_in_ram6635892_arg\(32 to 47));
                  \$17891\ := work.Print.print_newline(clk,eclat_unit);
                  \$v6663\ := \$ram_lock\;
                  if \$v6663\(0) = '1' then
                    state_var7461 := Q_WAIT6662;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17734_copy_root_in_ram6635892_arg\(32 to 47)));
                    \$ram_write\ <= \$17879_hd\; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6661;
                  end if;
                when PAUSE_GET6668 =>
                  \$17874_w\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v6667\ := eclat_if(work.Bool.lnot(""&\$17874_w\(31)) & 
                              eclat_if(work.Int.le(\$17734_copy_root_in_ram6635892_arg\(64 to 79), eclat_resize(\$17874_w\(0 to 30),16)) & 
                              work.Int.lt(eclat_resize(\$17874_w\(0 to 30),16), 
                                          work.Int.add(\$17734_copy_root_in_ram6635892_arg\(64 to 79), X"1770")) & eclat_false) & eclat_false);
                  if \$v6667\(0) = '1' then
                    \$17753\ := \$17874_w\ & \$17734_copy_root_in_ram6635892_arg\(32 to 47);
                    \$v6654\ := \$ram_lock\;
                    if \$v6654\(0) = '1' then
                      state_var7461 := Q_WAIT6653;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(\$17734_copy_root_in_ram6635892_arg\(0 to 15)));
                      \$ram_write\ <= \$17753\(0 to 31); \$ram_write_request\ <= '1';
                      state_var7461 := PAUSE_SET6652;
                    end if;
                  else
                    \$v6666\ := \$ram_lock\;
                    if \$v6666\(0) = '1' then
                      state_var7461 := Q_WAIT6665;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$17749\(0 to 30),16)));
                      state_var7461 := PAUSE_GET6664;
                    end if;
                  end if;
                when PAUSE_GET6672 =>
                  \$17749\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v6671\ := work.Bool.lnot(eclat_if(work.Bool.lnot(
                                                      ""&\$17749\(31)) & 
                                             eclat_if(work.Int.le(\$17734_copy_root_in_ram6635892_arg\(48 to 63), eclat_resize(\$17749\(0 to 30),16)) & 
                                             work.Int.lt(eclat_resize(\$17749\(0 to 30),16), 
                                                         work.Int.add(
                                                         \$17734_copy_root_in_ram6635892_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false));
                  if \$v6671\(0) = '1' then
                    \$17753\ := \$17749\ & \$17734_copy_root_in_ram6635892_arg\(32 to 47);
                    \$v6654\ := \$ram_lock\;
                    if \$v6654\(0) = '1' then
                      state_var7461 := Q_WAIT6653;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(\$17734_copy_root_in_ram6635892_arg\(0 to 15)));
                      \$ram_write\ <= \$17753\(0 to 31); \$ram_write_request\ <= '1';
                      state_var7461 := PAUSE_SET6652;
                    end if;
                  else
                    \$v6670\ := \$ram_lock\;
                    if \$v6670\(0) = '1' then
                      state_var7461 := Q_WAIT6669;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                        eclat_resize(\$17749\(0 to 30),16), X"000" & X"1")));
                      state_var7461 := PAUSE_GET6668;
                    end if;
                  end if;
                when PAUSE_GET6685 =>
                  \$17957_hd\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$17961\ := work.Print.print_string(clk,of_string("bloc "));
                  \$17962\ := work.Int.print(clk,eclat_resize(\$13922_wait662_arg\(33 to 63),16));
                  \$17963\ := work.Print.print_string(clk,of_string(" of size "));
                  \$17964\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                              work.Int.lsr(
                                                              \$17957_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$17965\ := work.Print.print_string(clk,of_string(" from "));
                  \$17966\ := work.Int.print(clk,eclat_resize(\$13922_wait662_arg\(33 to 63),16));
                  \$17967\ := work.Print.print_string(clk,of_string(" to "));
                  \$17968\ := work.Int.print(clk,\$17470\(32 to 47));
                  \$17969\ := work.Print.print_newline(clk,eclat_unit);
                  \$v6684\ := \$ram_lock\;
                  if \$v6684\(0) = '1' then
                    state_var7461 := Q_WAIT6683;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17470\(32 to 47)));
                    \$ram_write\ <= \$17957_hd\; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6682;
                  end if;
                when PAUSE_GET6689 =>
                  \$17952_w\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v6688\ := eclat_if(work.Bool.lnot(""&\$17952_w\(31)) & 
                              eclat_if(work.Int.le(\$17444\(112 to 127), eclat_resize(\$17952_w\(0 to 30),16)) & 
                              work.Int.lt(eclat_resize(\$17952_w\(0 to 30),16), 
                                          work.Int.add(\$17444\(112 to 127), X"1770")) & eclat_false) & eclat_false);
                  if \$v6688\(0) = '1' then
                    \$17487\ := \$17952_w\ & \$17470\(32 to 47);
                    \$17734_copy_root_in_ram6635892_id\ := "000000110000";
                    \$17734_copy_root_in_ram6635892_arg\ := X"0" & X"3e8" & \$13922_wait662_arg\(65 to 80) & \$17487\(32 to 47) & \$17444\(96 to 111) & \$17444\(112 to 127);
                    state_var7461 := \$17734_COPY_ROOT_IN_RAM6635892\;
                  else
                    \$v6687\ := \$ram_lock\;
                    if \$v6687\(0) = '1' then
                      state_var7461 := Q_WAIT6686;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$13922_wait662_arg\(33 to 63),16)));
                      state_var7461 := PAUSE_GET6685;
                    end if;
                  end if;
                when PAUSE_GET6702 =>
                  \$18035_hd\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$18039\ := work.Print.print_string(clk,of_string("bloc "));
                  \$18040\ := work.Int.print(clk,eclat_resize(\$13922_wait662_arg\(1 to 31),16));
                  \$18041\ := work.Print.print_string(clk,of_string(" of size "));
                  \$18042\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                              work.Int.lsr(
                                                              \$18035_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$18043\ := work.Print.print_string(clk,of_string(" from "));
                  \$18044\ := work.Int.print(clk,eclat_resize(\$13922_wait662_arg\(1 to 31),16));
                  \$18045\ := work.Print.print_string(clk,of_string(" to "));
                  \$18046\ := work.Int.print(clk,\$17444\(112 to 127));
                  \$18047\ := work.Print.print_newline(clk,eclat_unit);
                  \$v6701\ := \$ram_lock\;
                  if \$v6701\(0) = '1' then
                    state_var7461 := Q_WAIT6700;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17444\(112 to 127)));
                    \$ram_write\ <= \$18035_hd\; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6699;
                  end if;
                when PAUSE_GET6706 =>
                  \$18030_w\ := \$ram_value\;
                  release(\$ram_lock\);
                  \$v6705\ := eclat_if(work.Bool.lnot(""&\$18030_w\(31)) & 
                              eclat_if(work.Int.le(\$17444\(112 to 127), eclat_resize(\$18030_w\(0 to 30),16)) & 
                              work.Int.lt(eclat_resize(\$18030_w\(0 to 30),16), 
                                          work.Int.add(\$17444\(112 to 127), X"1770")) & eclat_false) & eclat_false);
                  if \$v6705\(0) = '1' then
                    \$17470\ := \$18030_w\ & \$17444\(112 to 127);
                    \$v6692\ := work.Bool.lnot(eclat_if(work.Bool.lnot(
                                                        ""&\$13922_wait662_arg\(64)) & 
                                               eclat_if(work.Int.le(\$17444\(96 to 111), eclat_resize(\$13922_wait662_arg\(33 to 63),16)) & 
                                               work.Int.lt(eclat_resize(\$13922_wait662_arg\(33 to 63),16), 
                                                           work.Int.add(
                                                           \$17444\(96 to 111), X"1770")) & eclat_false) & eclat_false));
                    if \$v6692\(0) = '1' then
                      \$17487\ := \$13922_wait662_arg\(33 to 64) & \$17470\(32 to 47);
                      \$17734_copy_root_in_ram6635892_id\ := "000000110000";
                      \$17734_copy_root_in_ram6635892_arg\ := X"0" & X"3e8" & \$13922_wait662_arg\(65 to 80) & \$17487\(32 to 47) & \$17444\(96 to 111) & \$17444\(112 to 127);
                      state_var7461 := \$17734_COPY_ROOT_IN_RAM6635892\;
                    else
                      \$v6691\ := \$ram_lock\;
                      if \$v6691\(0) = '1' then
                        state_var7461 := Q_WAIT6690;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$13922_wait662_arg\(33 to 63),16), X"000" & X"1")));
                        state_var7461 := PAUSE_GET6689;
                      end if;
                    end if;
                  else
                    \$v6704\ := \$ram_lock\;
                    if \$v6704\(0) = '1' then
                      state_var7461 := Q_WAIT6703;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$13922_wait662_arg\(1 to 31),16)));
                      state_var7461 := PAUSE_GET6702;
                    end if;
                  end if;
                when PAUSE_SET6506 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$18422\ := eclat_unit;
                  \$17455_loop666_arg\ := work.Int.add(\$17455_loop666_arg\(0 to 15), X"000" & X"1") & \$17455_loop666_arg\(16 to 31) & \$17455_loop666_arg\(32 to 47) & \$17455_loop666_arg\(48 to 63);
                  state_var7461 := \$17455_LOOP666\;
                when PAUSE_SET6513 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$18326\ := eclat_unit;
                  \$17456_loop665_arg\ := work.Int.add(\$17456_loop665_arg\(0 to 15), X"000" & X"1") & \$18323\(32 to 47) & \$17456_loop665_arg\(32 to 47) & \$17456_loop665_arg\(48 to 63) & \$17456_loop665_arg\(64 to 79) & \$17456_loop665_arg\(80 to 95);
                  state_var7461 := \$17456_LOOP665\;
                when PAUSE_SET6516 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$18356\ := eclat_unit;
                  \$18323\ := eclat_resize(\$17456_loop665_arg\(16 to 31),31) & eclat_false & 
                  work.Int.add(\$17456_loop665_arg\(16 to 31), work.Int.add(
                                                               eclat_resize(
                                                               work.Int.lsr(
                                                               \$18340_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$v6515\ := \$ram_lock\;
                  if \$v6515\(0) = '1' then
                    state_var7461 := Q_WAIT6514;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            \$17456_loop665_arg\(64 to 79), \$17456_loop665_arg\(0 to 15))));
                    \$ram_write\ <= \$18323\(0 to 31); \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6513;
                  end if;
                when PAUSE_SET6519 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$18355\ := eclat_unit;
                  \$v6518\ := \$ram_lock\;
                  if \$v6518\(0) = '1' then
                    state_var7461 := Q_WAIT6517;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$18319\(0 to 30),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$17456_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6516;
                  end if;
                when PAUSE_SET6522 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$18353\ := eclat_unit;
                  \$17455_loop666_id\ := "000000100001";
                  \$17455_loop666_arg\ := X"000" & X"1" & \$17456_loop665_arg\(16 to 31) & eclat_resize(\$18319\(0 to 30),16) & eclat_resize(
                  work.Int.lsr(\$18340_hd\(0 to 30), X"0000000" & X"2"),16);
                  state_var7461 := \$17455_LOOP666\;
                when PAUSE_SET6541 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$18262\ := eclat_unit;
                  \$17458_loop666_arg\ := work.Int.add(\$17458_loop666_arg\(0 to 15), X"000" & X"1") & \$17458_loop666_arg\(16 to 31) & \$17458_loop666_arg\(32 to 47) & \$17458_loop666_arg\(48 to 63);
                  state_var7461 := \$17458_LOOP666\;
                when PAUSE_SET6548 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$18166\ := eclat_unit;
                  \$17459_loop665_arg\ := work.Int.add(\$17459_loop665_arg\(0 to 15), X"000" & X"1") & \$18163\(32 to 47) & \$17459_loop665_arg\(32 to 47) & \$17459_loop665_arg\(48 to 63) & \$17459_loop665_arg\(64 to 79) & \$17459_loop665_arg\(80 to 95);
                  state_var7461 := \$17459_LOOP665\;
                when PAUSE_SET6551 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$18196\ := eclat_unit;
                  \$18163\ := eclat_resize(\$17459_loop665_arg\(16 to 31),31) & eclat_false & 
                  work.Int.add(\$17459_loop665_arg\(16 to 31), work.Int.add(
                                                               eclat_resize(
                                                               work.Int.lsr(
                                                               \$18180_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$v6550\ := \$ram_lock\;
                  if \$v6550\(0) = '1' then
                    state_var7461 := Q_WAIT6549;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            \$17459_loop665_arg\(64 to 79), \$17459_loop665_arg\(0 to 15))));
                    \$ram_write\ <= \$18163\(0 to 31); \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6548;
                  end if;
                when PAUSE_SET6554 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$18195\ := eclat_unit;
                  \$v6553\ := \$ram_lock\;
                  if \$v6553\(0) = '1' then
                    state_var7461 := Q_WAIT6552;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$18159\(0 to 30),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$17459_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6551;
                  end if;
                when PAUSE_SET6557 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$18193\ := eclat_unit;
                  \$17458_loop666_id\ := "000000100011";
                  \$17458_loop666_arg\ := X"000" & X"1" & \$17459_loop665_arg\(16 to 31) & eclat_resize(\$18159\(0 to 30),16) & eclat_resize(
                  work.Int.lsr(\$18180_hd\(0 to 30), X"0000000" & X"2"),16);
                  state_var7461 := \$17458_LOOP666\;
                when PAUSE_SET6577 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$17569\ := eclat_unit;
                  \$17570\ := work.Print.print_string(clk,of_string(" next="));
                  \$17571\ := work.Int.print(clk,\$17566\(32 to 47));
                  \$17572\ := work.Print.print_newline(clk,eclat_unit);
                  \$17547_copy_root_in_ram6635891_arg\ := work.Int.add(
                                                          \$17547_copy_root_in_ram6635891_arg\(0 to 15), X"000" & X"1") & \$17547_copy_root_in_ram6635891_arg\(16 to 31) & \$17566\(32 to 47) & \$17547_copy_root_in_ram6635891_arg\(48 to 63) & \$17547_copy_root_in_ram6635891_arg\(64 to 79);
                  state_var7461 := \$17547_COPY_ROOT_IN_RAM6635891\;
                when PAUSE_SET6580 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$17601\ := eclat_unit;
                  \$17566\ := eclat_resize(\$17547_copy_root_in_ram6635891_arg\(32 to 47),31) & eclat_false & 
                  work.Int.add(\$17547_copy_root_in_ram6635891_arg\(32 to 47), 
                               work.Int.add(eclat_resize(work.Int.lsr(
                                                         \$17585_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$v6579\ := \$ram_lock\;
                  if \$v6579\(0) = '1' then
                    state_var7461 := Q_WAIT6578;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17547_copy_root_in_ram6635891_arg\(0 to 15)));
                    \$ram_write\ <= \$17566\(0 to 31); \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6577;
                  end if;
                when PAUSE_SET6583 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$17600\ := eclat_unit;
                  \$v6582\ := \$ram_lock\;
                  if \$v6582\(0) = '1' then
                    state_var7461 := Q_WAIT6581;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$17562\(0 to 30),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$17547_copy_root_in_ram6635891_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6580;
                  end if;
                when PAUSE_SET6586 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$17598\ := eclat_unit;
                  \$17458_loop666_id\ := "000000101001";
                  \$17458_loop666_arg\ := X"000" & X"1" & \$17547_copy_root_in_ram6635891_arg\(32 to 47) & eclat_resize(\$17562\(0 to 30),16) & eclat_resize(
                  work.Int.lsr(\$17585_hd\(0 to 30), X"0000000" & X"2"),16);
                  state_var7461 := \$17458_LOOP666\;
                when PAUSE_SET6601 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$17542\ := eclat_unit;
                  \$17543\ := work.Print.print_string(clk,of_string(" next="));
                  \$17544\ := work.Int.print(clk,\$17539\(32 to 47));
                  \$17545\ := work.Print.print_newline(clk,eclat_unit);
                  \$17547_copy_root_in_ram6635891_id\ := "000000101010";
                  \$17547_copy_root_in_ram6635891_arg\ := work.Int.add(
                                                          \$17520_copy_root_in_ram6635893_arg\(0 to 15), X"000" & X"1") & \$17520_copy_root_in_ram6635893_arg\(16 to 31) & \$17539\(32 to 47) & \$17520_copy_root_in_ram6635893_arg\(48 to 63) & \$17520_copy_root_in_ram6635893_arg\(64 to 79);
                  state_var7461 := \$17547_COPY_ROOT_IN_RAM6635891\;
                when PAUSE_SET6604 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$17681\ := eclat_unit;
                  \$17539\ := eclat_resize(\$17520_copy_root_in_ram6635893_arg\(32 to 47),31) & eclat_false & 
                  work.Int.add(\$17520_copy_root_in_ram6635893_arg\(32 to 47), 
                               work.Int.add(eclat_resize(work.Int.lsr(
                                                         \$17665_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$v6603\ := \$ram_lock\;
                  if \$v6603\(0) = '1' then
                    state_var7461 := Q_WAIT6602;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17520_copy_root_in_ram6635893_arg\(0 to 15)));
                    \$ram_write\ <= \$17539\(0 to 31); \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6601;
                  end if;
                when PAUSE_SET6607 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$17680\ := eclat_unit;
                  \$v6606\ := \$ram_lock\;
                  if \$v6606\(0) = '1' then
                    state_var7461 := Q_WAIT6605;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$17535\(0 to 30),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$17520_copy_root_in_ram6635893_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6604;
                  end if;
                when PAUSE_SET6610 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$17678\ := eclat_unit;
                  \$17458_loop666_id\ := "000000101011";
                  \$17458_loop666_arg\ := X"000" & X"1" & \$17520_copy_root_in_ram6635893_arg\(32 to 47) & eclat_resize(\$17535\(0 to 30),16) & eclat_resize(
                  work.Int.lsr(\$17665_hd\(0 to 30), X"0000000" & X"2"),16);
                  state_var7461 := \$17458_LOOP666\;
                when PAUSE_SET6628 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$17783\ := eclat_unit;
                  \$17784\ := work.Print.print_string(clk,of_string(" next="));
                  \$17785\ := work.Int.print(clk,\$17780\(32 to 47));
                  \$17786\ := work.Print.print_newline(clk,eclat_unit);
                  \$17761_copy_root_in_ram6635891_arg\ := work.Int.add(
                                                          \$17761_copy_root_in_ram6635891_arg\(0 to 15), X"000" & X"1") & \$17761_copy_root_in_ram6635891_arg\(16 to 31) & \$17780\(32 to 47) & \$17761_copy_root_in_ram6635891_arg\(48 to 63) & \$17761_copy_root_in_ram6635891_arg\(64 to 79);
                  state_var7461 := \$17761_COPY_ROOT_IN_RAM6635891\;
                when PAUSE_SET6631 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$17815\ := eclat_unit;
                  \$17780\ := eclat_resize(\$17761_copy_root_in_ram6635891_arg\(32 to 47),31) & eclat_false & 
                  work.Int.add(\$17761_copy_root_in_ram6635891_arg\(32 to 47), 
                               work.Int.add(eclat_resize(work.Int.lsr(
                                                         \$17799_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$v6630\ := \$ram_lock\;
                  if \$v6630\(0) = '1' then
                    state_var7461 := Q_WAIT6629;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17761_copy_root_in_ram6635891_arg\(0 to 15)));
                    \$ram_write\ <= \$17780\(0 to 31); \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6628;
                  end if;
                when PAUSE_SET6634 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$17814\ := eclat_unit;
                  \$v6633\ := \$ram_lock\;
                  if \$v6633\(0) = '1' then
                    state_var7461 := Q_WAIT6632;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$17776\(0 to 30),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$17761_copy_root_in_ram6635891_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6631;
                  end if;
                when PAUSE_SET6637 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$17812\ := eclat_unit;
                  \$17458_loop666_id\ := "000000101101";
                  \$17458_loop666_arg\ := X"000" & X"1" & \$17761_copy_root_in_ram6635891_arg\(32 to 47) & eclat_resize(\$17776\(0 to 30),16) & eclat_resize(
                  work.Int.lsr(\$17799_hd\(0 to 30), X"0000000" & X"2"),16);
                  state_var7461 := \$17458_LOOP666\;
                when PAUSE_SET6652 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$17756\ := eclat_unit;
                  \$17757\ := work.Print.print_string(clk,of_string(" next="));
                  \$17758\ := work.Int.print(clk,\$17753\(32 to 47));
                  \$17759\ := work.Print.print_newline(clk,eclat_unit);
                  \$17761_copy_root_in_ram6635891_id\ := "000000101110";
                  \$17761_copy_root_in_ram6635891_arg\ := work.Int.add(
                                                          \$17734_copy_root_in_ram6635892_arg\(0 to 15), X"000" & X"1") & \$17734_copy_root_in_ram6635892_arg\(16 to 31) & \$17753\(32 to 47) & \$17734_copy_root_in_ram6635892_arg\(48 to 63) & \$17734_copy_root_in_ram6635892_arg\(64 to 79);
                  state_var7461 := \$17761_COPY_ROOT_IN_RAM6635891\;
                when PAUSE_SET6655 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$17895\ := eclat_unit;
                  \$17753\ := eclat_resize(\$17734_copy_root_in_ram6635892_arg\(32 to 47),31) & eclat_false & 
                  work.Int.add(\$17734_copy_root_in_ram6635892_arg\(32 to 47), 
                               work.Int.add(eclat_resize(work.Int.lsr(
                                                         \$17879_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$v6654\ := \$ram_lock\;
                  if \$v6654\(0) = '1' then
                    state_var7461 := Q_WAIT6653;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17734_copy_root_in_ram6635892_arg\(0 to 15)));
                    \$ram_write\ <= \$17753\(0 to 31); \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6652;
                  end if;
                when PAUSE_SET6658 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$17894\ := eclat_unit;
                  \$v6657\ := \$ram_lock\;
                  if \$v6657\(0) = '1' then
                    state_var7461 := Q_WAIT6656;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$17749\(0 to 30),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$17734_copy_root_in_ram6635892_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6655;
                  end if;
                when PAUSE_SET6661 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$17892\ := eclat_unit;
                  \$17458_loop666_id\ := "000000101111";
                  \$17458_loop666_arg\ := X"000" & X"1" & \$17734_copy_root_in_ram6635892_arg\(32 to 47) & eclat_resize(\$17749\(0 to 30),16) & eclat_resize(
                  work.Int.lsr(\$17879_hd\(0 to 30), X"0000000" & X"2"),16);
                  state_var7461 := \$17458_LOOP666\;
                when PAUSE_SET6676 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$17973\ := eclat_unit;
                  \$17487\ := eclat_resize(\$17470\(32 to 47),31) & eclat_false & 
                  work.Int.add(\$17470\(32 to 47), work.Int.add(eclat_resize(
                                                                work.Int.lsr(
                                                                \$17957_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$17734_copy_root_in_ram6635892_id\ := "000000110000";
                  \$17734_copy_root_in_ram6635892_arg\ := X"0" & X"3e8" & \$13922_wait662_arg\(65 to 80) & \$17487\(32 to 47) & \$17444\(96 to 111) & \$17444\(112 to 127);
                  state_var7461 := \$17734_COPY_ROOT_IN_RAM6635892\;
                when PAUSE_SET6679 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$17972\ := eclat_unit;
                  \$v6678\ := \$ram_lock\;
                  if \$v6678\(0) = '1' then
                    state_var7461 := Q_WAIT6677;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$13922_wait662_arg\(33 to 63),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$17470\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6676;
                  end if;
                when PAUSE_SET6682 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$17970\ := eclat_unit;
                  \$17458_loop666_id\ := "000000110001";
                  \$17458_loop666_arg\ := X"000" & X"1" & \$17470\(32 to 47) & eclat_resize(\$13922_wait662_arg\(33 to 63),16) & eclat_resize(
                  work.Int.lsr(\$17957_hd\(0 to 30), X"0000000" & X"2"),16);
                  state_var7461 := \$17458_LOOP666\;
                when PAUSE_SET6693 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$18051\ := eclat_unit;
                  \$17470\ := eclat_resize(\$17444\(112 to 127),31) & eclat_false & 
                  work.Int.add(\$17444\(112 to 127), work.Int.add(eclat_resize(
                                                                  work.Int.lsr(
                                                                  \$18035_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                  \$v6692\ := work.Bool.lnot(eclat_if(work.Bool.lnot(
                                                      ""&\$13922_wait662_arg\(64)) & 
                                             eclat_if(work.Int.le(\$17444\(96 to 111), eclat_resize(\$13922_wait662_arg\(33 to 63),16)) & 
                                             work.Int.lt(eclat_resize(\$13922_wait662_arg\(33 to 63),16), 
                                                         work.Int.add(
                                                         \$17444\(96 to 111), X"1770")) & eclat_false) & eclat_false));
                  if \$v6692\(0) = '1' then
                    \$17487\ := \$13922_wait662_arg\(33 to 64) & \$17470\(32 to 47);
                    \$17734_copy_root_in_ram6635892_id\ := "000000110000";
                    \$17734_copy_root_in_ram6635892_arg\ := X"0" & X"3e8" & \$13922_wait662_arg\(65 to 80) & \$17487\(32 to 47) & \$17444\(96 to 111) & \$17444\(112 to 127);
                    state_var7461 := \$17734_COPY_ROOT_IN_RAM6635892\;
                  else
                    \$v6691\ := \$ram_lock\;
                    if \$v6691\(0) = '1' then
                      state_var7461 := Q_WAIT6690;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                        eclat_resize(\$13922_wait662_arg\(33 to 63),16), X"000" & X"1")));
                      state_var7461 := PAUSE_GET6689;
                    end if;
                  end if;
                when PAUSE_SET6696 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$18050\ := eclat_unit;
                  \$v6695\ := \$ram_lock\;
                  if \$v6695\(0) = '1' then
                    state_var7461 := Q_WAIT6694;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$13922_wait662_arg\(1 to 31),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$17444\(112 to 127),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6693;
                  end if;
                when PAUSE_SET6699 =>
                  \$ram_write_request\ <= '0';
                  release(\$ram_lock\);
                  \$18048\ := eclat_unit;
                  \$17458_loop666_id\ := "000000110010";
                  \$17458_loop666_arg\ := X"000" & X"1" & \$17444\(112 to 127) & eclat_resize(\$13922_wait662_arg\(1 to 31),16) & eclat_resize(
                  work.Int.lsr(\$18035_hd\(0 to 30), X"0000000" & X"2"),16);
                  state_var7461 := \$17458_LOOP666\;
                when Q_WAIT6507 =>
                  \$v6508\ := \$ram_lock\;
                  if \$v6508\(0) = '1' then
                    state_var7461 := Q_WAIT6507;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            \$17455_loop666_arg\(16 to 31), \$17455_loop666_arg\(0 to 15))));
                    \$ram_write\ <= \$18421\; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6506;
                  end if;
                when Q_WAIT6510 =>
                  \$v6511\ := \$ram_lock\;
                  if \$v6511\(0) = '1' then
                    state_var7461 := Q_WAIT6510;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$17455_loop666_arg\(32 to 47), \$17455_loop666_arg\(0 to 15))));
                    state_var7461 := PAUSE_GET6509;
                  end if;
                when Q_WAIT6514 =>
                  \$v6515\ := \$ram_lock\;
                  if \$v6515\(0) = '1' then
                    state_var7461 := Q_WAIT6514;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            \$17456_loop665_arg\(64 to 79), \$17456_loop665_arg\(0 to 15))));
                    \$ram_write\ <= \$18323\(0 to 31); \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6513;
                  end if;
                when Q_WAIT6517 =>
                  \$v6518\ := \$ram_lock\;
                  if \$v6518\(0) = '1' then
                    state_var7461 := Q_WAIT6517;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$18319\(0 to 30),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$17456_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6516;
                  end if;
                when Q_WAIT6520 =>
                  \$v6521\ := \$ram_lock\;
                  if \$v6521\(0) = '1' then
                    state_var7461 := Q_WAIT6520;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18319\(0 to 30),16)));
                    \$ram_write\ <= eclat_resize(\$17456_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6519;
                  end if;
                when Q_WAIT6523 =>
                  \$v6524\ := \$ram_lock\;
                  if \$v6524\(0) = '1' then
                    state_var7461 := Q_WAIT6523;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17456_loop665_arg\(16 to 31)));
                    \$ram_write\ <= \$18340_hd\; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6522;
                  end if;
                when Q_WAIT6526 =>
                  \$v6527\ := \$ram_lock\;
                  if \$v6527\(0) = '1' then
                    state_var7461 := Q_WAIT6526;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18319\(0 to 30),16)));
                    state_var7461 := PAUSE_GET6525;
                  end if;
                when Q_WAIT6530 =>
                  \$v6531\ := \$ram_lock\;
                  if \$v6531\(0) = '1' then
                    state_var7461 := Q_WAIT6530;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18319\(0 to 30),16), X"000" & X"1")));
                    state_var7461 := PAUSE_GET6529;
                  end if;
                when Q_WAIT6534 =>
                  \$v6535\ := \$ram_lock\;
                  if \$v6535\(0) = '1' then
                    state_var7461 := Q_WAIT6534;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$17456_loop665_arg\(64 to 79), \$17456_loop665_arg\(0 to 15))));
                    state_var7461 := PAUSE_GET6533;
                  end if;
                when Q_WAIT6538 =>
                  \$v6539\ := \$ram_lock\;
                  if \$v6539\(0) = '1' then
                    state_var7461 := Q_WAIT6538;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(\$17457_aux664_arg\(0 to 15)));
                    state_var7461 := PAUSE_GET6537;
                  end if;
                when Q_WAIT6542 =>
                  \$v6543\ := \$ram_lock\;
                  if \$v6543\(0) = '1' then
                    state_var7461 := Q_WAIT6542;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            \$17458_loop666_arg\(16 to 31), \$17458_loop666_arg\(0 to 15))));
                    \$ram_write\ <= \$18261\; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6541;
                  end if;
                when Q_WAIT6545 =>
                  \$v6546\ := \$ram_lock\;
                  if \$v6546\(0) = '1' then
                    state_var7461 := Q_WAIT6545;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$17458_loop666_arg\(32 to 47), \$17458_loop666_arg\(0 to 15))));
                    state_var7461 := PAUSE_GET6544;
                  end if;
                when Q_WAIT6549 =>
                  \$v6550\ := \$ram_lock\;
                  if \$v6550\(0) = '1' then
                    state_var7461 := Q_WAIT6549;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            \$17459_loop665_arg\(64 to 79), \$17459_loop665_arg\(0 to 15))));
                    \$ram_write\ <= \$18163\(0 to 31); \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6548;
                  end if;
                when Q_WAIT6552 =>
                  \$v6553\ := \$ram_lock\;
                  if \$v6553\(0) = '1' then
                    state_var7461 := Q_WAIT6552;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$18159\(0 to 30),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$17459_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6551;
                  end if;
                when Q_WAIT6555 =>
                  \$v6556\ := \$ram_lock\;
                  if \$v6556\(0) = '1' then
                    state_var7461 := Q_WAIT6555;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18159\(0 to 30),16)));
                    \$ram_write\ <= eclat_resize(\$17459_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6554;
                  end if;
                when Q_WAIT6558 =>
                  \$v6559\ := \$ram_lock\;
                  if \$v6559\(0) = '1' then
                    state_var7461 := Q_WAIT6558;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17459_loop665_arg\(16 to 31)));
                    \$ram_write\ <= \$18180_hd\; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6557;
                  end if;
                when Q_WAIT6561 =>
                  \$v6562\ := \$ram_lock\;
                  if \$v6562\(0) = '1' then
                    state_var7461 := Q_WAIT6561;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18159\(0 to 30),16)));
                    state_var7461 := PAUSE_GET6560;
                  end if;
                when Q_WAIT6565 =>
                  \$v6566\ := \$ram_lock\;
                  if \$v6566\(0) = '1' then
                    state_var7461 := Q_WAIT6565;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18159\(0 to 30),16), X"000" & X"1")));
                    state_var7461 := PAUSE_GET6564;
                  end if;
                when Q_WAIT6569 =>
                  \$v6570\ := \$ram_lock\;
                  if \$v6570\(0) = '1' then
                    state_var7461 := Q_WAIT6569;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$17459_loop665_arg\(64 to 79), \$17459_loop665_arg\(0 to 15))));
                    state_var7461 := PAUSE_GET6568;
                  end if;
                when Q_WAIT6573 =>
                  \$v6574\ := \$ram_lock\;
                  if \$v6574\(0) = '1' then
                    state_var7461 := Q_WAIT6573;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(\$17460_aux664_arg\(0 to 15)));
                    state_var7461 := PAUSE_GET6572;
                  end if;
                when Q_WAIT6578 =>
                  \$v6579\ := \$ram_lock\;
                  if \$v6579\(0) = '1' then
                    state_var7461 := Q_WAIT6578;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17547_copy_root_in_ram6635891_arg\(0 to 15)));
                    \$ram_write\ <= \$17566\(0 to 31); \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6577;
                  end if;
                when Q_WAIT6581 =>
                  \$v6582\ := \$ram_lock\;
                  if \$v6582\(0) = '1' then
                    state_var7461 := Q_WAIT6581;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$17562\(0 to 30),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$17547_copy_root_in_ram6635891_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6580;
                  end if;
                when Q_WAIT6584 =>
                  \$v6585\ := \$ram_lock\;
                  if \$v6585\(0) = '1' then
                    state_var7461 := Q_WAIT6584;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$17562\(0 to 30),16)));
                    \$ram_write\ <= eclat_resize(\$17547_copy_root_in_ram6635891_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6583;
                  end if;
                when Q_WAIT6587 =>
                  \$v6588\ := \$ram_lock\;
                  if \$v6588\(0) = '1' then
                    state_var7461 := Q_WAIT6587;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17547_copy_root_in_ram6635891_arg\(32 to 47)));
                    \$ram_write\ <= \$17585_hd\; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6586;
                  end if;
                when Q_WAIT6590 =>
                  \$v6591\ := \$ram_lock\;
                  if \$v6591\(0) = '1' then
                    state_var7461 := Q_WAIT6590;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$17562\(0 to 30),16)));
                    state_var7461 := PAUSE_GET6589;
                  end if;
                when Q_WAIT6594 =>
                  \$v6595\ := \$ram_lock\;
                  if \$v6595\(0) = '1' then
                    state_var7461 := Q_WAIT6594;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$17562\(0 to 30),16), X"000" & X"1")));
                    state_var7461 := PAUSE_GET6593;
                  end if;
                when Q_WAIT6598 =>
                  \$v6599\ := \$ram_lock\;
                  if \$v6599\(0) = '1' then
                    state_var7461 := Q_WAIT6598;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(\$17547_copy_root_in_ram6635891_arg\(0 to 15)));
                    state_var7461 := PAUSE_GET6597;
                  end if;
                when Q_WAIT6602 =>
                  \$v6603\ := \$ram_lock\;
                  if \$v6603\(0) = '1' then
                    state_var7461 := Q_WAIT6602;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17520_copy_root_in_ram6635893_arg\(0 to 15)));
                    \$ram_write\ <= \$17539\(0 to 31); \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6601;
                  end if;
                when Q_WAIT6605 =>
                  \$v6606\ := \$ram_lock\;
                  if \$v6606\(0) = '1' then
                    state_var7461 := Q_WAIT6605;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$17535\(0 to 30),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$17520_copy_root_in_ram6635893_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6604;
                  end if;
                when Q_WAIT6608 =>
                  \$v6609\ := \$ram_lock\;
                  if \$v6609\(0) = '1' then
                    state_var7461 := Q_WAIT6608;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$17535\(0 to 30),16)));
                    \$ram_write\ <= eclat_resize(\$17520_copy_root_in_ram6635893_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6607;
                  end if;
                when Q_WAIT6611 =>
                  \$v6612\ := \$ram_lock\;
                  if \$v6612\(0) = '1' then
                    state_var7461 := Q_WAIT6611;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17520_copy_root_in_ram6635893_arg\(32 to 47)));
                    \$ram_write\ <= \$17665_hd\; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6610;
                  end if;
                when Q_WAIT6614 =>
                  \$v6615\ := \$ram_lock\;
                  if \$v6615\(0) = '1' then
                    state_var7461 := Q_WAIT6614;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$17535\(0 to 30),16)));
                    state_var7461 := PAUSE_GET6613;
                  end if;
                when Q_WAIT6618 =>
                  \$v6619\ := \$ram_lock\;
                  if \$v6619\(0) = '1' then
                    state_var7461 := Q_WAIT6618;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$17535\(0 to 30),16), X"000" & X"1")));
                    state_var7461 := PAUSE_GET6617;
                  end if;
                when Q_WAIT6622 =>
                  \$v6623\ := \$ram_lock\;
                  if \$v6623\(0) = '1' then
                    state_var7461 := Q_WAIT6622;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(\$17520_copy_root_in_ram6635893_arg\(0 to 15)));
                    state_var7461 := PAUSE_GET6621;
                  end if;
                when Q_WAIT6626 =>
                  \$v6627\ := \$global_end_lock\;
                  if \$v6627\(0) = '1' then
                    state_var7461 := Q_WAIT6626;
                  else
                    acquire(\$global_end_lock\);
                    \$global_end_ptr\ <= 0;
                    state_var7461 := PAUSE_GET6625;
                  end if;
                when Q_WAIT6629 =>
                  \$v6630\ := \$ram_lock\;
                  if \$v6630\(0) = '1' then
                    state_var7461 := Q_WAIT6629;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17761_copy_root_in_ram6635891_arg\(0 to 15)));
                    \$ram_write\ <= \$17780\(0 to 31); \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6628;
                  end if;
                when Q_WAIT6632 =>
                  \$v6633\ := \$ram_lock\;
                  if \$v6633\(0) = '1' then
                    state_var7461 := Q_WAIT6632;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$17776\(0 to 30),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$17761_copy_root_in_ram6635891_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6631;
                  end if;
                when Q_WAIT6635 =>
                  \$v6636\ := \$ram_lock\;
                  if \$v6636\(0) = '1' then
                    state_var7461 := Q_WAIT6635;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$17776\(0 to 30),16)));
                    \$ram_write\ <= eclat_resize(\$17761_copy_root_in_ram6635891_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6634;
                  end if;
                when Q_WAIT6638 =>
                  \$v6639\ := \$ram_lock\;
                  if \$v6639\(0) = '1' then
                    state_var7461 := Q_WAIT6638;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17761_copy_root_in_ram6635891_arg\(32 to 47)));
                    \$ram_write\ <= \$17799_hd\; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6637;
                  end if;
                when Q_WAIT6641 =>
                  \$v6642\ := \$ram_lock\;
                  if \$v6642\(0) = '1' then
                    state_var7461 := Q_WAIT6641;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$17776\(0 to 30),16)));
                    state_var7461 := PAUSE_GET6640;
                  end if;
                when Q_WAIT6645 =>
                  \$v6646\ := \$ram_lock\;
                  if \$v6646\(0) = '1' then
                    state_var7461 := Q_WAIT6645;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$17776\(0 to 30),16), X"000" & X"1")));
                    state_var7461 := PAUSE_GET6644;
                  end if;
                when Q_WAIT6649 =>
                  \$v6650\ := \$ram_lock\;
                  if \$v6650\(0) = '1' then
                    state_var7461 := Q_WAIT6649;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(\$17761_copy_root_in_ram6635891_arg\(0 to 15)));
                    state_var7461 := PAUSE_GET6648;
                  end if;
                when Q_WAIT6653 =>
                  \$v6654\ := \$ram_lock\;
                  if \$v6654\(0) = '1' then
                    state_var7461 := Q_WAIT6653;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17734_copy_root_in_ram6635892_arg\(0 to 15)));
                    \$ram_write\ <= \$17753\(0 to 31); \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6652;
                  end if;
                when Q_WAIT6656 =>
                  \$v6657\ := \$ram_lock\;
                  if \$v6657\(0) = '1' then
                    state_var7461 := Q_WAIT6656;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$17749\(0 to 30),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$17734_copy_root_in_ram6635892_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6655;
                  end if;
                when Q_WAIT6659 =>
                  \$v6660\ := \$ram_lock\;
                  if \$v6660\(0) = '1' then
                    state_var7461 := Q_WAIT6659;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$17749\(0 to 30),16)));
                    \$ram_write\ <= eclat_resize(\$17734_copy_root_in_ram6635892_arg\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6658;
                  end if;
                when Q_WAIT6662 =>
                  \$v6663\ := \$ram_lock\;
                  if \$v6663\(0) = '1' then
                    state_var7461 := Q_WAIT6662;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17734_copy_root_in_ram6635892_arg\(32 to 47)));
                    \$ram_write\ <= \$17879_hd\; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6661;
                  end if;
                when Q_WAIT6665 =>
                  \$v6666\ := \$ram_lock\;
                  if \$v6666\(0) = '1' then
                    state_var7461 := Q_WAIT6665;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$17749\(0 to 30),16)));
                    state_var7461 := PAUSE_GET6664;
                  end if;
                when Q_WAIT6669 =>
                  \$v6670\ := \$ram_lock\;
                  if \$v6670\(0) = '1' then
                    state_var7461 := Q_WAIT6669;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$17749\(0 to 30),16), X"000" & X"1")));
                    state_var7461 := PAUSE_GET6668;
                  end if;
                when Q_WAIT6673 =>
                  \$v6674\ := \$ram_lock\;
                  if \$v6674\(0) = '1' then
                    state_var7461 := Q_WAIT6673;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(\$17734_copy_root_in_ram6635892_arg\(0 to 15)));
                    state_var7461 := PAUSE_GET6672;
                  end if;
                when Q_WAIT6677 =>
                  \$v6678\ := \$ram_lock\;
                  if \$v6678\(0) = '1' then
                    state_var7461 := Q_WAIT6677;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$13922_wait662_arg\(33 to 63),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$17470\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6676;
                  end if;
                when Q_WAIT6680 =>
                  \$v6681\ := \$ram_lock\;
                  if \$v6681\(0) = '1' then
                    state_var7461 := Q_WAIT6680;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$13922_wait662_arg\(33 to 63),16)));
                    \$ram_write\ <= eclat_resize(\$17470\(32 to 47),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6679;
                  end if;
                when Q_WAIT6683 =>
                  \$v6684\ := \$ram_lock\;
                  if \$v6684\(0) = '1' then
                    state_var7461 := Q_WAIT6683;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17470\(32 to 47)));
                    \$ram_write\ <= \$17957_hd\; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6682;
                  end if;
                when Q_WAIT6686 =>
                  \$v6687\ := \$ram_lock\;
                  if \$v6687\(0) = '1' then
                    state_var7461 := Q_WAIT6686;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$13922_wait662_arg\(33 to 63),16)));
                    state_var7461 := PAUSE_GET6685;
                  end if;
                when Q_WAIT6690 =>
                  \$v6691\ := \$ram_lock\;
                  if \$v6691\(0) = '1' then
                    state_var7461 := Q_WAIT6690;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$13922_wait662_arg\(33 to 63),16), X"000" & X"1")));
                    state_var7461 := PAUSE_GET6689;
                  end if;
                when Q_WAIT6694 =>
                  \$v6695\ := \$ram_lock\;
                  if \$v6695\(0) = '1' then
                    state_var7461 := Q_WAIT6694;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$13922_wait662_arg\(1 to 31),16), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(\$17444\(112 to 127),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6693;
                  end if;
                when Q_WAIT6697 =>
                  \$v6698\ := \$ram_lock\;
                  if \$v6698\(0) = '1' then
                    state_var7461 := Q_WAIT6697;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$13922_wait662_arg\(1 to 31),16)));
                    \$ram_write\ <= eclat_resize(\$17444\(112 to 127),31) & eclat_false; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6696;
                  end if;
                when Q_WAIT6700 =>
                  \$v6701\ := \$ram_lock\;
                  if \$v6701\(0) = '1' then
                    state_var7461 := Q_WAIT6700;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17444\(112 to 127)));
                    \$ram_write\ <= \$18035_hd\; \$ram_write_request\ <= '1';
                    state_var7461 := PAUSE_SET6699;
                  end if;
                when Q_WAIT6703 =>
                  \$v6704\ := \$ram_lock\;
                  if \$v6704\(0) = '1' then
                    state_var7461 := Q_WAIT6703;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$13922_wait662_arg\(1 to 31),16)));
                    state_var7461 := PAUSE_GET6702;
                  end if;
                when Q_WAIT6707 =>
                  \$v6708\ := \$ram_lock\;
                  if \$v6708\(0) = '1' then
                    state_var7461 := Q_WAIT6707;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$13922_wait662_arg\(1 to 31),16), X"000" & X"1")));
                    state_var7461 := PAUSE_GET6706;
                  end if;
                when IDLE6505 =>
                  rdy6504 := eclat_false;
                  \$v6710\ := work.Int.gt(work.Int.add(\$17444\(80 to 95), \$13922_wait662_arg\(81 to 96)), 
                                          work.Int.add(\$17444\(96 to 111), X"1770"));
                  if \$v6710\(0) = '1' then
                    \$17463\ := work.Print.print_newline(clk,eclat_unit);
                    \$17464\ := work.Print.print_newline(clk,eclat_unit);
                    \$17465\ := work.Print.print_string(clk,of_string("[================= GC START ======================]"));
                    \$18104\ := work.Print.print_newline(clk,eclat_unit);
                    \$17466\ := work.Print.print_newline(clk,eclat_unit);
                    \$v6709\ := work.Bool.lnot(eclat_if(work.Bool.lnot(
                                                        ""&\$13922_wait662_arg\(32)) & 
                                               eclat_if(work.Int.le(\$17444\(96 to 111), eclat_resize(\$13922_wait662_arg\(1 to 31),16)) & 
                                               work.Int.lt(eclat_resize(\$13922_wait662_arg\(1 to 31),16), 
                                                           work.Int.add(
                                                           \$17444\(96 to 111), X"1770")) & eclat_false) & eclat_false));
                    if \$v6709\(0) = '1' then
                      \$17470\ := \$13922_wait662_arg\(1 to 32) & \$17444\(112 to 127);
                      \$v6692\ := work.Bool.lnot(eclat_if(work.Bool.lnot(
                                                          ""&\$13922_wait662_arg\(64)) & 
                                                 eclat_if(work.Int.le(
                                                          \$17444\(96 to 111), eclat_resize(\$13922_wait662_arg\(33 to 63),16)) & 
                                                 work.Int.lt(eclat_resize(\$13922_wait662_arg\(33 to 63),16), 
                                                             work.Int.add(
                                                             \$17444\(96 to 111), X"1770")) & eclat_false) & eclat_false));
                      if \$v6692\(0) = '1' then
                        \$17487\ := \$13922_wait662_arg\(33 to 64) & \$17470\(32 to 47);
                        \$17734_copy_root_in_ram6635892_id\ := "000000110000";
                        \$17734_copy_root_in_ram6635892_arg\ := X"0" & X"3e8" & \$13922_wait662_arg\(65 to 80) & \$17487\(32 to 47) & \$17444\(96 to 111) & \$17444\(112 to 127);
                        state_var7461 := \$17734_COPY_ROOT_IN_RAM6635892\;
                      else
                        \$v6691\ := \$ram_lock\;
                        if \$v6691\(0) = '1' then
                          state_var7461 := Q_WAIT6690;
                        else
                          acquire(\$ram_lock\);
                          \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                            eclat_resize(\$13922_wait662_arg\(33 to 63),16), X"000" & X"1")));
                          state_var7461 := PAUSE_GET6689;
                        end if;
                      end if;
                    else
                      \$v6708\ := \$ram_lock\;
                      if \$v6708\(0) = '1' then
                        state_var7461 := Q_WAIT6707;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$13922_wait662_arg\(1 to 31),16), X"000" & X"1")));
                        state_var7461 := PAUSE_GET6706;
                      end if;
                    end if;
                  else
                    result6503 := \$13922_wait662_arg\(1 to 32) & \$13922_wait662_arg\(33 to 64) & \$17444\(80 to 95) & 
                    work.Int.add(\$17444\(80 to 95), \$13922_wait662_arg\(81 to 96)) & \$17444\(96 to 111) & \$17444\(112 to 127);
                    rdy6504 := eclat_true;
                    state_var7461 := IDLE6505;
                  end if;
                end case;
                
                if rdy6504(0) = '1' then
                  
                else
                  result6503 := \$17444\(0 to 31) & \$17444\(32 to 63) & \$17444\(64 to 79) & \$17444\(80 to 95) & \$17444\(96 to 111) & \$17444\(112 to 127);
                end if;
                \$17444\ := result6503 & rdy6504;
                \$17434\ := \$17444\;
                \$v6502\ := ""&\$17434\(128);
                if \$v6502\(0) = '1' then
                  \$13922_wait662_result\ := \$17434\(0 to 31) & \$17434\(32 to 63) & \$17434\(64 to 79);
                  \$17389\ := \$13922_wait662_result\;
                  \$17393\ := work.Print.print_string(clk,of_string("size:"));
                  \$17394\ := work.Int.print(clk,eclat_if(work.Int.eq(
                                                          \$13923_make_block579_arg\(88 to 103), X"000" & X"0") & X"000" & X"1" & \$13923_make_block579_arg\(88 to 103)));
                  \$17395\ := work.Print.print_newline(clk,eclat_unit);
                  \$v6714\ := \$ram_lock\;
                  if \$v6714\(0) = '1' then
                    state_var7460 := Q_WAIT6713;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17389\(64 to 79)));
                    \$ram_write\ <= work.Int.lor(work.Int.lsl(eclat_resize(\$13923_make_block579_arg\(80 to 87),31), X"000000" & X"18"), 
                                                 work.Int.lsl(eclat_resize(
                                                              eclat_if(
                                                              work.Int.eq(
                                                              \$13923_make_block579_arg\(88 to 103), X"000" & X"0") & X"000" & X"1" & \$13923_make_block579_arg\(88 to 103)),31), X"0000000" & X"2")) & eclat_true; \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET6712;
                  end if;
                else
                  \$13922_wait662_arg\ := eclat_unit & \$13922_wait662_arg\(1 to 32) & \$13922_wait662_arg\(33 to 64) & \$13922_wait662_arg\(65 to 80) & \$13922_wait662_arg\(81 to 96);
                  state_var7460 := \$13922_WAIT662\;
                end if;
              when \$13923_MAKE_BLOCK579\ =>
                \$17386\ := work.Print.print_string(clk,of_string("GC-ALLOC:(size="));
                \$17387\ := work.Int.print(clk,work.Int.add(eclat_if(
                                                            work.Int.eq(
                                                            \$13923_make_block579_arg\(88 to 103), X"000" & X"0") & X"000" & X"1" & \$13923_make_block579_arg\(88 to 103)), X"000" & X"1"));
                \$17388\ := work.Print.print_string(clk,of_string(")"));
                \$17412\ := work.Print.print_newline(clk,eclat_unit);
                \$13922_wait662_id\ := "000000110011";
                \$13922_wait662_arg\ := eclat_unit & \$13923_make_block579_arg\(16 to 47) & \$13923_make_block579_arg\(48 to 79) & \$13923_make_block579_arg\(0 to 15) & 
                work.Int.add(eclat_if(work.Int.eq(\$13923_make_block579_arg\(88 to 103), X"000" & X"0") & X"000" & X"1" & \$13923_make_block579_arg\(88 to 103)), X"000" & X"1");
                state_var7460 := \$13922_WAIT662\;
              when \$13924_APPLY638\ =>
                \$17310\ := work.Print.print_string(clk,of_string("ENV:"));
                \$17314\ := work.Int.print(clk,\$13924_apply638_arg\(110 to 140));
                \$17315\ := work.Print.print_string(clk,of_string("<"));
                \$v6752\ := ""&\$13924_apply638_arg\(141);
                if \$v6752\(0) = '1' then
                  \$17377\ := work.Print.print_string(clk,of_string("int"));
                  \$17319\ := work.Print.print_string(clk,of_string(">"));
                  \$17320\ := work.Print.print_newline(clk,eclat_unit);
                  \$v6751\ := ""&\$13924_apply638_arg\(0);
                  if \$v6751\(0) = '1' then
                    \$v6750\ := \$ram_lock\;
                    if \$v6750\(0) = '1' then
                      state_var7460 := Q_WAIT6749;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(
                                                        \$13924_apply638_arg\(92 to 107), X"000" & X"1")));
                      state_var7460 := PAUSE_GET6748;
                    end if;
                  else
                    \$17321\ := "000"& X"000000" & X"1" & eclat_true & \$13924_apply638_arg\(92 to 107);
                    \$v6747\ := ""&\$13924_apply638_arg\(1);
                    if \$v6747\(0) = '1' then
                      \$v6746\ := \$ram_lock\;
                      if \$v6746\(0) = '1' then
                        state_var7460 := Q_WAIT6745;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(
                                                          \$17321\(32 to 47), X"000" & X"1")));
                        state_var7460 := PAUSE_GET6744;
                      end if;
                    else
                      \$17324\ := "000"& X"000000" & X"1" & eclat_true & \$17321\(32 to 47);
                      \$v6743\ := ""&\$13924_apply638_arg\(2);
                      if \$v6743\(0) = '1' then
                        \$v6742\ := \$ram_lock\;
                        if \$v6742\(0) = '1' then
                          state_var7460 := Q_WAIT6741;
                        else
                          acquire(\$ram_lock\);
                          \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(
                                                            \$17324\(32 to 47), X"000" & X"1")));
                          state_var7460 := PAUSE_GET6740;
                        end if;
                      else
                        \$17327\ := "000"& X"000000" & X"1" & eclat_true & \$17324\(32 to 47);
                        \$v6739\ := ""&\$13924_apply638_arg\(11);
                        if \$v6739\(0) = '1' then
                          \$17330_sp\ := work.Int.add(work.Int.sub(\$17327\(32 to 47), \$13924_apply638_arg\(12 to 27)), \$13924_apply638_arg\(28 to 43));
                          \$v6729\ := ""&\$13924_apply638_arg\(2);
                          if \$v6729\(0) = '1' then
                            \$v6728\ := \$ram_lock\;
                            if \$v6728\(0) = '1' then
                              state_var7460 := Q_WAIT6727;
                            else
                              acquire(\$ram_lock\);
                              \$ram_ptr_write\ <= to_integer(unsigned(\$17330_sp\));
                              \$ram_write\ <= \$17327\(0 to 31); \$ram_write_request\ <= '1';
                              state_var7460 := PAUSE_SET6726;
                            end if;
                          else
                            \$17331_sp\ := \$17330_sp\;
                            \$v6725\ := ""&\$13924_apply638_arg\(1);
                            if \$v6725\(0) = '1' then
                              \$v6724\ := \$ram_lock\;
                              if \$v6724\(0) = '1' then
                                state_var7460 := Q_WAIT6723;
                              else
                                acquire(\$ram_lock\);
                                \$ram_ptr_write\ <= to_integer(unsigned(\$17331_sp\));
                                \$ram_write\ <= \$17324\(0 to 31); \$ram_write_request\ <= '1';
                                state_var7460 := PAUSE_SET6722;
                              end if;
                            else
                              \$17332_sp\ := \$17331_sp\;
                              \$v6721\ := ""&\$13924_apply638_arg\(0);
                              if \$v6721\(0) = '1' then
                                \$v6720\ := \$ram_lock\;
                                if \$v6720\(0) = '1' then
                                  state_var7460 := Q_WAIT6719;
                                else
                                  acquire(\$ram_lock\);
                                  \$ram_ptr_write\ <= to_integer(unsigned(\$17332_sp\));
                                  \$ram_write\ <= \$17321\(0 to 31); \$ram_write_request\ <= '1';
                                  state_var7460 := PAUSE_SET6718;
                                end if;
                              else
                                \$17333_sp\ := \$17332_sp\;
                                \$v6717\ := \$ram_lock\;
                                if \$v6717\(0) = '1' then
                                  state_var7460 := Q_WAIT6716;
                                else
                                  acquire(\$ram_lock\);
                                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                                    work.Int.add(
                                                                    eclat_resize(\$13924_apply638_arg\(60 to 90),16), X"000" & X"0"), X"000" & X"1")));
                                  state_var7460 := PAUSE_GET6715;
                                end if;
                              end if;
                            end if;
                          end if;
                        else
                          \$v6738\ := \$ram_lock\;
                          if \$v6738\(0) = '1' then
                            state_var7460 := Q_WAIT6737;
                          else
                            acquire(\$ram_lock\);
                            \$ram_ptr_write\ <= to_integer(unsigned(\$17327\(32 to 47)));
                            \$ram_write\ <= eclat_resize(\$13924_apply638_arg\(142 to 149),31) & eclat_true; \$ram_write_request\ <= '1';
                            state_var7460 := PAUSE_SET6736;
                          end if;
                        end if;
                      end if;
                    end if;
                  end if;
                else
                  \$17377\ := work.Print.print_string(clk,of_string("ptr"));
                  \$17319\ := work.Print.print_string(clk,of_string(">"));
                  \$17320\ := work.Print.print_newline(clk,eclat_unit);
                  \$v6751\ := ""&\$13924_apply638_arg\(0);
                  if \$v6751\(0) = '1' then
                    \$v6750\ := \$ram_lock\;
                    if \$v6750\(0) = '1' then
                      state_var7460 := Q_WAIT6749;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(
                                                        \$13924_apply638_arg\(92 to 107), X"000" & X"1")));
                      state_var7460 := PAUSE_GET6748;
                    end if;
                  else
                    \$17321\ := "000"& X"000000" & X"1" & eclat_true & \$13924_apply638_arg\(92 to 107);
                    \$v6747\ := ""&\$13924_apply638_arg\(1);
                    if \$v6747\(0) = '1' then
                      \$v6746\ := \$ram_lock\;
                      if \$v6746\(0) = '1' then
                        state_var7460 := Q_WAIT6745;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(
                                                          \$17321\(32 to 47), X"000" & X"1")));
                        state_var7460 := PAUSE_GET6744;
                      end if;
                    else
                      \$17324\ := "000"& X"000000" & X"1" & eclat_true & \$17321\(32 to 47);
                      \$v6743\ := ""&\$13924_apply638_arg\(2);
                      if \$v6743\(0) = '1' then
                        \$v6742\ := \$ram_lock\;
                        if \$v6742\(0) = '1' then
                          state_var7460 := Q_WAIT6741;
                        else
                          acquire(\$ram_lock\);
                          \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(
                                                            \$17324\(32 to 47), X"000" & X"1")));
                          state_var7460 := PAUSE_GET6740;
                        end if;
                      else
                        \$17327\ := "000"& X"000000" & X"1" & eclat_true & \$17324\(32 to 47);
                        \$v6739\ := ""&\$13924_apply638_arg\(11);
                        if \$v6739\(0) = '1' then
                          \$17330_sp\ := work.Int.add(work.Int.sub(\$17327\(32 to 47), \$13924_apply638_arg\(12 to 27)), \$13924_apply638_arg\(28 to 43));
                          \$v6729\ := ""&\$13924_apply638_arg\(2);
                          if \$v6729\(0) = '1' then
                            \$v6728\ := \$ram_lock\;
                            if \$v6728\(0) = '1' then
                              state_var7460 := Q_WAIT6727;
                            else
                              acquire(\$ram_lock\);
                              \$ram_ptr_write\ <= to_integer(unsigned(\$17330_sp\));
                              \$ram_write\ <= \$17327\(0 to 31); \$ram_write_request\ <= '1';
                              state_var7460 := PAUSE_SET6726;
                            end if;
                          else
                            \$17331_sp\ := \$17330_sp\;
                            \$v6725\ := ""&\$13924_apply638_arg\(1);
                            if \$v6725\(0) = '1' then
                              \$v6724\ := \$ram_lock\;
                              if \$v6724\(0) = '1' then
                                state_var7460 := Q_WAIT6723;
                              else
                                acquire(\$ram_lock\);
                                \$ram_ptr_write\ <= to_integer(unsigned(\$17331_sp\));
                                \$ram_write\ <= \$17324\(0 to 31); \$ram_write_request\ <= '1';
                                state_var7460 := PAUSE_SET6722;
                              end if;
                            else
                              \$17332_sp\ := \$17331_sp\;
                              \$v6721\ := ""&\$13924_apply638_arg\(0);
                              if \$v6721\(0) = '1' then
                                \$v6720\ := \$ram_lock\;
                                if \$v6720\(0) = '1' then
                                  state_var7460 := Q_WAIT6719;
                                else
                                  acquire(\$ram_lock\);
                                  \$ram_ptr_write\ <= to_integer(unsigned(\$17332_sp\));
                                  \$ram_write\ <= \$17321\(0 to 31); \$ram_write_request\ <= '1';
                                  state_var7460 := PAUSE_SET6718;
                                end if;
                              else
                                \$17333_sp\ := \$17332_sp\;
                                \$v6717\ := \$ram_lock\;
                                if \$v6717\(0) = '1' then
                                  state_var7460 := Q_WAIT6716;
                                else
                                  acquire(\$ram_lock\);
                                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                                    work.Int.add(
                                                                    eclat_resize(\$13924_apply638_arg\(60 to 90),16), X"000" & X"0"), X"000" & X"1")));
                                  state_var7460 := PAUSE_GET6715;
                                end if;
                              end if;
                            end if;
                          end if;
                        else
                          \$v6738\ := \$ram_lock\;
                          if \$v6738\(0) = '1' then
                            state_var7460 := Q_WAIT6737;
                          else
                            acquire(\$ram_lock\);
                            \$ram_ptr_write\ <= to_integer(unsigned(\$17327\(32 to 47)));
                            \$ram_write\ <= eclat_resize(\$13924_apply638_arg\(142 to 149),31) & eclat_true; \$ram_write_request\ <= '1';
                            state_var7460 := PAUSE_SET6736;
                          end if;
                        end if;
                      end if;
                    end if;
                  end if;
                end if;
              when \$13925_OFFSETCLOSURE_N639\ =>
                \$13925_offsetclosure_n639_result\ := \$13925_offsetclosure_n639_arg\(0 to 15) & eclat_resize(
                work.Int.add(eclat_resize(\$13925_offsetclosure_n639_arg\(106 to 136),16), \$13925_offsetclosure_n639_arg\(32 to 47)),31) & eclat_false & \$13925_offsetclosure_n639_arg\(16 to 31) & \$13925_offsetclosure_n639_arg\(48 to 103) & \$13925_offsetclosure_n639_arg\(104 to 105);
                result6468 := \$13925_offsetclosure_n639_result\;
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when \$13926_MAKE_BLOCK_N646\ =>
                \$13923_make_block579_id\ := "000000110100";
                \$13923_make_block579_arg\ := \$13926_make_block_n646_arg\(16 to 31) & \$13926_make_block_n646_arg\(82 to 113) & \$13926_make_block_n646_arg\(116 to 147) & eclat_resize(\$13926_make_block_n646_arg\(35 to 65),8) & \$13926_make_block_n646_arg\(66 to 81);
                state_var7460 := \$13923_MAKE_BLOCK579\;
              when \$13927_BRANCH_IF648\ =>
                \$v6774\ := eclat_if(""&\$13927_branch_if648_arg\(0) & 
                            work.Bool.lnot(work.Int.neq(\$13927_branch_if648_arg\(17 to 47), "000"& X"000000" & X"0")) & 
                            work.Int.neq(\$13927_branch_if648_arg\(17 to 47), "000"& X"000000" & X"0"));
                if \$v6774\(0) = '1' then
                  \$v6773\ := \$code_lock\;
                  if \$v6773\(0) = '1' then
                    state_var7460 := Q_WAIT6772;
                  else
                    acquire(\$code_lock\);
                    \$code_ptr\ <= to_integer(unsigned(work.Int.add(\$13927_branch_if648_arg\(1 to 16), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6771;
                  end if;
                else
                  \$13927_branch_if648_result\ := work.Int.add(\$13927_branch_if648_arg\(1 to 16), X"000" & X"2") & \$13927_branch_if648_arg\(17 to 48) & \$13927_branch_if648_arg\(49 to 64) & \$13927_branch_if648_arg\(65 to 120) & \$13927_branch_if648_arg\(121 to 122);
                  result6468 := \$13927_branch_if648_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                end if;
              when \$13928_W652\ =>
                \$v6781\ := work.Int.gt(\$13928_w652_arg\(0 to 15), \$13928_w652_arg\(32 to 47));
                if \$v6781\(0) = '1' then
                  \$13928_w652_result\ := eclat_unit;
                  \$16626\ := \$13928_w652_result\;
                  \$v7358\ := \$ram_lock\;
                  if \$v7358\(0) = '1' then
                    state_var7460 := Q_WAIT7357;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$13911\(16 to 46),16), X"000" & X"0"), X"000" & X"1")));
                    state_var7460 := PAUSE_GET7356;
                  end if;
                else
                  \$v6780\ := \$ram_lock\;
                  if \$v6780\(0) = '1' then
                    state_var7460 := Q_WAIT6779;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13928_w652_arg\(16 to 31), \$13928_w652_arg\(0 to 15))));
                    state_var7460 := PAUSE_GET6778;
                  end if;
                end if;
              when \$14207_LOOP_PUSH6495899\ =>
                \$v6899\ := work.Int.ge(\$14207_loop_push6495899_arg\(16 to 23), 
                                        work.Int.sub(\$14207_loop_push6495899_arg\(56 to 63), "00000010"));
                if \$v6899\(0) = '1' then
                  \$14207_loop_push6495899_result\ := \$14207_loop_push6495899_arg\(0 to 15);
                  \$14181_sp\ := \$14207_loop_push6495899_result\;
                  \$v6892\ := \$ram_lock\;
                  if \$v6892\(0) = '1' then
                    state_var7460 := Q_WAIT6891;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$13911\(64 to 94),16), X"000" & X"1"), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6890;
                  end if;
                else
                  \$v6898\ := \$ram_lock\;
                  if \$v6898\(0) = '1' then
                    state_var7460 := Q_WAIT6897;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$14207_loop_push6495899_arg\(24 to 54),16), eclat_resize(
                                                                   work.Int.add(
                                                                   \$14207_loop_push6495899_arg\(16 to 23), "00000010"),16)), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6896;
                  end if;
                end if;
              when \$14564_BINOP_INT6435900\ =>
                \$v7020\ := \$ram_lock\;
                if \$v7020\(0) = '1' then
                  state_var7460 := Q_WAIT7019;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$14564_binop_int6435900_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7018;
                end if;
              when \$14589_MODULO6685895\ =>
                \$v7012\ := work.Int.lt(\$14589_modulo6685895_arg\(0 to 30), \$14589_modulo6685895_arg\(31 to 61));
                if \$v7012\(0) = '1' then
                  \$14589_modulo6685895_result\ := \$14589_modulo6685895_arg\(0 to 30);
                  \$14586_r\ := \$14589_modulo6685895_result\;
                  \$14582_res\ := eclat_if(work.Int.lt(\$14564_binop_int6435900_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$14586_r\) & \$14586_r\);
                  \$14564_binop_int6435900_result\ := work.Int.add(\$14564_binop_int6435900_arg\(32 to 47), X"000" & X"1") & \$14582_res\ & eclat_true & 
                  work.Int.sub(\$14564_binop_int6435900_arg\(80 to 95), X"000" & X"1") & \$14564_binop_int6435900_arg\(96 to 151) & \$14564_binop_int6435900_arg\(152 to 153);
                  result6468 := \$14564_binop_int6435900_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$14597_modulo6685888_id\ := "000001000011";
                  \$14597_modulo6685888_arg\ := work.Int.sub(\$14589_modulo6685895_arg\(0 to 30), \$14589_modulo6685895_arg\(31 to 61)) & \$14589_modulo6685895_arg\(31 to 61);
                  state_var7460 := \$14597_MODULO6685888\;
                end if;
              when \$14597_MODULO6685888\ =>
                \$v7011\ := work.Int.lt(\$14597_modulo6685888_arg\(0 to 30), \$14597_modulo6685888_arg\(31 to 61));
                if \$v7011\(0) = '1' then
                  \$14597_modulo6685888_result\ := \$14597_modulo6685888_arg\(0 to 30);
                  \$14589_modulo6685895_result\ := \$14597_modulo6685888_result\;
                  \$14586_r\ := \$14589_modulo6685895_result\;
                  \$14582_res\ := eclat_if(work.Int.lt(\$14564_binop_int6435900_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$14586_r\) & \$14586_r\);
                  \$14564_binop_int6435900_result\ := work.Int.add(\$14564_binop_int6435900_arg\(32 to 47), X"000" & X"1") & \$14582_res\ & eclat_true & 
                  work.Int.sub(\$14564_binop_int6435900_arg\(80 to 95), X"000" & X"1") & \$14564_binop_int6435900_arg\(96 to 151) & \$14564_binop_int6435900_arg\(152 to 153);
                  result6468 := \$14564_binop_int6435900_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$14597_modulo6685888_arg\ := work.Int.sub(\$14597_modulo6685888_arg\(0 to 30), \$14597_modulo6685888_arg\(31 to 61)) & \$14597_modulo6685888_arg\(31 to 61);
                  state_var7460 := \$14597_MODULO6685888\;
                end if;
              when \$14613_MODULO6685896\ =>
                \$v7015\ := work.Int.lt(\$14613_modulo6685896_arg\(0 to 30), \$14613_modulo6685896_arg\(31 to 61));
                if \$v7015\(0) = '1' then
                  \$14613_modulo6685896_result\ := \$14613_modulo6685896_arg\(0 to 30);
                  \$14610_r\ := \$14613_modulo6685896_result\;
                  \$14582_res\ := eclat_if(work.Int.lt(\$14564_binop_int6435900_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$14610_r\) & \$14610_r\);
                  \$14564_binop_int6435900_result\ := work.Int.add(\$14564_binop_int6435900_arg\(32 to 47), X"000" & X"1") & \$14582_res\ & eclat_true & 
                  work.Int.sub(\$14564_binop_int6435900_arg\(80 to 95), X"000" & X"1") & \$14564_binop_int6435900_arg\(96 to 151) & \$14564_binop_int6435900_arg\(152 to 153);
                  result6468 := \$14564_binop_int6435900_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$14621_modulo6685888_id\ := "000001000101";
                  \$14621_modulo6685888_arg\ := work.Int.sub(\$14613_modulo6685896_arg\(0 to 30), \$14613_modulo6685896_arg\(31 to 61)) & \$14613_modulo6685896_arg\(31 to 61);
                  state_var7460 := \$14621_MODULO6685888\;
                end if;
              when \$14621_MODULO6685888\ =>
                \$v7014\ := work.Int.lt(\$14621_modulo6685888_arg\(0 to 30), \$14621_modulo6685888_arg\(31 to 61));
                if \$v7014\(0) = '1' then
                  \$14621_modulo6685888_result\ := \$14621_modulo6685888_arg\(0 to 30);
                  \$14613_modulo6685896_result\ := \$14621_modulo6685888_result\;
                  \$14610_r\ := \$14613_modulo6685896_result\;
                  \$14582_res\ := eclat_if(work.Int.lt(\$14564_binop_int6435900_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$14610_r\) & \$14610_r\);
                  \$14564_binop_int6435900_result\ := work.Int.add(\$14564_binop_int6435900_arg\(32 to 47), X"000" & X"1") & \$14582_res\ & eclat_true & 
                  work.Int.sub(\$14564_binop_int6435900_arg\(80 to 95), X"000" & X"1") & \$14564_binop_int6435900_arg\(96 to 151) & \$14564_binop_int6435900_arg\(152 to 153);
                  result6468 := \$14564_binop_int6435900_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$14621_modulo6685888_arg\ := work.Int.sub(\$14621_modulo6685888_arg\(0 to 30), \$14621_modulo6685888_arg\(31 to 61)) & \$14621_modulo6685888_arg\(31 to 61);
                  state_var7460 := \$14621_MODULO6685888\;
                end if;
              when \$14644_BINOP_INT6435901\ =>
                \$v7030\ := \$ram_lock\;
                if \$v7030\(0) = '1' then
                  state_var7460 := Q_WAIT7029;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$14644_binop_int6435901_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7028;
                end if;
              when \$14669_MODULO6685895\ =>
                \$v7022\ := work.Int.lt(\$14669_modulo6685895_arg\(0 to 30), \$14669_modulo6685895_arg\(31 to 61));
                if \$v7022\(0) = '1' then
                  \$14669_modulo6685895_result\ := \$14669_modulo6685895_arg\(0 to 30);
                  \$14666_r\ := \$14669_modulo6685895_result\;
                  \$14662_res\ := eclat_if(work.Int.lt(\$14644_binop_int6435901_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$14666_r\) & \$14666_r\);
                  \$14644_binop_int6435901_result\ := work.Int.add(\$14644_binop_int6435901_arg\(32 to 47), X"000" & X"1") & \$14662_res\ & eclat_true & 
                  work.Int.sub(\$14644_binop_int6435901_arg\(80 to 95), X"000" & X"1") & \$14644_binop_int6435901_arg\(96 to 151) & \$14644_binop_int6435901_arg\(152 to 153);
                  result6468 := \$14644_binop_int6435901_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$14677_modulo6685888_id\ := "000001001000";
                  \$14677_modulo6685888_arg\ := work.Int.sub(\$14669_modulo6685895_arg\(0 to 30), \$14669_modulo6685895_arg\(31 to 61)) & \$14669_modulo6685895_arg\(31 to 61);
                  state_var7460 := \$14677_MODULO6685888\;
                end if;
              when \$14677_MODULO6685888\ =>
                \$v7021\ := work.Int.lt(\$14677_modulo6685888_arg\(0 to 30), \$14677_modulo6685888_arg\(31 to 61));
                if \$v7021\(0) = '1' then
                  \$14677_modulo6685888_result\ := \$14677_modulo6685888_arg\(0 to 30);
                  \$14669_modulo6685895_result\ := \$14677_modulo6685888_result\;
                  \$14666_r\ := \$14669_modulo6685895_result\;
                  \$14662_res\ := eclat_if(work.Int.lt(\$14644_binop_int6435901_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$14666_r\) & \$14666_r\);
                  \$14644_binop_int6435901_result\ := work.Int.add(\$14644_binop_int6435901_arg\(32 to 47), X"000" & X"1") & \$14662_res\ & eclat_true & 
                  work.Int.sub(\$14644_binop_int6435901_arg\(80 to 95), X"000" & X"1") & \$14644_binop_int6435901_arg\(96 to 151) & \$14644_binop_int6435901_arg\(152 to 153);
                  result6468 := \$14644_binop_int6435901_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$14677_modulo6685888_arg\ := work.Int.sub(\$14677_modulo6685888_arg\(0 to 30), \$14677_modulo6685888_arg\(31 to 61)) & \$14677_modulo6685888_arg\(31 to 61);
                  state_var7460 := \$14677_MODULO6685888\;
                end if;
              when \$14693_MODULO6685896\ =>
                \$v7025\ := work.Int.lt(\$14693_modulo6685896_arg\(0 to 30), \$14693_modulo6685896_arg\(31 to 61));
                if \$v7025\(0) = '1' then
                  \$14693_modulo6685896_result\ := \$14693_modulo6685896_arg\(0 to 30);
                  \$14690_r\ := \$14693_modulo6685896_result\;
                  \$14662_res\ := eclat_if(work.Int.lt(\$14644_binop_int6435901_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$14690_r\) & \$14690_r\);
                  \$14644_binop_int6435901_result\ := work.Int.add(\$14644_binop_int6435901_arg\(32 to 47), X"000" & X"1") & \$14662_res\ & eclat_true & 
                  work.Int.sub(\$14644_binop_int6435901_arg\(80 to 95), X"000" & X"1") & \$14644_binop_int6435901_arg\(96 to 151) & \$14644_binop_int6435901_arg\(152 to 153);
                  result6468 := \$14644_binop_int6435901_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$14701_modulo6685888_id\ := "000001001010";
                  \$14701_modulo6685888_arg\ := work.Int.sub(\$14693_modulo6685896_arg\(0 to 30), \$14693_modulo6685896_arg\(31 to 61)) & \$14693_modulo6685896_arg\(31 to 61);
                  state_var7460 := \$14701_MODULO6685888\;
                end if;
              when \$14701_MODULO6685888\ =>
                \$v7024\ := work.Int.lt(\$14701_modulo6685888_arg\(0 to 30), \$14701_modulo6685888_arg\(31 to 61));
                if \$v7024\(0) = '1' then
                  \$14701_modulo6685888_result\ := \$14701_modulo6685888_arg\(0 to 30);
                  \$14693_modulo6685896_result\ := \$14701_modulo6685888_result\;
                  \$14690_r\ := \$14693_modulo6685896_result\;
                  \$14662_res\ := eclat_if(work.Int.lt(\$14644_binop_int6435901_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$14690_r\) & \$14690_r\);
                  \$14644_binop_int6435901_result\ := work.Int.add(\$14644_binop_int6435901_arg\(32 to 47), X"000" & X"1") & \$14662_res\ & eclat_true & 
                  work.Int.sub(\$14644_binop_int6435901_arg\(80 to 95), X"000" & X"1") & \$14644_binop_int6435901_arg\(96 to 151) & \$14644_binop_int6435901_arg\(152 to 153);
                  result6468 := \$14644_binop_int6435901_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$14701_modulo6685888_arg\ := work.Int.sub(\$14701_modulo6685888_arg\(0 to 30), \$14701_modulo6685888_arg\(31 to 61)) & \$14701_modulo6685888_arg\(31 to 61);
                  state_var7460 := \$14701_MODULO6685888\;
                end if;
              when \$14724_BINOP_INT6435902\ =>
                \$v7040\ := \$ram_lock\;
                if \$v7040\(0) = '1' then
                  state_var7460 := Q_WAIT7039;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$14724_binop_int6435902_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7038;
                end if;
              when \$14749_MODULO6685895\ =>
                \$v7032\ := work.Int.lt(\$14749_modulo6685895_arg\(0 to 30), \$14749_modulo6685895_arg\(31 to 61));
                if \$v7032\(0) = '1' then
                  \$14749_modulo6685895_result\ := \$14749_modulo6685895_arg\(0 to 30);
                  \$14746_r\ := \$14749_modulo6685895_result\;
                  \$14742_res\ := eclat_if(work.Int.lt(\$14724_binop_int6435902_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$14746_r\) & \$14746_r\);
                  \$14724_binop_int6435902_result\ := work.Int.add(\$14724_binop_int6435902_arg\(32 to 47), X"000" & X"1") & \$14742_res\ & eclat_true & 
                  work.Int.sub(\$14724_binop_int6435902_arg\(80 to 95), X"000" & X"1") & \$14724_binop_int6435902_arg\(96 to 151) & \$14724_binop_int6435902_arg\(152 to 153);
                  result6468 := \$14724_binop_int6435902_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$14757_modulo6685888_id\ := "000001001101";
                  \$14757_modulo6685888_arg\ := work.Int.sub(\$14749_modulo6685895_arg\(0 to 30), \$14749_modulo6685895_arg\(31 to 61)) & \$14749_modulo6685895_arg\(31 to 61);
                  state_var7460 := \$14757_MODULO6685888\;
                end if;
              when \$14757_MODULO6685888\ =>
                \$v7031\ := work.Int.lt(\$14757_modulo6685888_arg\(0 to 30), \$14757_modulo6685888_arg\(31 to 61));
                if \$v7031\(0) = '1' then
                  \$14757_modulo6685888_result\ := \$14757_modulo6685888_arg\(0 to 30);
                  \$14749_modulo6685895_result\ := \$14757_modulo6685888_result\;
                  \$14746_r\ := \$14749_modulo6685895_result\;
                  \$14742_res\ := eclat_if(work.Int.lt(\$14724_binop_int6435902_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$14746_r\) & \$14746_r\);
                  \$14724_binop_int6435902_result\ := work.Int.add(\$14724_binop_int6435902_arg\(32 to 47), X"000" & X"1") & \$14742_res\ & eclat_true & 
                  work.Int.sub(\$14724_binop_int6435902_arg\(80 to 95), X"000" & X"1") & \$14724_binop_int6435902_arg\(96 to 151) & \$14724_binop_int6435902_arg\(152 to 153);
                  result6468 := \$14724_binop_int6435902_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$14757_modulo6685888_arg\ := work.Int.sub(\$14757_modulo6685888_arg\(0 to 30), \$14757_modulo6685888_arg\(31 to 61)) & \$14757_modulo6685888_arg\(31 to 61);
                  state_var7460 := \$14757_MODULO6685888\;
                end if;
              when \$14773_MODULO6685896\ =>
                \$v7035\ := work.Int.lt(\$14773_modulo6685896_arg\(0 to 30), \$14773_modulo6685896_arg\(31 to 61));
                if \$v7035\(0) = '1' then
                  \$14773_modulo6685896_result\ := \$14773_modulo6685896_arg\(0 to 30);
                  \$14770_r\ := \$14773_modulo6685896_result\;
                  \$14742_res\ := eclat_if(work.Int.lt(\$14724_binop_int6435902_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$14770_r\) & \$14770_r\);
                  \$14724_binop_int6435902_result\ := work.Int.add(\$14724_binop_int6435902_arg\(32 to 47), X"000" & X"1") & \$14742_res\ & eclat_true & 
                  work.Int.sub(\$14724_binop_int6435902_arg\(80 to 95), X"000" & X"1") & \$14724_binop_int6435902_arg\(96 to 151) & \$14724_binop_int6435902_arg\(152 to 153);
                  result6468 := \$14724_binop_int6435902_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$14781_modulo6685888_id\ := "000001001111";
                  \$14781_modulo6685888_arg\ := work.Int.sub(\$14773_modulo6685896_arg\(0 to 30), \$14773_modulo6685896_arg\(31 to 61)) & \$14773_modulo6685896_arg\(31 to 61);
                  state_var7460 := \$14781_MODULO6685888\;
                end if;
              when \$14781_MODULO6685888\ =>
                \$v7034\ := work.Int.lt(\$14781_modulo6685888_arg\(0 to 30), \$14781_modulo6685888_arg\(31 to 61));
                if \$v7034\(0) = '1' then
                  \$14781_modulo6685888_result\ := \$14781_modulo6685888_arg\(0 to 30);
                  \$14773_modulo6685896_result\ := \$14781_modulo6685888_result\;
                  \$14770_r\ := \$14773_modulo6685896_result\;
                  \$14742_res\ := eclat_if(work.Int.lt(\$14724_binop_int6435902_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$14770_r\) & \$14770_r\);
                  \$14724_binop_int6435902_result\ := work.Int.add(\$14724_binop_int6435902_arg\(32 to 47), X"000" & X"1") & \$14742_res\ & eclat_true & 
                  work.Int.sub(\$14724_binop_int6435902_arg\(80 to 95), X"000" & X"1") & \$14724_binop_int6435902_arg\(96 to 151) & \$14724_binop_int6435902_arg\(152 to 153);
                  result6468 := \$14724_binop_int6435902_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$14781_modulo6685888_arg\ := work.Int.sub(\$14781_modulo6685888_arg\(0 to 30), \$14781_modulo6685888_arg\(31 to 61)) & \$14781_modulo6685888_arg\(31 to 61);
                  state_var7460 := \$14781_MODULO6685888\;
                end if;
              when \$14804_BINOP_INT6435903\ =>
                \$v7050\ := \$ram_lock\;
                if \$v7050\(0) = '1' then
                  state_var7460 := Q_WAIT7049;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$14804_binop_int6435903_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7048;
                end if;
              when \$14829_MODULO6685895\ =>
                \$v7042\ := work.Int.lt(\$14829_modulo6685895_arg\(0 to 30), \$14829_modulo6685895_arg\(31 to 61));
                if \$v7042\(0) = '1' then
                  \$14829_modulo6685895_result\ := \$14829_modulo6685895_arg\(0 to 30);
                  \$14826_r\ := \$14829_modulo6685895_result\;
                  \$14822_res\ := eclat_if(work.Int.lt(\$14804_binop_int6435903_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$14826_r\) & \$14826_r\);
                  \$14804_binop_int6435903_result\ := work.Int.add(\$14804_binop_int6435903_arg\(32 to 47), X"000" & X"1") & \$14822_res\ & eclat_true & 
                  work.Int.sub(\$14804_binop_int6435903_arg\(80 to 95), X"000" & X"1") & \$14804_binop_int6435903_arg\(96 to 151) & \$14804_binop_int6435903_arg\(152 to 153);
                  result6468 := \$14804_binop_int6435903_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$14837_modulo6685888_id\ := "000001010010";
                  \$14837_modulo6685888_arg\ := work.Int.sub(\$14829_modulo6685895_arg\(0 to 30), \$14829_modulo6685895_arg\(31 to 61)) & \$14829_modulo6685895_arg\(31 to 61);
                  state_var7460 := \$14837_MODULO6685888\;
                end if;
              when \$14837_MODULO6685888\ =>
                \$v7041\ := work.Int.lt(\$14837_modulo6685888_arg\(0 to 30), \$14837_modulo6685888_arg\(31 to 61));
                if \$v7041\(0) = '1' then
                  \$14837_modulo6685888_result\ := \$14837_modulo6685888_arg\(0 to 30);
                  \$14829_modulo6685895_result\ := \$14837_modulo6685888_result\;
                  \$14826_r\ := \$14829_modulo6685895_result\;
                  \$14822_res\ := eclat_if(work.Int.lt(\$14804_binop_int6435903_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$14826_r\) & \$14826_r\);
                  \$14804_binop_int6435903_result\ := work.Int.add(\$14804_binop_int6435903_arg\(32 to 47), X"000" & X"1") & \$14822_res\ & eclat_true & 
                  work.Int.sub(\$14804_binop_int6435903_arg\(80 to 95), X"000" & X"1") & \$14804_binop_int6435903_arg\(96 to 151) & \$14804_binop_int6435903_arg\(152 to 153);
                  result6468 := \$14804_binop_int6435903_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$14837_modulo6685888_arg\ := work.Int.sub(\$14837_modulo6685888_arg\(0 to 30), \$14837_modulo6685888_arg\(31 to 61)) & \$14837_modulo6685888_arg\(31 to 61);
                  state_var7460 := \$14837_MODULO6685888\;
                end if;
              when \$14853_MODULO6685896\ =>
                \$v7045\ := work.Int.lt(\$14853_modulo6685896_arg\(0 to 30), \$14853_modulo6685896_arg\(31 to 61));
                if \$v7045\(0) = '1' then
                  \$14853_modulo6685896_result\ := \$14853_modulo6685896_arg\(0 to 30);
                  \$14850_r\ := \$14853_modulo6685896_result\;
                  \$14822_res\ := eclat_if(work.Int.lt(\$14804_binop_int6435903_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$14850_r\) & \$14850_r\);
                  \$14804_binop_int6435903_result\ := work.Int.add(\$14804_binop_int6435903_arg\(32 to 47), X"000" & X"1") & \$14822_res\ & eclat_true & 
                  work.Int.sub(\$14804_binop_int6435903_arg\(80 to 95), X"000" & X"1") & \$14804_binop_int6435903_arg\(96 to 151) & \$14804_binop_int6435903_arg\(152 to 153);
                  result6468 := \$14804_binop_int6435903_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$14861_modulo6685888_id\ := "000001010100";
                  \$14861_modulo6685888_arg\ := work.Int.sub(\$14853_modulo6685896_arg\(0 to 30), \$14853_modulo6685896_arg\(31 to 61)) & \$14853_modulo6685896_arg\(31 to 61);
                  state_var7460 := \$14861_MODULO6685888\;
                end if;
              when \$14861_MODULO6685888\ =>
                \$v7044\ := work.Int.lt(\$14861_modulo6685888_arg\(0 to 30), \$14861_modulo6685888_arg\(31 to 61));
                if \$v7044\(0) = '1' then
                  \$14861_modulo6685888_result\ := \$14861_modulo6685888_arg\(0 to 30);
                  \$14853_modulo6685896_result\ := \$14861_modulo6685888_result\;
                  \$14850_r\ := \$14853_modulo6685896_result\;
                  \$14822_res\ := eclat_if(work.Int.lt(\$14804_binop_int6435903_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$14850_r\) & \$14850_r\);
                  \$14804_binop_int6435903_result\ := work.Int.add(\$14804_binop_int6435903_arg\(32 to 47), X"000" & X"1") & \$14822_res\ & eclat_true & 
                  work.Int.sub(\$14804_binop_int6435903_arg\(80 to 95), X"000" & X"1") & \$14804_binop_int6435903_arg\(96 to 151) & \$14804_binop_int6435903_arg\(152 to 153);
                  result6468 := \$14804_binop_int6435903_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$14861_modulo6685888_arg\ := work.Int.sub(\$14861_modulo6685888_arg\(0 to 30), \$14861_modulo6685888_arg\(31 to 61)) & \$14861_modulo6685888_arg\(31 to 61);
                  state_var7460 := \$14861_MODULO6685888\;
                end if;
              when \$14884_BINOP_INT6435904\ =>
                \$v7060\ := \$ram_lock\;
                if \$v7060\(0) = '1' then
                  state_var7460 := Q_WAIT7059;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$14884_binop_int6435904_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7058;
                end if;
              when \$14909_MODULO6685895\ =>
                \$v7052\ := work.Int.lt(\$14909_modulo6685895_arg\(0 to 30), \$14909_modulo6685895_arg\(31 to 61));
                if \$v7052\(0) = '1' then
                  \$14909_modulo6685895_result\ := \$14909_modulo6685895_arg\(0 to 30);
                  \$14906_r\ := \$14909_modulo6685895_result\;
                  \$14902_res\ := eclat_if(work.Int.lt(\$14884_binop_int6435904_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$14906_r\) & \$14906_r\);
                  \$14884_binop_int6435904_result\ := work.Int.add(\$14884_binop_int6435904_arg\(32 to 47), X"000" & X"1") & \$14902_res\ & eclat_true & 
                  work.Int.sub(\$14884_binop_int6435904_arg\(80 to 95), X"000" & X"1") & \$14884_binop_int6435904_arg\(96 to 151) & \$14884_binop_int6435904_arg\(152 to 153);
                  result6468 := \$14884_binop_int6435904_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$14917_modulo6685888_id\ := "000001010111";
                  \$14917_modulo6685888_arg\ := work.Int.sub(\$14909_modulo6685895_arg\(0 to 30), \$14909_modulo6685895_arg\(31 to 61)) & \$14909_modulo6685895_arg\(31 to 61);
                  state_var7460 := \$14917_MODULO6685888\;
                end if;
              when \$14917_MODULO6685888\ =>
                \$v7051\ := work.Int.lt(\$14917_modulo6685888_arg\(0 to 30), \$14917_modulo6685888_arg\(31 to 61));
                if \$v7051\(0) = '1' then
                  \$14917_modulo6685888_result\ := \$14917_modulo6685888_arg\(0 to 30);
                  \$14909_modulo6685895_result\ := \$14917_modulo6685888_result\;
                  \$14906_r\ := \$14909_modulo6685895_result\;
                  \$14902_res\ := eclat_if(work.Int.lt(\$14884_binop_int6435904_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$14906_r\) & \$14906_r\);
                  \$14884_binop_int6435904_result\ := work.Int.add(\$14884_binop_int6435904_arg\(32 to 47), X"000" & X"1") & \$14902_res\ & eclat_true & 
                  work.Int.sub(\$14884_binop_int6435904_arg\(80 to 95), X"000" & X"1") & \$14884_binop_int6435904_arg\(96 to 151) & \$14884_binop_int6435904_arg\(152 to 153);
                  result6468 := \$14884_binop_int6435904_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$14917_modulo6685888_arg\ := work.Int.sub(\$14917_modulo6685888_arg\(0 to 30), \$14917_modulo6685888_arg\(31 to 61)) & \$14917_modulo6685888_arg\(31 to 61);
                  state_var7460 := \$14917_MODULO6685888\;
                end if;
              when \$14933_MODULO6685896\ =>
                \$v7055\ := work.Int.lt(\$14933_modulo6685896_arg\(0 to 30), \$14933_modulo6685896_arg\(31 to 61));
                if \$v7055\(0) = '1' then
                  \$14933_modulo6685896_result\ := \$14933_modulo6685896_arg\(0 to 30);
                  \$14930_r\ := \$14933_modulo6685896_result\;
                  \$14902_res\ := eclat_if(work.Int.lt(\$14884_binop_int6435904_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$14930_r\) & \$14930_r\);
                  \$14884_binop_int6435904_result\ := work.Int.add(\$14884_binop_int6435904_arg\(32 to 47), X"000" & X"1") & \$14902_res\ & eclat_true & 
                  work.Int.sub(\$14884_binop_int6435904_arg\(80 to 95), X"000" & X"1") & \$14884_binop_int6435904_arg\(96 to 151) & \$14884_binop_int6435904_arg\(152 to 153);
                  result6468 := \$14884_binop_int6435904_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$14941_modulo6685888_id\ := "000001011001";
                  \$14941_modulo6685888_arg\ := work.Int.sub(\$14933_modulo6685896_arg\(0 to 30), \$14933_modulo6685896_arg\(31 to 61)) & \$14933_modulo6685896_arg\(31 to 61);
                  state_var7460 := \$14941_MODULO6685888\;
                end if;
              when \$14941_MODULO6685888\ =>
                \$v7054\ := work.Int.lt(\$14941_modulo6685888_arg\(0 to 30), \$14941_modulo6685888_arg\(31 to 61));
                if \$v7054\(0) = '1' then
                  \$14941_modulo6685888_result\ := \$14941_modulo6685888_arg\(0 to 30);
                  \$14933_modulo6685896_result\ := \$14941_modulo6685888_result\;
                  \$14930_r\ := \$14933_modulo6685896_result\;
                  \$14902_res\ := eclat_if(work.Int.lt(\$14884_binop_int6435904_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$14930_r\) & \$14930_r\);
                  \$14884_binop_int6435904_result\ := work.Int.add(\$14884_binop_int6435904_arg\(32 to 47), X"000" & X"1") & \$14902_res\ & eclat_true & 
                  work.Int.sub(\$14884_binop_int6435904_arg\(80 to 95), X"000" & X"1") & \$14884_binop_int6435904_arg\(96 to 151) & \$14884_binop_int6435904_arg\(152 to 153);
                  result6468 := \$14884_binop_int6435904_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$14941_modulo6685888_arg\ := work.Int.sub(\$14941_modulo6685888_arg\(0 to 30), \$14941_modulo6685888_arg\(31 to 61)) & \$14941_modulo6685888_arg\(31 to 61);
                  state_var7460 := \$14941_MODULO6685888\;
                end if;
              when \$14964_BINOP_INT6435905\ =>
                \$v7070\ := \$ram_lock\;
                if \$v7070\(0) = '1' then
                  state_var7460 := Q_WAIT7069;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$14964_binop_int6435905_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7068;
                end if;
              when \$14989_MODULO6685895\ =>
                \$v7062\ := work.Int.lt(\$14989_modulo6685895_arg\(0 to 30), \$14989_modulo6685895_arg\(31 to 61));
                if \$v7062\(0) = '1' then
                  \$14989_modulo6685895_result\ := \$14989_modulo6685895_arg\(0 to 30);
                  \$14986_r\ := \$14989_modulo6685895_result\;
                  \$14982_res\ := eclat_if(work.Int.lt(\$14964_binop_int6435905_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$14986_r\) & \$14986_r\);
                  \$14964_binop_int6435905_result\ := work.Int.add(\$14964_binop_int6435905_arg\(32 to 47), X"000" & X"1") & \$14982_res\ & eclat_true & 
                  work.Int.sub(\$14964_binop_int6435905_arg\(80 to 95), X"000" & X"1") & \$14964_binop_int6435905_arg\(96 to 151) & \$14964_binop_int6435905_arg\(152 to 153);
                  result6468 := \$14964_binop_int6435905_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$14997_modulo6685888_id\ := "000001011100";
                  \$14997_modulo6685888_arg\ := work.Int.sub(\$14989_modulo6685895_arg\(0 to 30), \$14989_modulo6685895_arg\(31 to 61)) & \$14989_modulo6685895_arg\(31 to 61);
                  state_var7460 := \$14997_MODULO6685888\;
                end if;
              when \$14997_MODULO6685888\ =>
                \$v7061\ := work.Int.lt(\$14997_modulo6685888_arg\(0 to 30), \$14997_modulo6685888_arg\(31 to 61));
                if \$v7061\(0) = '1' then
                  \$14997_modulo6685888_result\ := \$14997_modulo6685888_arg\(0 to 30);
                  \$14989_modulo6685895_result\ := \$14997_modulo6685888_result\;
                  \$14986_r\ := \$14989_modulo6685895_result\;
                  \$14982_res\ := eclat_if(work.Int.lt(\$14964_binop_int6435905_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$14986_r\) & \$14986_r\);
                  \$14964_binop_int6435905_result\ := work.Int.add(\$14964_binop_int6435905_arg\(32 to 47), X"000" & X"1") & \$14982_res\ & eclat_true & 
                  work.Int.sub(\$14964_binop_int6435905_arg\(80 to 95), X"000" & X"1") & \$14964_binop_int6435905_arg\(96 to 151) & \$14964_binop_int6435905_arg\(152 to 153);
                  result6468 := \$14964_binop_int6435905_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$14997_modulo6685888_arg\ := work.Int.sub(\$14997_modulo6685888_arg\(0 to 30), \$14997_modulo6685888_arg\(31 to 61)) & \$14997_modulo6685888_arg\(31 to 61);
                  state_var7460 := \$14997_MODULO6685888\;
                end if;
              when \$15013_MODULO6685896\ =>
                \$v7065\ := work.Int.lt(\$15013_modulo6685896_arg\(0 to 30), \$15013_modulo6685896_arg\(31 to 61));
                if \$v7065\(0) = '1' then
                  \$15013_modulo6685896_result\ := \$15013_modulo6685896_arg\(0 to 30);
                  \$15010_r\ := \$15013_modulo6685896_result\;
                  \$14982_res\ := eclat_if(work.Int.lt(\$14964_binop_int6435905_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$15010_r\) & \$15010_r\);
                  \$14964_binop_int6435905_result\ := work.Int.add(\$14964_binop_int6435905_arg\(32 to 47), X"000" & X"1") & \$14982_res\ & eclat_true & 
                  work.Int.sub(\$14964_binop_int6435905_arg\(80 to 95), X"000" & X"1") & \$14964_binop_int6435905_arg\(96 to 151) & \$14964_binop_int6435905_arg\(152 to 153);
                  result6468 := \$14964_binop_int6435905_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$15021_modulo6685888_id\ := "000001011110";
                  \$15021_modulo6685888_arg\ := work.Int.sub(\$15013_modulo6685896_arg\(0 to 30), \$15013_modulo6685896_arg\(31 to 61)) & \$15013_modulo6685896_arg\(31 to 61);
                  state_var7460 := \$15021_MODULO6685888\;
                end if;
              when \$15021_MODULO6685888\ =>
                \$v7064\ := work.Int.lt(\$15021_modulo6685888_arg\(0 to 30), \$15021_modulo6685888_arg\(31 to 61));
                if \$v7064\(0) = '1' then
                  \$15021_modulo6685888_result\ := \$15021_modulo6685888_arg\(0 to 30);
                  \$15013_modulo6685896_result\ := \$15021_modulo6685888_result\;
                  \$15010_r\ := \$15013_modulo6685896_result\;
                  \$14982_res\ := eclat_if(work.Int.lt(\$14964_binop_int6435905_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$15010_r\) & \$15010_r\);
                  \$14964_binop_int6435905_result\ := work.Int.add(\$14964_binop_int6435905_arg\(32 to 47), X"000" & X"1") & \$14982_res\ & eclat_true & 
                  work.Int.sub(\$14964_binop_int6435905_arg\(80 to 95), X"000" & X"1") & \$14964_binop_int6435905_arg\(96 to 151) & \$14964_binop_int6435905_arg\(152 to 153);
                  result6468 := \$14964_binop_int6435905_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$15021_modulo6685888_arg\ := work.Int.sub(\$15021_modulo6685888_arg\(0 to 30), \$15021_modulo6685888_arg\(31 to 61)) & \$15021_modulo6685888_arg\(31 to 61);
                  state_var7460 := \$15021_MODULO6685888\;
                end if;
              when \$15044_BINOP_INT6435906\ =>
                \$v7080\ := \$ram_lock\;
                if \$v7080\(0) = '1' then
                  state_var7460 := Q_WAIT7079;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$15044_binop_int6435906_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7078;
                end if;
              when \$15069_MODULO6685895\ =>
                \$v7072\ := work.Int.lt(\$15069_modulo6685895_arg\(0 to 30), \$15069_modulo6685895_arg\(31 to 61));
                if \$v7072\(0) = '1' then
                  \$15069_modulo6685895_result\ := \$15069_modulo6685895_arg\(0 to 30);
                  \$15066_r\ := \$15069_modulo6685895_result\;
                  \$15062_res\ := eclat_if(work.Int.lt(\$15044_binop_int6435906_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$15066_r\) & \$15066_r\);
                  \$15044_binop_int6435906_result\ := work.Int.add(\$15044_binop_int6435906_arg\(32 to 47), X"000" & X"1") & \$15062_res\ & eclat_true & 
                  work.Int.sub(\$15044_binop_int6435906_arg\(80 to 95), X"000" & X"1") & \$15044_binop_int6435906_arg\(96 to 151) & \$15044_binop_int6435906_arg\(152 to 153);
                  result6468 := \$15044_binop_int6435906_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$15077_modulo6685888_id\ := "000001100001";
                  \$15077_modulo6685888_arg\ := work.Int.sub(\$15069_modulo6685895_arg\(0 to 30), \$15069_modulo6685895_arg\(31 to 61)) & \$15069_modulo6685895_arg\(31 to 61);
                  state_var7460 := \$15077_MODULO6685888\;
                end if;
              when \$15077_MODULO6685888\ =>
                \$v7071\ := work.Int.lt(\$15077_modulo6685888_arg\(0 to 30), \$15077_modulo6685888_arg\(31 to 61));
                if \$v7071\(0) = '1' then
                  \$15077_modulo6685888_result\ := \$15077_modulo6685888_arg\(0 to 30);
                  \$15069_modulo6685895_result\ := \$15077_modulo6685888_result\;
                  \$15066_r\ := \$15069_modulo6685895_result\;
                  \$15062_res\ := eclat_if(work.Int.lt(\$15044_binop_int6435906_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$15066_r\) & \$15066_r\);
                  \$15044_binop_int6435906_result\ := work.Int.add(\$15044_binop_int6435906_arg\(32 to 47), X"000" & X"1") & \$15062_res\ & eclat_true & 
                  work.Int.sub(\$15044_binop_int6435906_arg\(80 to 95), X"000" & X"1") & \$15044_binop_int6435906_arg\(96 to 151) & \$15044_binop_int6435906_arg\(152 to 153);
                  result6468 := \$15044_binop_int6435906_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$15077_modulo6685888_arg\ := work.Int.sub(\$15077_modulo6685888_arg\(0 to 30), \$15077_modulo6685888_arg\(31 to 61)) & \$15077_modulo6685888_arg\(31 to 61);
                  state_var7460 := \$15077_MODULO6685888\;
                end if;
              when \$15093_MODULO6685896\ =>
                \$v7075\ := work.Int.lt(\$15093_modulo6685896_arg\(0 to 30), \$15093_modulo6685896_arg\(31 to 61));
                if \$v7075\(0) = '1' then
                  \$15093_modulo6685896_result\ := \$15093_modulo6685896_arg\(0 to 30);
                  \$15090_r\ := \$15093_modulo6685896_result\;
                  \$15062_res\ := eclat_if(work.Int.lt(\$15044_binop_int6435906_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$15090_r\) & \$15090_r\);
                  \$15044_binop_int6435906_result\ := work.Int.add(\$15044_binop_int6435906_arg\(32 to 47), X"000" & X"1") & \$15062_res\ & eclat_true & 
                  work.Int.sub(\$15044_binop_int6435906_arg\(80 to 95), X"000" & X"1") & \$15044_binop_int6435906_arg\(96 to 151) & \$15044_binop_int6435906_arg\(152 to 153);
                  result6468 := \$15044_binop_int6435906_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$15101_modulo6685888_id\ := "000001100011";
                  \$15101_modulo6685888_arg\ := work.Int.sub(\$15093_modulo6685896_arg\(0 to 30), \$15093_modulo6685896_arg\(31 to 61)) & \$15093_modulo6685896_arg\(31 to 61);
                  state_var7460 := \$15101_MODULO6685888\;
                end if;
              when \$15101_MODULO6685888\ =>
                \$v7074\ := work.Int.lt(\$15101_modulo6685888_arg\(0 to 30), \$15101_modulo6685888_arg\(31 to 61));
                if \$v7074\(0) = '1' then
                  \$15101_modulo6685888_result\ := \$15101_modulo6685888_arg\(0 to 30);
                  \$15093_modulo6685896_result\ := \$15101_modulo6685888_result\;
                  \$15090_r\ := \$15093_modulo6685896_result\;
                  \$15062_res\ := eclat_if(work.Int.lt(\$15044_binop_int6435906_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$15090_r\) & \$15090_r\);
                  \$15044_binop_int6435906_result\ := work.Int.add(\$15044_binop_int6435906_arg\(32 to 47), X"000" & X"1") & \$15062_res\ & eclat_true & 
                  work.Int.sub(\$15044_binop_int6435906_arg\(80 to 95), X"000" & X"1") & \$15044_binop_int6435906_arg\(96 to 151) & \$15044_binop_int6435906_arg\(152 to 153);
                  result6468 := \$15044_binop_int6435906_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$15101_modulo6685888_arg\ := work.Int.sub(\$15101_modulo6685888_arg\(0 to 30), \$15101_modulo6685888_arg\(31 to 61)) & \$15101_modulo6685888_arg\(31 to 61);
                  state_var7460 := \$15101_MODULO6685888\;
                end if;
              when \$15124_BINOP_INT6435907\ =>
                \$v7090\ := \$ram_lock\;
                if \$v7090\(0) = '1' then
                  state_var7460 := Q_WAIT7089;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$15124_binop_int6435907_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7088;
                end if;
              when \$15149_MODULO6685895\ =>
                \$v7082\ := work.Int.lt(\$15149_modulo6685895_arg\(0 to 30), \$15149_modulo6685895_arg\(31 to 61));
                if \$v7082\(0) = '1' then
                  \$15149_modulo6685895_result\ := \$15149_modulo6685895_arg\(0 to 30);
                  \$15146_r\ := \$15149_modulo6685895_result\;
                  \$15142_res\ := eclat_if(work.Int.lt(\$15124_binop_int6435907_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$15146_r\) & \$15146_r\);
                  \$15124_binop_int6435907_result\ := work.Int.add(\$15124_binop_int6435907_arg\(32 to 47), X"000" & X"1") & \$15142_res\ & eclat_true & 
                  work.Int.sub(\$15124_binop_int6435907_arg\(80 to 95), X"000" & X"1") & \$15124_binop_int6435907_arg\(96 to 151) & \$15124_binop_int6435907_arg\(152 to 153);
                  result6468 := \$15124_binop_int6435907_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$15157_modulo6685888_id\ := "000001100110";
                  \$15157_modulo6685888_arg\ := work.Int.sub(\$15149_modulo6685895_arg\(0 to 30), \$15149_modulo6685895_arg\(31 to 61)) & \$15149_modulo6685895_arg\(31 to 61);
                  state_var7460 := \$15157_MODULO6685888\;
                end if;
              when \$15157_MODULO6685888\ =>
                \$v7081\ := work.Int.lt(\$15157_modulo6685888_arg\(0 to 30), \$15157_modulo6685888_arg\(31 to 61));
                if \$v7081\(0) = '1' then
                  \$15157_modulo6685888_result\ := \$15157_modulo6685888_arg\(0 to 30);
                  \$15149_modulo6685895_result\ := \$15157_modulo6685888_result\;
                  \$15146_r\ := \$15149_modulo6685895_result\;
                  \$15142_res\ := eclat_if(work.Int.lt(\$15124_binop_int6435907_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$15146_r\) & \$15146_r\);
                  \$15124_binop_int6435907_result\ := work.Int.add(\$15124_binop_int6435907_arg\(32 to 47), X"000" & X"1") & \$15142_res\ & eclat_true & 
                  work.Int.sub(\$15124_binop_int6435907_arg\(80 to 95), X"000" & X"1") & \$15124_binop_int6435907_arg\(96 to 151) & \$15124_binop_int6435907_arg\(152 to 153);
                  result6468 := \$15124_binop_int6435907_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$15157_modulo6685888_arg\ := work.Int.sub(\$15157_modulo6685888_arg\(0 to 30), \$15157_modulo6685888_arg\(31 to 61)) & \$15157_modulo6685888_arg\(31 to 61);
                  state_var7460 := \$15157_MODULO6685888\;
                end if;
              when \$15173_MODULO6685896\ =>
                \$v7085\ := work.Int.lt(\$15173_modulo6685896_arg\(0 to 30), \$15173_modulo6685896_arg\(31 to 61));
                if \$v7085\(0) = '1' then
                  \$15173_modulo6685896_result\ := \$15173_modulo6685896_arg\(0 to 30);
                  \$15170_r\ := \$15173_modulo6685896_result\;
                  \$15142_res\ := eclat_if(work.Int.lt(\$15124_binop_int6435907_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$15170_r\) & \$15170_r\);
                  \$15124_binop_int6435907_result\ := work.Int.add(\$15124_binop_int6435907_arg\(32 to 47), X"000" & X"1") & \$15142_res\ & eclat_true & 
                  work.Int.sub(\$15124_binop_int6435907_arg\(80 to 95), X"000" & X"1") & \$15124_binop_int6435907_arg\(96 to 151) & \$15124_binop_int6435907_arg\(152 to 153);
                  result6468 := \$15124_binop_int6435907_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$15181_modulo6685888_id\ := "000001101000";
                  \$15181_modulo6685888_arg\ := work.Int.sub(\$15173_modulo6685896_arg\(0 to 30), \$15173_modulo6685896_arg\(31 to 61)) & \$15173_modulo6685896_arg\(31 to 61);
                  state_var7460 := \$15181_MODULO6685888\;
                end if;
              when \$15181_MODULO6685888\ =>
                \$v7084\ := work.Int.lt(\$15181_modulo6685888_arg\(0 to 30), \$15181_modulo6685888_arg\(31 to 61));
                if \$v7084\(0) = '1' then
                  \$15181_modulo6685888_result\ := \$15181_modulo6685888_arg\(0 to 30);
                  \$15173_modulo6685896_result\ := \$15181_modulo6685888_result\;
                  \$15170_r\ := \$15173_modulo6685896_result\;
                  \$15142_res\ := eclat_if(work.Int.lt(\$15124_binop_int6435907_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$15170_r\) & \$15170_r\);
                  \$15124_binop_int6435907_result\ := work.Int.add(\$15124_binop_int6435907_arg\(32 to 47), X"000" & X"1") & \$15142_res\ & eclat_true & 
                  work.Int.sub(\$15124_binop_int6435907_arg\(80 to 95), X"000" & X"1") & \$15124_binop_int6435907_arg\(96 to 151) & \$15124_binop_int6435907_arg\(152 to 153);
                  result6468 := \$15124_binop_int6435907_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$15181_modulo6685888_arg\ := work.Int.sub(\$15181_modulo6685888_arg\(0 to 30), \$15181_modulo6685888_arg\(31 to 61)) & \$15181_modulo6685888_arg\(31 to 61);
                  state_var7460 := \$15181_MODULO6685888\;
                end if;
              when \$15204_BINOP_INT6435908\ =>
                \$v7100\ := \$ram_lock\;
                if \$v7100\(0) = '1' then
                  state_var7460 := Q_WAIT7099;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$15204_binop_int6435908_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7098;
                end if;
              when \$15229_MODULO6685895\ =>
                \$v7092\ := work.Int.lt(\$15229_modulo6685895_arg\(0 to 30), \$15229_modulo6685895_arg\(31 to 61));
                if \$v7092\(0) = '1' then
                  \$15229_modulo6685895_result\ := \$15229_modulo6685895_arg\(0 to 30);
                  \$15226_r\ := \$15229_modulo6685895_result\;
                  \$15222_res\ := eclat_if(work.Int.lt(\$15204_binop_int6435908_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$15226_r\) & \$15226_r\);
                  \$15204_binop_int6435908_result\ := work.Int.add(\$15204_binop_int6435908_arg\(32 to 47), X"000" & X"1") & \$15222_res\ & eclat_true & 
                  work.Int.sub(\$15204_binop_int6435908_arg\(80 to 95), X"000" & X"1") & \$15204_binop_int6435908_arg\(96 to 151) & \$15204_binop_int6435908_arg\(152 to 153);
                  result6468 := \$15204_binop_int6435908_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$15237_modulo6685888_id\ := "000001101011";
                  \$15237_modulo6685888_arg\ := work.Int.sub(\$15229_modulo6685895_arg\(0 to 30), \$15229_modulo6685895_arg\(31 to 61)) & \$15229_modulo6685895_arg\(31 to 61);
                  state_var7460 := \$15237_MODULO6685888\;
                end if;
              when \$15237_MODULO6685888\ =>
                \$v7091\ := work.Int.lt(\$15237_modulo6685888_arg\(0 to 30), \$15237_modulo6685888_arg\(31 to 61));
                if \$v7091\(0) = '1' then
                  \$15237_modulo6685888_result\ := \$15237_modulo6685888_arg\(0 to 30);
                  \$15229_modulo6685895_result\ := \$15237_modulo6685888_result\;
                  \$15226_r\ := \$15229_modulo6685895_result\;
                  \$15222_res\ := eclat_if(work.Int.lt(\$15204_binop_int6435908_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$15226_r\) & \$15226_r\);
                  \$15204_binop_int6435908_result\ := work.Int.add(\$15204_binop_int6435908_arg\(32 to 47), X"000" & X"1") & \$15222_res\ & eclat_true & 
                  work.Int.sub(\$15204_binop_int6435908_arg\(80 to 95), X"000" & X"1") & \$15204_binop_int6435908_arg\(96 to 151) & \$15204_binop_int6435908_arg\(152 to 153);
                  result6468 := \$15204_binop_int6435908_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$15237_modulo6685888_arg\ := work.Int.sub(\$15237_modulo6685888_arg\(0 to 30), \$15237_modulo6685888_arg\(31 to 61)) & \$15237_modulo6685888_arg\(31 to 61);
                  state_var7460 := \$15237_MODULO6685888\;
                end if;
              when \$15253_MODULO6685896\ =>
                \$v7095\ := work.Int.lt(\$15253_modulo6685896_arg\(0 to 30), \$15253_modulo6685896_arg\(31 to 61));
                if \$v7095\(0) = '1' then
                  \$15253_modulo6685896_result\ := \$15253_modulo6685896_arg\(0 to 30);
                  \$15250_r\ := \$15253_modulo6685896_result\;
                  \$15222_res\ := eclat_if(work.Int.lt(\$15204_binop_int6435908_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$15250_r\) & \$15250_r\);
                  \$15204_binop_int6435908_result\ := work.Int.add(\$15204_binop_int6435908_arg\(32 to 47), X"000" & X"1") & \$15222_res\ & eclat_true & 
                  work.Int.sub(\$15204_binop_int6435908_arg\(80 to 95), X"000" & X"1") & \$15204_binop_int6435908_arg\(96 to 151) & \$15204_binop_int6435908_arg\(152 to 153);
                  result6468 := \$15204_binop_int6435908_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$15261_modulo6685888_id\ := "000001101101";
                  \$15261_modulo6685888_arg\ := work.Int.sub(\$15253_modulo6685896_arg\(0 to 30), \$15253_modulo6685896_arg\(31 to 61)) & \$15253_modulo6685896_arg\(31 to 61);
                  state_var7460 := \$15261_MODULO6685888\;
                end if;
              when \$15261_MODULO6685888\ =>
                \$v7094\ := work.Int.lt(\$15261_modulo6685888_arg\(0 to 30), \$15261_modulo6685888_arg\(31 to 61));
                if \$v7094\(0) = '1' then
                  \$15261_modulo6685888_result\ := \$15261_modulo6685888_arg\(0 to 30);
                  \$15253_modulo6685896_result\ := \$15261_modulo6685888_result\;
                  \$15250_r\ := \$15253_modulo6685896_result\;
                  \$15222_res\ := eclat_if(work.Int.lt(\$15204_binop_int6435908_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$15250_r\) & \$15250_r\);
                  \$15204_binop_int6435908_result\ := work.Int.add(\$15204_binop_int6435908_arg\(32 to 47), X"000" & X"1") & \$15222_res\ & eclat_true & 
                  work.Int.sub(\$15204_binop_int6435908_arg\(80 to 95), X"000" & X"1") & \$15204_binop_int6435908_arg\(96 to 151) & \$15204_binop_int6435908_arg\(152 to 153);
                  result6468 := \$15204_binop_int6435908_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$15261_modulo6685888_arg\ := work.Int.sub(\$15261_modulo6685888_arg\(0 to 30), \$15261_modulo6685888_arg\(31 to 61)) & \$15261_modulo6685888_arg\(31 to 61);
                  state_var7460 := \$15261_MODULO6685888\;
                end if;
              when \$15284_BINOP_INT6435909\ =>
                \$v7110\ := \$ram_lock\;
                if \$v7110\(0) = '1' then
                  state_var7460 := Q_WAIT7109;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$15284_binop_int6435909_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7108;
                end if;
              when \$15309_MODULO6685895\ =>
                \$v7102\ := work.Int.lt(\$15309_modulo6685895_arg\(0 to 30), \$15309_modulo6685895_arg\(31 to 61));
                if \$v7102\(0) = '1' then
                  \$15309_modulo6685895_result\ := \$15309_modulo6685895_arg\(0 to 30);
                  \$15306_r\ := \$15309_modulo6685895_result\;
                  \$15302_res\ := eclat_if(work.Int.lt(\$15284_binop_int6435909_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$15306_r\) & \$15306_r\);
                  \$15284_binop_int6435909_result\ := work.Int.add(\$15284_binop_int6435909_arg\(32 to 47), X"000" & X"1") & \$15302_res\ & eclat_true & 
                  work.Int.sub(\$15284_binop_int6435909_arg\(80 to 95), X"000" & X"1") & \$15284_binop_int6435909_arg\(96 to 151) & \$15284_binop_int6435909_arg\(152 to 153);
                  result6468 := \$15284_binop_int6435909_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$15317_modulo6685888_id\ := "000001110000";
                  \$15317_modulo6685888_arg\ := work.Int.sub(\$15309_modulo6685895_arg\(0 to 30), \$15309_modulo6685895_arg\(31 to 61)) & \$15309_modulo6685895_arg\(31 to 61);
                  state_var7460 := \$15317_MODULO6685888\;
                end if;
              when \$15317_MODULO6685888\ =>
                \$v7101\ := work.Int.lt(\$15317_modulo6685888_arg\(0 to 30), \$15317_modulo6685888_arg\(31 to 61));
                if \$v7101\(0) = '1' then
                  \$15317_modulo6685888_result\ := \$15317_modulo6685888_arg\(0 to 30);
                  \$15309_modulo6685895_result\ := \$15317_modulo6685888_result\;
                  \$15306_r\ := \$15309_modulo6685895_result\;
                  \$15302_res\ := eclat_if(work.Int.lt(\$15284_binop_int6435909_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$15306_r\) & \$15306_r\);
                  \$15284_binop_int6435909_result\ := work.Int.add(\$15284_binop_int6435909_arg\(32 to 47), X"000" & X"1") & \$15302_res\ & eclat_true & 
                  work.Int.sub(\$15284_binop_int6435909_arg\(80 to 95), X"000" & X"1") & \$15284_binop_int6435909_arg\(96 to 151) & \$15284_binop_int6435909_arg\(152 to 153);
                  result6468 := \$15284_binop_int6435909_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$15317_modulo6685888_arg\ := work.Int.sub(\$15317_modulo6685888_arg\(0 to 30), \$15317_modulo6685888_arg\(31 to 61)) & \$15317_modulo6685888_arg\(31 to 61);
                  state_var7460 := \$15317_MODULO6685888\;
                end if;
              when \$15333_MODULO6685896\ =>
                \$v7105\ := work.Int.lt(\$15333_modulo6685896_arg\(0 to 30), \$15333_modulo6685896_arg\(31 to 61));
                if \$v7105\(0) = '1' then
                  \$15333_modulo6685896_result\ := \$15333_modulo6685896_arg\(0 to 30);
                  \$15330_r\ := \$15333_modulo6685896_result\;
                  \$15302_res\ := eclat_if(work.Int.lt(\$15284_binop_int6435909_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$15330_r\) & \$15330_r\);
                  \$15284_binop_int6435909_result\ := work.Int.add(\$15284_binop_int6435909_arg\(32 to 47), X"000" & X"1") & \$15302_res\ & eclat_true & 
                  work.Int.sub(\$15284_binop_int6435909_arg\(80 to 95), X"000" & X"1") & \$15284_binop_int6435909_arg\(96 to 151) & \$15284_binop_int6435909_arg\(152 to 153);
                  result6468 := \$15284_binop_int6435909_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$15341_modulo6685888_id\ := "000001110010";
                  \$15341_modulo6685888_arg\ := work.Int.sub(\$15333_modulo6685896_arg\(0 to 30), \$15333_modulo6685896_arg\(31 to 61)) & \$15333_modulo6685896_arg\(31 to 61);
                  state_var7460 := \$15341_MODULO6685888\;
                end if;
              when \$15341_MODULO6685888\ =>
                \$v7104\ := work.Int.lt(\$15341_modulo6685888_arg\(0 to 30), \$15341_modulo6685888_arg\(31 to 61));
                if \$v7104\(0) = '1' then
                  \$15341_modulo6685888_result\ := \$15341_modulo6685888_arg\(0 to 30);
                  \$15333_modulo6685896_result\ := \$15341_modulo6685888_result\;
                  \$15330_r\ := \$15333_modulo6685896_result\;
                  \$15302_res\ := eclat_if(work.Int.lt(\$15284_binop_int6435909_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$15330_r\) & \$15330_r\);
                  \$15284_binop_int6435909_result\ := work.Int.add(\$15284_binop_int6435909_arg\(32 to 47), X"000" & X"1") & \$15302_res\ & eclat_true & 
                  work.Int.sub(\$15284_binop_int6435909_arg\(80 to 95), X"000" & X"1") & \$15284_binop_int6435909_arg\(96 to 151) & \$15284_binop_int6435909_arg\(152 to 153);
                  result6468 := \$15284_binop_int6435909_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$15341_modulo6685888_arg\ := work.Int.sub(\$15341_modulo6685888_arg\(0 to 30), \$15341_modulo6685888_arg\(31 to 61)) & \$15341_modulo6685888_arg\(31 to 61);
                  state_var7460 := \$15341_MODULO6685888\;
                end if;
              when \$15364_BINOP_INT6435910\ =>
                \$v7120\ := \$ram_lock\;
                if \$v7120\(0) = '1' then
                  state_var7460 := Q_WAIT7119;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$15364_binop_int6435910_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7118;
                end if;
              when \$15389_MODULO6685895\ =>
                \$v7112\ := work.Int.lt(\$15389_modulo6685895_arg\(0 to 30), \$15389_modulo6685895_arg\(31 to 61));
                if \$v7112\(0) = '1' then
                  \$15389_modulo6685895_result\ := \$15389_modulo6685895_arg\(0 to 30);
                  \$15386_r\ := \$15389_modulo6685895_result\;
                  \$15382_res\ := eclat_if(work.Int.lt(\$15364_binop_int6435910_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$15386_r\) & \$15386_r\);
                  \$15364_binop_int6435910_result\ := work.Int.add(\$15364_binop_int6435910_arg\(32 to 47), X"000" & X"1") & \$15382_res\ & eclat_true & 
                  work.Int.sub(\$15364_binop_int6435910_arg\(80 to 95), X"000" & X"1") & \$15364_binop_int6435910_arg\(96 to 151) & \$15364_binop_int6435910_arg\(152 to 153);
                  result6468 := \$15364_binop_int6435910_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$15397_modulo6685888_id\ := "000001110101";
                  \$15397_modulo6685888_arg\ := work.Int.sub(\$15389_modulo6685895_arg\(0 to 30), \$15389_modulo6685895_arg\(31 to 61)) & \$15389_modulo6685895_arg\(31 to 61);
                  state_var7460 := \$15397_MODULO6685888\;
                end if;
              when \$15397_MODULO6685888\ =>
                \$v7111\ := work.Int.lt(\$15397_modulo6685888_arg\(0 to 30), \$15397_modulo6685888_arg\(31 to 61));
                if \$v7111\(0) = '1' then
                  \$15397_modulo6685888_result\ := \$15397_modulo6685888_arg\(0 to 30);
                  \$15389_modulo6685895_result\ := \$15397_modulo6685888_result\;
                  \$15386_r\ := \$15389_modulo6685895_result\;
                  \$15382_res\ := eclat_if(work.Int.lt(\$15364_binop_int6435910_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$15386_r\) & \$15386_r\);
                  \$15364_binop_int6435910_result\ := work.Int.add(\$15364_binop_int6435910_arg\(32 to 47), X"000" & X"1") & \$15382_res\ & eclat_true & 
                  work.Int.sub(\$15364_binop_int6435910_arg\(80 to 95), X"000" & X"1") & \$15364_binop_int6435910_arg\(96 to 151) & \$15364_binop_int6435910_arg\(152 to 153);
                  result6468 := \$15364_binop_int6435910_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$15397_modulo6685888_arg\ := work.Int.sub(\$15397_modulo6685888_arg\(0 to 30), \$15397_modulo6685888_arg\(31 to 61)) & \$15397_modulo6685888_arg\(31 to 61);
                  state_var7460 := \$15397_MODULO6685888\;
                end if;
              when \$15413_MODULO6685896\ =>
                \$v7115\ := work.Int.lt(\$15413_modulo6685896_arg\(0 to 30), \$15413_modulo6685896_arg\(31 to 61));
                if \$v7115\(0) = '1' then
                  \$15413_modulo6685896_result\ := \$15413_modulo6685896_arg\(0 to 30);
                  \$15410_r\ := \$15413_modulo6685896_result\;
                  \$15382_res\ := eclat_if(work.Int.lt(\$15364_binop_int6435910_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$15410_r\) & \$15410_r\);
                  \$15364_binop_int6435910_result\ := work.Int.add(\$15364_binop_int6435910_arg\(32 to 47), X"000" & X"1") & \$15382_res\ & eclat_true & 
                  work.Int.sub(\$15364_binop_int6435910_arg\(80 to 95), X"000" & X"1") & \$15364_binop_int6435910_arg\(96 to 151) & \$15364_binop_int6435910_arg\(152 to 153);
                  result6468 := \$15364_binop_int6435910_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$15421_modulo6685888_id\ := "000001110111";
                  \$15421_modulo6685888_arg\ := work.Int.sub(\$15413_modulo6685896_arg\(0 to 30), \$15413_modulo6685896_arg\(31 to 61)) & \$15413_modulo6685896_arg\(31 to 61);
                  state_var7460 := \$15421_MODULO6685888\;
                end if;
              when \$15421_MODULO6685888\ =>
                \$v7114\ := work.Int.lt(\$15421_modulo6685888_arg\(0 to 30), \$15421_modulo6685888_arg\(31 to 61));
                if \$v7114\(0) = '1' then
                  \$15421_modulo6685888_result\ := \$15421_modulo6685888_arg\(0 to 30);
                  \$15413_modulo6685896_result\ := \$15421_modulo6685888_result\;
                  \$15410_r\ := \$15413_modulo6685896_result\;
                  \$15382_res\ := eclat_if(work.Int.lt(\$15364_binop_int6435910_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$15410_r\) & \$15410_r\);
                  \$15364_binop_int6435910_result\ := work.Int.add(\$15364_binop_int6435910_arg\(32 to 47), X"000" & X"1") & \$15382_res\ & eclat_true & 
                  work.Int.sub(\$15364_binop_int6435910_arg\(80 to 95), X"000" & X"1") & \$15364_binop_int6435910_arg\(96 to 151) & \$15364_binop_int6435910_arg\(152 to 153);
                  result6468 := \$15364_binop_int6435910_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$15421_modulo6685888_arg\ := work.Int.sub(\$15421_modulo6685888_arg\(0 to 30), \$15421_modulo6685888_arg\(31 to 61)) & \$15421_modulo6685888_arg\(31 to 61);
                  state_var7460 := \$15421_MODULO6685888\;
                end if;
              when \$15447_FOREVER6705911\ =>
                \$15447_forever6705911_arg\ := eclat_unit;
                state_var7460 := \$15447_FOREVER6705911\;
              when \$15451_BINOP_INT6435912\ =>
                \$v7130\ := \$ram_lock\;
                if \$v7130\(0) = '1' then
                  state_var7460 := Q_WAIT7129;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$15451_binop_int6435912_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7128;
                end if;
              when \$15476_MODULO6685895\ =>
                \$v7122\ := work.Int.lt(\$15476_modulo6685895_arg\(0 to 30), \$15476_modulo6685895_arg\(31 to 61));
                if \$v7122\(0) = '1' then
                  \$15476_modulo6685895_result\ := \$15476_modulo6685895_arg\(0 to 30);
                  \$15473_r\ := \$15476_modulo6685895_result\;
                  \$15469_res\ := eclat_if(work.Int.lt(\$15451_binop_int6435912_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$15473_r\) & \$15473_r\);
                  \$15451_binop_int6435912_result\ := work.Int.add(\$15451_binop_int6435912_arg\(32 to 47), X"000" & X"1") & \$15469_res\ & eclat_true & 
                  work.Int.sub(\$15451_binop_int6435912_arg\(80 to 95), X"000" & X"1") & \$15451_binop_int6435912_arg\(96 to 151) & \$15451_binop_int6435912_arg\(152 to 153);
                  result6468 := \$15451_binop_int6435912_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$15484_modulo6685888_id\ := "000001111011";
                  \$15484_modulo6685888_arg\ := work.Int.sub(\$15476_modulo6685895_arg\(0 to 30), \$15476_modulo6685895_arg\(31 to 61)) & \$15476_modulo6685895_arg\(31 to 61);
                  state_var7460 := \$15484_MODULO6685888\;
                end if;
              when \$15484_MODULO6685888\ =>
                \$v7121\ := work.Int.lt(\$15484_modulo6685888_arg\(0 to 30), \$15484_modulo6685888_arg\(31 to 61));
                if \$v7121\(0) = '1' then
                  \$15484_modulo6685888_result\ := \$15484_modulo6685888_arg\(0 to 30);
                  \$15476_modulo6685895_result\ := \$15484_modulo6685888_result\;
                  \$15473_r\ := \$15476_modulo6685895_result\;
                  \$15469_res\ := eclat_if(work.Int.lt(\$15451_binop_int6435912_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$15473_r\) & \$15473_r\);
                  \$15451_binop_int6435912_result\ := work.Int.add(\$15451_binop_int6435912_arg\(32 to 47), X"000" & X"1") & \$15469_res\ & eclat_true & 
                  work.Int.sub(\$15451_binop_int6435912_arg\(80 to 95), X"000" & X"1") & \$15451_binop_int6435912_arg\(96 to 151) & \$15451_binop_int6435912_arg\(152 to 153);
                  result6468 := \$15451_binop_int6435912_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$15484_modulo6685888_arg\ := work.Int.sub(\$15484_modulo6685888_arg\(0 to 30), \$15484_modulo6685888_arg\(31 to 61)) & \$15484_modulo6685888_arg\(31 to 61);
                  state_var7460 := \$15484_MODULO6685888\;
                end if;
              when \$15500_MODULO6685896\ =>
                \$v7125\ := work.Int.lt(\$15500_modulo6685896_arg\(0 to 30), \$15500_modulo6685896_arg\(31 to 61));
                if \$v7125\(0) = '1' then
                  \$15500_modulo6685896_result\ := \$15500_modulo6685896_arg\(0 to 30);
                  \$15497_r\ := \$15500_modulo6685896_result\;
                  \$15469_res\ := eclat_if(work.Int.lt(\$15451_binop_int6435912_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$15497_r\) & \$15497_r\);
                  \$15451_binop_int6435912_result\ := work.Int.add(\$15451_binop_int6435912_arg\(32 to 47), X"000" & X"1") & \$15469_res\ & eclat_true & 
                  work.Int.sub(\$15451_binop_int6435912_arg\(80 to 95), X"000" & X"1") & \$15451_binop_int6435912_arg\(96 to 151) & \$15451_binop_int6435912_arg\(152 to 153);
                  result6468 := \$15451_binop_int6435912_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$15508_modulo6685888_id\ := "000001111101";
                  \$15508_modulo6685888_arg\ := work.Int.sub(\$15500_modulo6685896_arg\(0 to 30), \$15500_modulo6685896_arg\(31 to 61)) & \$15500_modulo6685896_arg\(31 to 61);
                  state_var7460 := \$15508_MODULO6685888\;
                end if;
              when \$15508_MODULO6685888\ =>
                \$v7124\ := work.Int.lt(\$15508_modulo6685888_arg\(0 to 30), \$15508_modulo6685888_arg\(31 to 61));
                if \$v7124\(0) = '1' then
                  \$15508_modulo6685888_result\ := \$15508_modulo6685888_arg\(0 to 30);
                  \$15500_modulo6685896_result\ := \$15508_modulo6685888_result\;
                  \$15497_r\ := \$15500_modulo6685896_result\;
                  \$15469_res\ := eclat_if(work.Int.lt(\$15451_binop_int6435912_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$15497_r\) & \$15497_r\);
                  \$15451_binop_int6435912_result\ := work.Int.add(\$15451_binop_int6435912_arg\(32 to 47), X"000" & X"1") & \$15469_res\ & eclat_true & 
                  work.Int.sub(\$15451_binop_int6435912_arg\(80 to 95), X"000" & X"1") & \$15451_binop_int6435912_arg\(96 to 151) & \$15451_binop_int6435912_arg\(152 to 153);
                  result6468 := \$15451_binop_int6435912_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$15508_modulo6685888_arg\ := work.Int.sub(\$15508_modulo6685888_arg\(0 to 30), \$15508_modulo6685888_arg\(31 to 61)) & \$15508_modulo6685888_arg\(31 to 61);
                  state_var7460 := \$15508_MODULO6685888\;
                end if;
              when \$15531_BINOP_INT6435913\ =>
                \$v7140\ := \$ram_lock\;
                if \$v7140\(0) = '1' then
                  state_var7460 := Q_WAIT7139;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$15531_binop_int6435913_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7138;
                end if;
              when \$15556_MODULO6685895\ =>
                \$v7132\ := work.Int.lt(\$15556_modulo6685895_arg\(0 to 30), \$15556_modulo6685895_arg\(31 to 61));
                if \$v7132\(0) = '1' then
                  \$15556_modulo6685895_result\ := \$15556_modulo6685895_arg\(0 to 30);
                  \$15553_r\ := \$15556_modulo6685895_result\;
                  \$15549_res\ := eclat_if(work.Int.lt(\$15531_binop_int6435913_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$15553_r\) & \$15553_r\);
                  \$15531_binop_int6435913_result\ := work.Int.add(\$15531_binop_int6435913_arg\(32 to 47), X"000" & X"1") & \$15549_res\ & eclat_true & 
                  work.Int.sub(\$15531_binop_int6435913_arg\(80 to 95), X"000" & X"1") & \$15531_binop_int6435913_arg\(96 to 151) & \$15531_binop_int6435913_arg\(152 to 153);
                  result6468 := \$15531_binop_int6435913_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$15564_modulo6685888_id\ := "000010000000";
                  \$15564_modulo6685888_arg\ := work.Int.sub(\$15556_modulo6685895_arg\(0 to 30), \$15556_modulo6685895_arg\(31 to 61)) & \$15556_modulo6685895_arg\(31 to 61);
                  state_var7460 := \$15564_MODULO6685888\;
                end if;
              when \$15564_MODULO6685888\ =>
                \$v7131\ := work.Int.lt(\$15564_modulo6685888_arg\(0 to 30), \$15564_modulo6685888_arg\(31 to 61));
                if \$v7131\(0) = '1' then
                  \$15564_modulo6685888_result\ := \$15564_modulo6685888_arg\(0 to 30);
                  \$15556_modulo6685895_result\ := \$15564_modulo6685888_result\;
                  \$15553_r\ := \$15556_modulo6685895_result\;
                  \$15549_res\ := eclat_if(work.Int.lt(\$15531_binop_int6435913_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$15553_r\) & \$15553_r\);
                  \$15531_binop_int6435913_result\ := work.Int.add(\$15531_binop_int6435913_arg\(32 to 47), X"000" & X"1") & \$15549_res\ & eclat_true & 
                  work.Int.sub(\$15531_binop_int6435913_arg\(80 to 95), X"000" & X"1") & \$15531_binop_int6435913_arg\(96 to 151) & \$15531_binop_int6435913_arg\(152 to 153);
                  result6468 := \$15531_binop_int6435913_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$15564_modulo6685888_arg\ := work.Int.sub(\$15564_modulo6685888_arg\(0 to 30), \$15564_modulo6685888_arg\(31 to 61)) & \$15564_modulo6685888_arg\(31 to 61);
                  state_var7460 := \$15564_MODULO6685888\;
                end if;
              when \$15580_MODULO6685896\ =>
                \$v7135\ := work.Int.lt(\$15580_modulo6685896_arg\(0 to 30), \$15580_modulo6685896_arg\(31 to 61));
                if \$v7135\(0) = '1' then
                  \$15580_modulo6685896_result\ := \$15580_modulo6685896_arg\(0 to 30);
                  \$15577_r\ := \$15580_modulo6685896_result\;
                  \$15549_res\ := eclat_if(work.Int.lt(\$15531_binop_int6435913_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$15577_r\) & \$15577_r\);
                  \$15531_binop_int6435913_result\ := work.Int.add(\$15531_binop_int6435913_arg\(32 to 47), X"000" & X"1") & \$15549_res\ & eclat_true & 
                  work.Int.sub(\$15531_binop_int6435913_arg\(80 to 95), X"000" & X"1") & \$15531_binop_int6435913_arg\(96 to 151) & \$15531_binop_int6435913_arg\(152 to 153);
                  result6468 := \$15531_binop_int6435913_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$15588_modulo6685888_id\ := "000010000010";
                  \$15588_modulo6685888_arg\ := work.Int.sub(\$15580_modulo6685896_arg\(0 to 30), \$15580_modulo6685896_arg\(31 to 61)) & \$15580_modulo6685896_arg\(31 to 61);
                  state_var7460 := \$15588_MODULO6685888\;
                end if;
              when \$15588_MODULO6685888\ =>
                \$v7134\ := work.Int.lt(\$15588_modulo6685888_arg\(0 to 30), \$15588_modulo6685888_arg\(31 to 61));
                if \$v7134\(0) = '1' then
                  \$15588_modulo6685888_result\ := \$15588_modulo6685888_arg\(0 to 30);
                  \$15580_modulo6685896_result\ := \$15588_modulo6685888_result\;
                  \$15577_r\ := \$15580_modulo6685896_result\;
                  \$15549_res\ := eclat_if(work.Int.lt(\$15531_binop_int6435913_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  work.Int.sub("000"& X"000000" & X"0", \$15577_r\) & \$15577_r\);
                  \$15531_binop_int6435913_result\ := work.Int.add(\$15531_binop_int6435913_arg\(32 to 47), X"000" & X"1") & \$15549_res\ & eclat_true & 
                  work.Int.sub(\$15531_binop_int6435913_arg\(80 to 95), X"000" & X"1") & \$15531_binop_int6435913_arg\(96 to 151) & \$15531_binop_int6435913_arg\(152 to 153);
                  result6468 := \$15531_binop_int6435913_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$15588_modulo6685888_arg\ := work.Int.sub(\$15588_modulo6685888_arg\(0 to 30), \$15588_modulo6685888_arg\(31 to 61)) & \$15588_modulo6685888_arg\(31 to 61);
                  state_var7460 := \$15588_MODULO6685888\;
                end if;
              when \$15614_FOREVER6705914\ =>
                \$15614_forever6705914_arg\ := eclat_unit;
                state_var7460 := \$15614_FOREVER6705914\;
              when \$15621_FOREVER6705915\ =>
                \$15621_forever6705915_arg\ := eclat_unit;
                state_var7460 := \$15621_FOREVER6705915\;
              when \$15625_BINOP_COMPARE6455916\ =>
                \$v7144\ := \$ram_lock\;
                if \$v7144\(0) = '1' then
                  state_var7460 := Q_WAIT7143;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$15625_binop_compare6455916_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7142;
                end if;
              when \$15648_COMPARE6445897\ =>
                \$v7141\ := \$15648_compare6445897_arg\(0 to 31);
                case \$v7141\ is
                when X"0000000" & X"0" =>
                  \$15648_compare6445897_result\ := work.Int.eq(\$15648_compare6445897_arg\(32 to 62), \$15648_compare6445897_arg\(63 to 93));
                when X"0000000" & X"1" =>
                  \$15648_compare6445897_result\ := work.Bool.lnot(work.Int.eq(
                                                                   \$15648_compare6445897_arg\(32 to 62), \$15648_compare6445897_arg\(63 to 93)));
                when X"0000000" & X"2" =>
                  \$15648_compare6445897_result\ := work.Int.lt(\$15648_compare6445897_arg\(32 to 62), \$15648_compare6445897_arg\(63 to 93));
                when X"0000000" & X"3" =>
                  \$15648_compare6445897_result\ := eclat_if(work.Int.lt(
                                                             \$15648_compare6445897_arg\(32 to 62), \$15648_compare6445897_arg\(63 to 93)) & eclat_true & 
                                                    work.Int.eq(\$15648_compare6445897_arg\(32 to 62), \$15648_compare6445897_arg\(63 to 93)));
                when X"0000000" & X"4" =>
                  \$15648_compare6445897_result\ := work.Bool.lnot(eclat_if(
                                                                   work.Int.lt(
                                                                   \$15648_compare6445897_arg\(32 to 62), \$15648_compare6445897_arg\(63 to 93)) & eclat_true & 
                                                                   work.Int.eq(
                                                                   \$15648_compare6445897_arg\(32 to 62), \$15648_compare6445897_arg\(63 to 93))));
                when X"0000000" & X"5" =>
                  \$15648_compare6445897_result\ := work.Bool.lnot(work.Int.lt(
                                                                   \$15648_compare6445897_arg\(32 to 62), \$15648_compare6445897_arg\(63 to 93)));
                when others =>
                  \$15648_compare6445897_result\ := eclat_false;
                end case;
                \$15643_res\ := \$15648_compare6445897_result\;
                \$15625_binop_compare6455916_result\ := work.Int.add(
                                                        \$15625_binop_compare6455916_arg\(32 to 47), X"000" & X"1") & 
                eclat_if(\$15643_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & 
                work.Int.sub(\$15625_binop_compare6455916_arg\(80 to 95), X"000" & X"1") & \$15625_binop_compare6455916_arg\(96 to 151) & \$15625_binop_compare6455916_arg\(152 to 153);
                result6468 := \$15625_binop_compare6455916_result\;
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when \$15661_BINOP_COMPARE6455917\ =>
                \$v7148\ := \$ram_lock\;
                if \$v7148\(0) = '1' then
                  state_var7460 := Q_WAIT7147;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$15661_binop_compare6455917_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7146;
                end if;
              when \$15684_COMPARE6445897\ =>
                \$v7145\ := \$15684_compare6445897_arg\(0 to 31);
                case \$v7145\ is
                when X"0000000" & X"0" =>
                  \$15684_compare6445897_result\ := work.Int.eq(\$15684_compare6445897_arg\(32 to 62), \$15684_compare6445897_arg\(63 to 93));
                when X"0000000" & X"1" =>
                  \$15684_compare6445897_result\ := work.Bool.lnot(work.Int.eq(
                                                                   \$15684_compare6445897_arg\(32 to 62), \$15684_compare6445897_arg\(63 to 93)));
                when X"0000000" & X"2" =>
                  \$15684_compare6445897_result\ := work.Int.lt(\$15684_compare6445897_arg\(32 to 62), \$15684_compare6445897_arg\(63 to 93));
                when X"0000000" & X"3" =>
                  \$15684_compare6445897_result\ := eclat_if(work.Int.lt(
                                                             \$15684_compare6445897_arg\(32 to 62), \$15684_compare6445897_arg\(63 to 93)) & eclat_true & 
                                                    work.Int.eq(\$15684_compare6445897_arg\(32 to 62), \$15684_compare6445897_arg\(63 to 93)));
                when X"0000000" & X"4" =>
                  \$15684_compare6445897_result\ := work.Bool.lnot(eclat_if(
                                                                   work.Int.lt(
                                                                   \$15684_compare6445897_arg\(32 to 62), \$15684_compare6445897_arg\(63 to 93)) & eclat_true & 
                                                                   work.Int.eq(
                                                                   \$15684_compare6445897_arg\(32 to 62), \$15684_compare6445897_arg\(63 to 93))));
                when X"0000000" & X"5" =>
                  \$15684_compare6445897_result\ := work.Bool.lnot(work.Int.lt(
                                                                   \$15684_compare6445897_arg\(32 to 62), \$15684_compare6445897_arg\(63 to 93)));
                when others =>
                  \$15684_compare6445897_result\ := eclat_false;
                end case;
                \$15679_res\ := \$15684_compare6445897_result\;
                \$15661_binop_compare6455917_result\ := work.Int.add(
                                                        \$15661_binop_compare6455917_arg\(32 to 47), X"000" & X"1") & 
                eclat_if(\$15679_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & 
                work.Int.sub(\$15661_binop_compare6455917_arg\(80 to 95), X"000" & X"1") & \$15661_binop_compare6455917_arg\(96 to 151) & \$15661_binop_compare6455917_arg\(152 to 153);
                result6468 := \$15661_binop_compare6455917_result\;
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when \$15697_BINOP_COMPARE6455918\ =>
                \$v7152\ := \$ram_lock\;
                if \$v7152\(0) = '1' then
                  state_var7460 := Q_WAIT7151;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$15697_binop_compare6455918_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7150;
                end if;
              when \$15720_COMPARE6445897\ =>
                \$v7149\ := \$15720_compare6445897_arg\(0 to 31);
                case \$v7149\ is
                when X"0000000" & X"0" =>
                  \$15720_compare6445897_result\ := work.Int.eq(\$15720_compare6445897_arg\(32 to 62), \$15720_compare6445897_arg\(63 to 93));
                when X"0000000" & X"1" =>
                  \$15720_compare6445897_result\ := work.Bool.lnot(work.Int.eq(
                                                                   \$15720_compare6445897_arg\(32 to 62), \$15720_compare6445897_arg\(63 to 93)));
                when X"0000000" & X"2" =>
                  \$15720_compare6445897_result\ := work.Int.lt(\$15720_compare6445897_arg\(32 to 62), \$15720_compare6445897_arg\(63 to 93));
                when X"0000000" & X"3" =>
                  \$15720_compare6445897_result\ := eclat_if(work.Int.lt(
                                                             \$15720_compare6445897_arg\(32 to 62), \$15720_compare6445897_arg\(63 to 93)) & eclat_true & 
                                                    work.Int.eq(\$15720_compare6445897_arg\(32 to 62), \$15720_compare6445897_arg\(63 to 93)));
                when X"0000000" & X"4" =>
                  \$15720_compare6445897_result\ := work.Bool.lnot(eclat_if(
                                                                   work.Int.lt(
                                                                   \$15720_compare6445897_arg\(32 to 62), \$15720_compare6445897_arg\(63 to 93)) & eclat_true & 
                                                                   work.Int.eq(
                                                                   \$15720_compare6445897_arg\(32 to 62), \$15720_compare6445897_arg\(63 to 93))));
                when X"0000000" & X"5" =>
                  \$15720_compare6445897_result\ := work.Bool.lnot(work.Int.lt(
                                                                   \$15720_compare6445897_arg\(32 to 62), \$15720_compare6445897_arg\(63 to 93)));
                when others =>
                  \$15720_compare6445897_result\ := eclat_false;
                end case;
                \$15715_res\ := \$15720_compare6445897_result\;
                \$15697_binop_compare6455918_result\ := work.Int.add(
                                                        \$15697_binop_compare6455918_arg\(32 to 47), X"000" & X"1") & 
                eclat_if(\$15715_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & 
                work.Int.sub(\$15697_binop_compare6455918_arg\(80 to 95), X"000" & X"1") & \$15697_binop_compare6455918_arg\(96 to 151) & \$15697_binop_compare6455918_arg\(152 to 153);
                result6468 := \$15697_binop_compare6455918_result\;
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when \$15733_BINOP_COMPARE6455919\ =>
                \$v7156\ := \$ram_lock\;
                if \$v7156\(0) = '1' then
                  state_var7460 := Q_WAIT7155;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$15733_binop_compare6455919_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7154;
                end if;
              when \$15756_COMPARE6445897\ =>
                \$v7153\ := \$15756_compare6445897_arg\(0 to 31);
                case \$v7153\ is
                when X"0000000" & X"0" =>
                  \$15756_compare6445897_result\ := work.Int.eq(\$15756_compare6445897_arg\(32 to 62), \$15756_compare6445897_arg\(63 to 93));
                when X"0000000" & X"1" =>
                  \$15756_compare6445897_result\ := work.Bool.lnot(work.Int.eq(
                                                                   \$15756_compare6445897_arg\(32 to 62), \$15756_compare6445897_arg\(63 to 93)));
                when X"0000000" & X"2" =>
                  \$15756_compare6445897_result\ := work.Int.lt(\$15756_compare6445897_arg\(32 to 62), \$15756_compare6445897_arg\(63 to 93));
                when X"0000000" & X"3" =>
                  \$15756_compare6445897_result\ := eclat_if(work.Int.lt(
                                                             \$15756_compare6445897_arg\(32 to 62), \$15756_compare6445897_arg\(63 to 93)) & eclat_true & 
                                                    work.Int.eq(\$15756_compare6445897_arg\(32 to 62), \$15756_compare6445897_arg\(63 to 93)));
                when X"0000000" & X"4" =>
                  \$15756_compare6445897_result\ := work.Bool.lnot(eclat_if(
                                                                   work.Int.lt(
                                                                   \$15756_compare6445897_arg\(32 to 62), \$15756_compare6445897_arg\(63 to 93)) & eclat_true & 
                                                                   work.Int.eq(
                                                                   \$15756_compare6445897_arg\(32 to 62), \$15756_compare6445897_arg\(63 to 93))));
                when X"0000000" & X"5" =>
                  \$15756_compare6445897_result\ := work.Bool.lnot(work.Int.lt(
                                                                   \$15756_compare6445897_arg\(32 to 62), \$15756_compare6445897_arg\(63 to 93)));
                when others =>
                  \$15756_compare6445897_result\ := eclat_false;
                end case;
                \$15751_res\ := \$15756_compare6445897_result\;
                \$15733_binop_compare6455919_result\ := work.Int.add(
                                                        \$15733_binop_compare6455919_arg\(32 to 47), X"000" & X"1") & 
                eclat_if(\$15751_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & 
                work.Int.sub(\$15733_binop_compare6455919_arg\(80 to 95), X"000" & X"1") & \$15733_binop_compare6455919_arg\(96 to 151) & \$15733_binop_compare6455919_arg\(152 to 153);
                result6468 := \$15733_binop_compare6455919_result\;
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when \$15769_BINOP_COMPARE6455920\ =>
                \$v7160\ := \$ram_lock\;
                if \$v7160\(0) = '1' then
                  state_var7460 := Q_WAIT7159;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$15769_binop_compare6455920_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7158;
                end if;
              when \$15792_COMPARE6445897\ =>
                \$v7157\ := \$15792_compare6445897_arg\(0 to 31);
                case \$v7157\ is
                when X"0000000" & X"0" =>
                  \$15792_compare6445897_result\ := work.Int.eq(\$15792_compare6445897_arg\(32 to 62), \$15792_compare6445897_arg\(63 to 93));
                when X"0000000" & X"1" =>
                  \$15792_compare6445897_result\ := work.Bool.lnot(work.Int.eq(
                                                                   \$15792_compare6445897_arg\(32 to 62), \$15792_compare6445897_arg\(63 to 93)));
                when X"0000000" & X"2" =>
                  \$15792_compare6445897_result\ := work.Int.lt(\$15792_compare6445897_arg\(32 to 62), \$15792_compare6445897_arg\(63 to 93));
                when X"0000000" & X"3" =>
                  \$15792_compare6445897_result\ := eclat_if(work.Int.lt(
                                                             \$15792_compare6445897_arg\(32 to 62), \$15792_compare6445897_arg\(63 to 93)) & eclat_true & 
                                                    work.Int.eq(\$15792_compare6445897_arg\(32 to 62), \$15792_compare6445897_arg\(63 to 93)));
                when X"0000000" & X"4" =>
                  \$15792_compare6445897_result\ := work.Bool.lnot(eclat_if(
                                                                   work.Int.lt(
                                                                   \$15792_compare6445897_arg\(32 to 62), \$15792_compare6445897_arg\(63 to 93)) & eclat_true & 
                                                                   work.Int.eq(
                                                                   \$15792_compare6445897_arg\(32 to 62), \$15792_compare6445897_arg\(63 to 93))));
                when X"0000000" & X"5" =>
                  \$15792_compare6445897_result\ := work.Bool.lnot(work.Int.lt(
                                                                   \$15792_compare6445897_arg\(32 to 62), \$15792_compare6445897_arg\(63 to 93)));
                when others =>
                  \$15792_compare6445897_result\ := eclat_false;
                end case;
                \$15787_res\ := \$15792_compare6445897_result\;
                \$15769_binop_compare6455920_result\ := work.Int.add(
                                                        \$15769_binop_compare6455920_arg\(32 to 47), X"000" & X"1") & 
                eclat_if(\$15787_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & 
                work.Int.sub(\$15769_binop_compare6455920_arg\(80 to 95), X"000" & X"1") & \$15769_binop_compare6455920_arg\(96 to 151) & \$15769_binop_compare6455920_arg\(152 to 153);
                result6468 := \$15769_binop_compare6455920_result\;
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when \$15805_BINOP_COMPARE6455921\ =>
                \$v7164\ := \$ram_lock\;
                if \$v7164\(0) = '1' then
                  state_var7460 := Q_WAIT7163;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$15805_binop_compare6455921_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7162;
                end if;
              when \$15828_COMPARE6445897\ =>
                \$v7161\ := \$15828_compare6445897_arg\(0 to 31);
                case \$v7161\ is
                when X"0000000" & X"0" =>
                  \$15828_compare6445897_result\ := work.Int.eq(\$15828_compare6445897_arg\(32 to 62), \$15828_compare6445897_arg\(63 to 93));
                when X"0000000" & X"1" =>
                  \$15828_compare6445897_result\ := work.Bool.lnot(work.Int.eq(
                                                                   \$15828_compare6445897_arg\(32 to 62), \$15828_compare6445897_arg\(63 to 93)));
                when X"0000000" & X"2" =>
                  \$15828_compare6445897_result\ := work.Int.lt(\$15828_compare6445897_arg\(32 to 62), \$15828_compare6445897_arg\(63 to 93));
                when X"0000000" & X"3" =>
                  \$15828_compare6445897_result\ := eclat_if(work.Int.lt(
                                                             \$15828_compare6445897_arg\(32 to 62), \$15828_compare6445897_arg\(63 to 93)) & eclat_true & 
                                                    work.Int.eq(\$15828_compare6445897_arg\(32 to 62), \$15828_compare6445897_arg\(63 to 93)));
                when X"0000000" & X"4" =>
                  \$15828_compare6445897_result\ := work.Bool.lnot(eclat_if(
                                                                   work.Int.lt(
                                                                   \$15828_compare6445897_arg\(32 to 62), \$15828_compare6445897_arg\(63 to 93)) & eclat_true & 
                                                                   work.Int.eq(
                                                                   \$15828_compare6445897_arg\(32 to 62), \$15828_compare6445897_arg\(63 to 93))));
                when X"0000000" & X"5" =>
                  \$15828_compare6445897_result\ := work.Bool.lnot(work.Int.lt(
                                                                   \$15828_compare6445897_arg\(32 to 62), \$15828_compare6445897_arg\(63 to 93)));
                when others =>
                  \$15828_compare6445897_result\ := eclat_false;
                end case;
                \$15823_res\ := \$15828_compare6445897_result\;
                \$15805_binop_compare6455921_result\ := work.Int.add(
                                                        \$15805_binop_compare6455921_arg\(32 to 47), X"000" & X"1") & 
                eclat_if(\$15823_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & 
                work.Int.sub(\$15805_binop_compare6455921_arg\(80 to 95), X"000" & X"1") & \$15805_binop_compare6455921_arg\(96 to 151) & \$15805_binop_compare6455921_arg\(152 to 153);
                result6468 := \$15805_binop_compare6455921_result\;
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when \$16063_W6515922\ =>
                \$v7226\ := work.Int.gt(\$16063_w6515922_arg\(0 to 7), \$16063_w6515922_arg\(24 to 31));
                if \$v7226\(0) = '1' then
                  \$16063_w6515922_result\ := \$16063_w6515922_arg\(8 to 23);
                  \$16036_sp\ := \$16063_w6515922_result\;
                  \$v7219\ := \$ram_lock\;
                  if \$v7219\(0) = '1' then
                    state_var7460 := Q_WAIT7218;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$16036_sp\, X"000" & X"1")));
                    state_var7460 := PAUSE_GET7217;
                  end if;
                else
                  \$v7225\ := \$ram_lock\;
                  if \$v7225\(0) = '1' then
                    state_var7460 := Q_WAIT7224;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$16063_w6515922_arg\(8 to 23), X"000" & X"1")));
                    state_var7460 := PAUSE_GET7223;
                  end if;
                end if;
              when \$16158_FOREVER6705923\ =>
                \$16158_forever6705923_arg\ := eclat_unit;
                state_var7460 := \$16158_FOREVER6705923\;
              when \$16195_FOREVER6705924\ =>
                \$16195_forever6705924_arg\ := eclat_unit;
                state_var7460 := \$16195_FOREVER6705924\;
              when \$16510_FOREVER6705925\ =>
                \$16510_forever6705925_arg\ := eclat_unit;
                state_var7460 := \$16510_FOREVER6705925\;
              when \$16551_COMPBRANCH6505926\ =>
                \$16574_compare6445898_id\ := "000010100010";
                \$16574_compare6445898_arg\ := \$16551_compbranch6505926_arg\(0 to 31) & \$16551_compbranch6505926_arg\(32 to 62) & \$16551_compbranch6505926_arg\(110 to 140);
                state_var7460 := \$16574_COMPARE6445898\;
              when \$16574_COMPARE6445898\ =>
                \$v7354\ := \$16574_compare6445898_arg\(0 to 31);
                case \$v7354\ is
                when X"0000000" & X"0" =>
                  \$16574_compare6445898_result\ := work.Int.eq(\$16574_compare6445898_arg\(32 to 62), \$16574_compare6445898_arg\(63 to 93));
                when X"0000000" & X"1" =>
                  \$16574_compare6445898_result\ := work.Bool.lnot(work.Int.eq(
                                                                   \$16574_compare6445898_arg\(32 to 62), \$16574_compare6445898_arg\(63 to 93)));
                when X"0000000" & X"2" =>
                  \$16574_compare6445898_result\ := work.Int.lt(\$16574_compare6445898_arg\(32 to 62), \$16574_compare6445898_arg\(63 to 93));
                when X"0000000" & X"3" =>
                  \$16574_compare6445898_result\ := eclat_if(work.Int.lt(
                                                             \$16574_compare6445898_arg\(32 to 62), \$16574_compare6445898_arg\(63 to 93)) & eclat_true & 
                                                    work.Int.eq(\$16574_compare6445898_arg\(32 to 62), \$16574_compare6445898_arg\(63 to 93)));
                when X"0000000" & X"4" =>
                  \$16574_compare6445898_result\ := work.Bool.lnot(eclat_if(
                                                                   work.Int.lt(
                                                                   \$16574_compare6445898_arg\(32 to 62), \$16574_compare6445898_arg\(63 to 93)) & eclat_true & 
                                                                   work.Int.eq(
                                                                   \$16574_compare6445898_arg\(32 to 62), \$16574_compare6445898_arg\(63 to 93))));
                when X"0000000" & X"5" =>
                  \$16574_compare6445898_result\ := work.Bool.lnot(work.Int.lt(
                                                                   \$16574_compare6445898_arg\(32 to 62), \$16574_compare6445898_arg\(63 to 93)));
                when others =>
                  \$16574_compare6445898_result\ := eclat_false;
                end case;
                \$16568_b\ := \$16574_compare6445898_result\;
                \$16551_compbranch6505926_result\ := eclat_if(\$16568_b\ & 
                                                     work.Int.add(work.Int.add(
                                                                  \$16551_compbranch6505926_arg\(94 to 109), X"000" & X"2"), eclat_resize(\$16551_compbranch6505926_arg\(63 to 93),16)) & \$16551_compbranch6505926_arg\(110 to 141) & \$16551_compbranch6505926_arg\(142 to 157) & \$16551_compbranch6505926_arg\(158 to 213) & \$16551_compbranch6505926_arg\(214 to 215) & 
                                                     work.Int.add(\$16551_compbranch6505926_arg\(94 to 109), X"000" & X"3") & \$16551_compbranch6505926_arg\(110 to 141) & \$16551_compbranch6505926_arg\(142 to 157) & \$16551_compbranch6505926_arg\(158 to 213) & \$16551_compbranch6505926_arg\(214 to 215));
                result6468 := \$16551_compbranch6505926_result\;
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when \$16589_COMPBRANCH6505927\ =>
                \$16612_compare6445898_id\ := "000010100100";
                \$16612_compare6445898_arg\ := \$16589_compbranch6505927_arg\(0 to 31) & \$16589_compbranch6505927_arg\(32 to 62) & \$16589_compbranch6505927_arg\(110 to 140);
                state_var7460 := \$16612_COMPARE6445898\;
              when \$16612_COMPARE6445898\ =>
                \$v7355\ := \$16612_compare6445898_arg\(0 to 31);
                case \$v7355\ is
                when X"0000000" & X"0" =>
                  \$16612_compare6445898_result\ := work.Int.eq(\$16612_compare6445898_arg\(32 to 62), \$16612_compare6445898_arg\(63 to 93));
                when X"0000000" & X"1" =>
                  \$16612_compare6445898_result\ := work.Bool.lnot(work.Int.eq(
                                                                   \$16612_compare6445898_arg\(32 to 62), \$16612_compare6445898_arg\(63 to 93)));
                when X"0000000" & X"2" =>
                  \$16612_compare6445898_result\ := work.Int.lt(\$16612_compare6445898_arg\(32 to 62), \$16612_compare6445898_arg\(63 to 93));
                when X"0000000" & X"3" =>
                  \$16612_compare6445898_result\ := eclat_if(work.Int.lt(
                                                             \$16612_compare6445898_arg\(32 to 62), \$16612_compare6445898_arg\(63 to 93)) & eclat_true & 
                                                    work.Int.eq(\$16612_compare6445898_arg\(32 to 62), \$16612_compare6445898_arg\(63 to 93)));
                when X"0000000" & X"4" =>
                  \$16612_compare6445898_result\ := work.Bool.lnot(eclat_if(
                                                                   work.Int.lt(
                                                                   \$16612_compare6445898_arg\(32 to 62), \$16612_compare6445898_arg\(63 to 93)) & eclat_true & 
                                                                   work.Int.eq(
                                                                   \$16612_compare6445898_arg\(32 to 62), \$16612_compare6445898_arg\(63 to 93))));
                when X"0000000" & X"5" =>
                  \$16612_compare6445898_result\ := work.Bool.lnot(work.Int.lt(
                                                                   \$16612_compare6445898_arg\(32 to 62), \$16612_compare6445898_arg\(63 to 93)));
                when others =>
                  \$16612_compare6445898_result\ := eclat_false;
                end case;
                \$16606_b\ := \$16612_compare6445898_result\;
                \$16589_compbranch6505927_result\ := eclat_if(\$16606_b\ & 
                                                     work.Int.add(work.Int.add(
                                                                  \$16589_compbranch6505927_arg\(94 to 109), X"000" & X"2"), eclat_resize(\$16589_compbranch6505927_arg\(63 to 93),16)) & \$16589_compbranch6505927_arg\(110 to 141) & \$16589_compbranch6505927_arg\(142 to 157) & \$16589_compbranch6505927_arg\(158 to 213) & \$16589_compbranch6505927_arg\(214 to 215) & 
                                                     work.Int.add(\$16589_compbranch6505927_arg\(94 to 109), X"000" & X"3") & \$16589_compbranch6505927_arg\(110 to 141) & \$16589_compbranch6505927_arg\(142 to 157) & \$16589_compbranch6505927_arg\(158 to 213) & \$16589_compbranch6505927_arg\(214 to 215));
                result6468 := \$16589_compbranch6505927_result\;
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when \$16662_FILL6535928\ =>
                \$v7365\ := work.Int.gt(\$16662_fill6535928_arg\(0 to 15), \$16662_fill6535928_arg\(32 to 47));
                if \$v7365\(0) = '1' then
                  \$16662_fill6535928_result\ := \$16662_fill6535928_arg\(16 to 31);
                  \$16659_sp\ := \$16662_fill6535928_result\;
                  result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"3") & \$16651\(64 to 95) & \$16659_sp\ & \$16651\(32 to 63) & \$13911\(96 to 103) & \$13911\(104 to 119) & \$13911\(120 to 121);
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$v7364\ := \$ram_lock\;
                  if \$v7364\(0) = '1' then
                    state_var7460 := Q_WAIT7363;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$16662_fill6535928_arg\(16 to 31), X"000" & X"1")));
                    state_var7460 := PAUSE_GET7362;
                  end if;
                end if;
              when \$16752_FILL6545929\ =>
                \$v7394\ := work.Int.ge(\$16752_fill6545929_arg\(0 to 15), \$16752_fill6545929_arg\(32 to 47));
                if \$v7394\(0) = '1' then
                  \$16752_fill6545929_result\ := \$16752_fill6545929_arg\(16 to 31);
                  \$16749_sp\ := \$16752_fill6545929_result\;
                  result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"3") & \$16741\(64 to 95) & \$16749_sp\ & \$16741\(32 to 63) & \$13911\(96 to 103) & \$13911\(104 to 119) & \$13911\(120 to 121);
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$v7393\ := \$ram_lock\;
                  if \$v7393\(0) = '1' then
                    state_var7460 := Q_WAIT7392;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$16752_fill6545929_arg\(16 to 31), X"000" & X"1")));
                    state_var7460 := PAUSE_GET7391;
                  end if;
                end if;
              when \$16788_COMPBRANCH6505930\ =>
                \$16811_compare6445898_id\ := "000010101011";
                \$16811_compare6445898_arg\ := \$16788_compbranch6505930_arg\(0 to 31) & \$16788_compbranch6505930_arg\(32 to 62) & \$16788_compbranch6505930_arg\(110 to 140);
                state_var7460 := \$16811_COMPARE6445898\;
              when \$16811_COMPARE6445898\ =>
                \$v7398\ := \$16811_compare6445898_arg\(0 to 31);
                case \$v7398\ is
                when X"0000000" & X"0" =>
                  \$16811_compare6445898_result\ := work.Int.eq(\$16811_compare6445898_arg\(32 to 62), \$16811_compare6445898_arg\(63 to 93));
                when X"0000000" & X"1" =>
                  \$16811_compare6445898_result\ := work.Bool.lnot(work.Int.eq(
                                                                   \$16811_compare6445898_arg\(32 to 62), \$16811_compare6445898_arg\(63 to 93)));
                when X"0000000" & X"2" =>
                  \$16811_compare6445898_result\ := work.Int.lt(\$16811_compare6445898_arg\(32 to 62), \$16811_compare6445898_arg\(63 to 93));
                when X"0000000" & X"3" =>
                  \$16811_compare6445898_result\ := eclat_if(work.Int.lt(
                                                             \$16811_compare6445898_arg\(32 to 62), \$16811_compare6445898_arg\(63 to 93)) & eclat_true & 
                                                    work.Int.eq(\$16811_compare6445898_arg\(32 to 62), \$16811_compare6445898_arg\(63 to 93)));
                when X"0000000" & X"4" =>
                  \$16811_compare6445898_result\ := work.Bool.lnot(eclat_if(
                                                                   work.Int.lt(
                                                                   \$16811_compare6445898_arg\(32 to 62), \$16811_compare6445898_arg\(63 to 93)) & eclat_true & 
                                                                   work.Int.eq(
                                                                   \$16811_compare6445898_arg\(32 to 62), \$16811_compare6445898_arg\(63 to 93))));
                when X"0000000" & X"5" =>
                  \$16811_compare6445898_result\ := work.Bool.lnot(work.Int.lt(
                                                                   \$16811_compare6445898_arg\(32 to 62), \$16811_compare6445898_arg\(63 to 93)));
                when others =>
                  \$16811_compare6445898_result\ := eclat_false;
                end case;
                \$16805_b\ := \$16811_compare6445898_result\;
                \$16788_compbranch6505930_result\ := eclat_if(\$16805_b\ & 
                                                     work.Int.add(work.Int.add(
                                                                  \$16788_compbranch6505930_arg\(94 to 109), X"000" & X"2"), eclat_resize(\$16788_compbranch6505930_arg\(63 to 93),16)) & \$16788_compbranch6505930_arg\(110 to 141) & \$16788_compbranch6505930_arg\(142 to 157) & \$16788_compbranch6505930_arg\(158 to 213) & \$16788_compbranch6505930_arg\(214 to 215) & 
                                                     work.Int.add(\$16788_compbranch6505930_arg\(94 to 109), X"000" & X"3") & \$16788_compbranch6505930_arg\(110 to 141) & \$16788_compbranch6505930_arg\(142 to 157) & \$16788_compbranch6505930_arg\(158 to 213) & \$16788_compbranch6505930_arg\(214 to 215));
                result6468 := \$16788_compbranch6505930_result\;
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when \$16823_COMPBRANCH6505931\ =>
                \$16846_compare6445898_id\ := "000010101101";
                \$16846_compare6445898_arg\ := \$16823_compbranch6505931_arg\(0 to 31) & \$16823_compbranch6505931_arg\(32 to 62) & \$16823_compbranch6505931_arg\(110 to 140);
                state_var7460 := \$16846_COMPARE6445898\;
              when \$16846_COMPARE6445898\ =>
                \$v7399\ := \$16846_compare6445898_arg\(0 to 31);
                case \$v7399\ is
                when X"0000000" & X"0" =>
                  \$16846_compare6445898_result\ := work.Int.eq(\$16846_compare6445898_arg\(32 to 62), \$16846_compare6445898_arg\(63 to 93));
                when X"0000000" & X"1" =>
                  \$16846_compare6445898_result\ := work.Bool.lnot(work.Int.eq(
                                                                   \$16846_compare6445898_arg\(32 to 62), \$16846_compare6445898_arg\(63 to 93)));
                when X"0000000" & X"2" =>
                  \$16846_compare6445898_result\ := work.Int.lt(\$16846_compare6445898_arg\(32 to 62), \$16846_compare6445898_arg\(63 to 93));
                when X"0000000" & X"3" =>
                  \$16846_compare6445898_result\ := eclat_if(work.Int.lt(
                                                             \$16846_compare6445898_arg\(32 to 62), \$16846_compare6445898_arg\(63 to 93)) & eclat_true & 
                                                    work.Int.eq(\$16846_compare6445898_arg\(32 to 62), \$16846_compare6445898_arg\(63 to 93)));
                when X"0000000" & X"4" =>
                  \$16846_compare6445898_result\ := work.Bool.lnot(eclat_if(
                                                                   work.Int.lt(
                                                                   \$16846_compare6445898_arg\(32 to 62), \$16846_compare6445898_arg\(63 to 93)) & eclat_true & 
                                                                   work.Int.eq(
                                                                   \$16846_compare6445898_arg\(32 to 62), \$16846_compare6445898_arg\(63 to 93))));
                when X"0000000" & X"5" =>
                  \$16846_compare6445898_result\ := work.Bool.lnot(work.Int.lt(
                                                                   \$16846_compare6445898_arg\(32 to 62), \$16846_compare6445898_arg\(63 to 93)));
                when others =>
                  \$16846_compare6445898_result\ := eclat_false;
                end case;
                \$16840_b\ := \$16846_compare6445898_result\;
                \$16823_compbranch6505931_result\ := eclat_if(\$16840_b\ & 
                                                     work.Int.add(work.Int.add(
                                                                  \$16823_compbranch6505931_arg\(94 to 109), X"000" & X"2"), eclat_resize(\$16823_compbranch6505931_arg\(63 to 93),16)) & \$16823_compbranch6505931_arg\(110 to 141) & \$16823_compbranch6505931_arg\(142 to 157) & \$16823_compbranch6505931_arg\(158 to 213) & \$16823_compbranch6505931_arg\(214 to 215) & 
                                                     work.Int.add(\$16823_compbranch6505931_arg\(94 to 109), X"000" & X"3") & \$16823_compbranch6505931_arg\(110 to 141) & \$16823_compbranch6505931_arg\(142 to 157) & \$16823_compbranch6505931_arg\(158 to 213) & \$16823_compbranch6505931_arg\(214 to 215));
                result6468 := \$16823_compbranch6505931_result\;
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when \$16858_COMPBRANCH6505932\ =>
                \$16881_compare6445898_id\ := "000010101111";
                \$16881_compare6445898_arg\ := \$16858_compbranch6505932_arg\(0 to 31) & \$16858_compbranch6505932_arg\(32 to 62) & \$16858_compbranch6505932_arg\(110 to 140);
                state_var7460 := \$16881_COMPARE6445898\;
              when \$16881_COMPARE6445898\ =>
                \$v7400\ := \$16881_compare6445898_arg\(0 to 31);
                case \$v7400\ is
                when X"0000000" & X"0" =>
                  \$16881_compare6445898_result\ := work.Int.eq(\$16881_compare6445898_arg\(32 to 62), \$16881_compare6445898_arg\(63 to 93));
                when X"0000000" & X"1" =>
                  \$16881_compare6445898_result\ := work.Bool.lnot(work.Int.eq(
                                                                   \$16881_compare6445898_arg\(32 to 62), \$16881_compare6445898_arg\(63 to 93)));
                when X"0000000" & X"2" =>
                  \$16881_compare6445898_result\ := work.Int.lt(\$16881_compare6445898_arg\(32 to 62), \$16881_compare6445898_arg\(63 to 93));
                when X"0000000" & X"3" =>
                  \$16881_compare6445898_result\ := eclat_if(work.Int.lt(
                                                             \$16881_compare6445898_arg\(32 to 62), \$16881_compare6445898_arg\(63 to 93)) & eclat_true & 
                                                    work.Int.eq(\$16881_compare6445898_arg\(32 to 62), \$16881_compare6445898_arg\(63 to 93)));
                when X"0000000" & X"4" =>
                  \$16881_compare6445898_result\ := work.Bool.lnot(eclat_if(
                                                                   work.Int.lt(
                                                                   \$16881_compare6445898_arg\(32 to 62), \$16881_compare6445898_arg\(63 to 93)) & eclat_true & 
                                                                   work.Int.eq(
                                                                   \$16881_compare6445898_arg\(32 to 62), \$16881_compare6445898_arg\(63 to 93))));
                when X"0000000" & X"5" =>
                  \$16881_compare6445898_result\ := work.Bool.lnot(work.Int.lt(
                                                                   \$16881_compare6445898_arg\(32 to 62), \$16881_compare6445898_arg\(63 to 93)));
                when others =>
                  \$16881_compare6445898_result\ := eclat_false;
                end case;
                \$16875_b\ := \$16881_compare6445898_result\;
                \$16858_compbranch6505932_result\ := eclat_if(\$16875_b\ & 
                                                     work.Int.add(work.Int.add(
                                                                  \$16858_compbranch6505932_arg\(94 to 109), X"000" & X"2"), eclat_resize(\$16858_compbranch6505932_arg\(63 to 93),16)) & \$16858_compbranch6505932_arg\(110 to 141) & \$16858_compbranch6505932_arg\(142 to 157) & \$16858_compbranch6505932_arg\(158 to 213) & \$16858_compbranch6505932_arg\(214 to 215) & 
                                                     work.Int.add(\$16858_compbranch6505932_arg\(94 to 109), X"000" & X"3") & \$16858_compbranch6505932_arg\(110 to 141) & \$16858_compbranch6505932_arg\(142 to 157) & \$16858_compbranch6505932_arg\(158 to 213) & \$16858_compbranch6505932_arg\(214 to 215));
                result6468 := \$16858_compbranch6505932_result\;
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when \$16893_COMPBRANCH6505933\ =>
                \$16916_compare6445898_id\ := "000010110001";
                \$16916_compare6445898_arg\ := \$16893_compbranch6505933_arg\(0 to 31) & \$16893_compbranch6505933_arg\(32 to 62) & \$16893_compbranch6505933_arg\(110 to 140);
                state_var7460 := \$16916_COMPARE6445898\;
              when \$16916_COMPARE6445898\ =>
                \$v7401\ := \$16916_compare6445898_arg\(0 to 31);
                case \$v7401\ is
                when X"0000000" & X"0" =>
                  \$16916_compare6445898_result\ := work.Int.eq(\$16916_compare6445898_arg\(32 to 62), \$16916_compare6445898_arg\(63 to 93));
                when X"0000000" & X"1" =>
                  \$16916_compare6445898_result\ := work.Bool.lnot(work.Int.eq(
                                                                   \$16916_compare6445898_arg\(32 to 62), \$16916_compare6445898_arg\(63 to 93)));
                when X"0000000" & X"2" =>
                  \$16916_compare6445898_result\ := work.Int.lt(\$16916_compare6445898_arg\(32 to 62), \$16916_compare6445898_arg\(63 to 93));
                when X"0000000" & X"3" =>
                  \$16916_compare6445898_result\ := eclat_if(work.Int.lt(
                                                             \$16916_compare6445898_arg\(32 to 62), \$16916_compare6445898_arg\(63 to 93)) & eclat_true & 
                                                    work.Int.eq(\$16916_compare6445898_arg\(32 to 62), \$16916_compare6445898_arg\(63 to 93)));
                when X"0000000" & X"4" =>
                  \$16916_compare6445898_result\ := work.Bool.lnot(eclat_if(
                                                                   work.Int.lt(
                                                                   \$16916_compare6445898_arg\(32 to 62), \$16916_compare6445898_arg\(63 to 93)) & eclat_true & 
                                                                   work.Int.eq(
                                                                   \$16916_compare6445898_arg\(32 to 62), \$16916_compare6445898_arg\(63 to 93))));
                when X"0000000" & X"5" =>
                  \$16916_compare6445898_result\ := work.Bool.lnot(work.Int.lt(
                                                                   \$16916_compare6445898_arg\(32 to 62), \$16916_compare6445898_arg\(63 to 93)));
                when others =>
                  \$16916_compare6445898_result\ := eclat_false;
                end case;
                \$16910_b\ := \$16916_compare6445898_result\;
                \$16893_compbranch6505933_result\ := eclat_if(\$16910_b\ & 
                                                     work.Int.add(work.Int.add(
                                                                  \$16893_compbranch6505933_arg\(94 to 109), X"000" & X"2"), eclat_resize(\$16893_compbranch6505933_arg\(63 to 93),16)) & \$16893_compbranch6505933_arg\(110 to 141) & \$16893_compbranch6505933_arg\(142 to 157) & \$16893_compbranch6505933_arg\(158 to 213) & \$16893_compbranch6505933_arg\(214 to 215) & 
                                                     work.Int.add(\$16893_compbranch6505933_arg\(94 to 109), X"000" & X"3") & \$16893_compbranch6505933_arg\(110 to 141) & \$16893_compbranch6505933_arg\(142 to 157) & \$16893_compbranch6505933_arg\(158 to 213) & \$16893_compbranch6505933_arg\(214 to 215));
                result6468 := \$16893_compbranch6505933_result\;
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when \$16928_COMPBRANCH6505934\ =>
                \$16951_compare6445898_id\ := "000010110011";
                \$16951_compare6445898_arg\ := \$16928_compbranch6505934_arg\(0 to 31) & \$16928_compbranch6505934_arg\(32 to 62) & \$16928_compbranch6505934_arg\(110 to 140);
                state_var7460 := \$16951_COMPARE6445898\;
              when \$16951_COMPARE6445898\ =>
                \$v7402\ := \$16951_compare6445898_arg\(0 to 31);
                case \$v7402\ is
                when X"0000000" & X"0" =>
                  \$16951_compare6445898_result\ := work.Int.eq(\$16951_compare6445898_arg\(32 to 62), \$16951_compare6445898_arg\(63 to 93));
                when X"0000000" & X"1" =>
                  \$16951_compare6445898_result\ := work.Bool.lnot(work.Int.eq(
                                                                   \$16951_compare6445898_arg\(32 to 62), \$16951_compare6445898_arg\(63 to 93)));
                when X"0000000" & X"2" =>
                  \$16951_compare6445898_result\ := work.Int.lt(\$16951_compare6445898_arg\(32 to 62), \$16951_compare6445898_arg\(63 to 93));
                when X"0000000" & X"3" =>
                  \$16951_compare6445898_result\ := eclat_if(work.Int.lt(
                                                             \$16951_compare6445898_arg\(32 to 62), \$16951_compare6445898_arg\(63 to 93)) & eclat_true & 
                                                    work.Int.eq(\$16951_compare6445898_arg\(32 to 62), \$16951_compare6445898_arg\(63 to 93)));
                when X"0000000" & X"4" =>
                  \$16951_compare6445898_result\ := work.Bool.lnot(eclat_if(
                                                                   work.Int.lt(
                                                                   \$16951_compare6445898_arg\(32 to 62), \$16951_compare6445898_arg\(63 to 93)) & eclat_true & 
                                                                   work.Int.eq(
                                                                   \$16951_compare6445898_arg\(32 to 62), \$16951_compare6445898_arg\(63 to 93))));
                when X"0000000" & X"5" =>
                  \$16951_compare6445898_result\ := work.Bool.lnot(work.Int.lt(
                                                                   \$16951_compare6445898_arg\(32 to 62), \$16951_compare6445898_arg\(63 to 93)));
                when others =>
                  \$16951_compare6445898_result\ := eclat_false;
                end case;
                \$16945_b\ := \$16951_compare6445898_result\;
                \$16928_compbranch6505934_result\ := eclat_if(\$16945_b\ & 
                                                     work.Int.add(work.Int.add(
                                                                  \$16928_compbranch6505934_arg\(94 to 109), X"000" & X"2"), eclat_resize(\$16928_compbranch6505934_arg\(63 to 93),16)) & \$16928_compbranch6505934_arg\(110 to 141) & \$16928_compbranch6505934_arg\(142 to 157) & \$16928_compbranch6505934_arg\(158 to 213) & \$16928_compbranch6505934_arg\(214 to 215) & 
                                                     work.Int.add(\$16928_compbranch6505934_arg\(94 to 109), X"000" & X"3") & \$16928_compbranch6505934_arg\(110 to 141) & \$16928_compbranch6505934_arg\(142 to 157) & \$16928_compbranch6505934_arg\(158 to 213) & \$16928_compbranch6505934_arg\(214 to 215));
                result6468 := \$16928_compbranch6505934_result\;
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when \$16963_COMPBRANCH6505935\ =>
                \$16986_compare6445898_id\ := "000010110101";
                \$16986_compare6445898_arg\ := \$16963_compbranch6505935_arg\(0 to 31) & \$16963_compbranch6505935_arg\(32 to 62) & \$16963_compbranch6505935_arg\(110 to 140);
                state_var7460 := \$16986_COMPARE6445898\;
              when \$16986_COMPARE6445898\ =>
                \$v7403\ := \$16986_compare6445898_arg\(0 to 31);
                case \$v7403\ is
                when X"0000000" & X"0" =>
                  \$16986_compare6445898_result\ := work.Int.eq(\$16986_compare6445898_arg\(32 to 62), \$16986_compare6445898_arg\(63 to 93));
                when X"0000000" & X"1" =>
                  \$16986_compare6445898_result\ := work.Bool.lnot(work.Int.eq(
                                                                   \$16986_compare6445898_arg\(32 to 62), \$16986_compare6445898_arg\(63 to 93)));
                when X"0000000" & X"2" =>
                  \$16986_compare6445898_result\ := work.Int.lt(\$16986_compare6445898_arg\(32 to 62), \$16986_compare6445898_arg\(63 to 93));
                when X"0000000" & X"3" =>
                  \$16986_compare6445898_result\ := eclat_if(work.Int.lt(
                                                             \$16986_compare6445898_arg\(32 to 62), \$16986_compare6445898_arg\(63 to 93)) & eclat_true & 
                                                    work.Int.eq(\$16986_compare6445898_arg\(32 to 62), \$16986_compare6445898_arg\(63 to 93)));
                when X"0000000" & X"4" =>
                  \$16986_compare6445898_result\ := work.Bool.lnot(eclat_if(
                                                                   work.Int.lt(
                                                                   \$16986_compare6445898_arg\(32 to 62), \$16986_compare6445898_arg\(63 to 93)) & eclat_true & 
                                                                   work.Int.eq(
                                                                   \$16986_compare6445898_arg\(32 to 62), \$16986_compare6445898_arg\(63 to 93))));
                when X"0000000" & X"5" =>
                  \$16986_compare6445898_result\ := work.Bool.lnot(work.Int.lt(
                                                                   \$16986_compare6445898_arg\(32 to 62), \$16986_compare6445898_arg\(63 to 93)));
                when others =>
                  \$16986_compare6445898_result\ := eclat_false;
                end case;
                \$16980_b\ := \$16986_compare6445898_result\;
                \$16963_compbranch6505935_result\ := eclat_if(\$16980_b\ & 
                                                     work.Int.add(work.Int.add(
                                                                  \$16963_compbranch6505935_arg\(94 to 109), X"000" & X"2"), eclat_resize(\$16963_compbranch6505935_arg\(63 to 93),16)) & \$16963_compbranch6505935_arg\(110 to 141) & \$16963_compbranch6505935_arg\(142 to 157) & \$16963_compbranch6505935_arg\(158 to 213) & \$16963_compbranch6505935_arg\(214 to 215) & 
                                                     work.Int.add(\$16963_compbranch6505935_arg\(94 to 109), X"000" & X"3") & \$16963_compbranch6505935_arg\(110 to 141) & \$16963_compbranch6505935_arg\(142 to 157) & \$16963_compbranch6505935_arg\(158 to 213) & \$16963_compbranch6505935_arg\(214 to 215));
                result6468 := \$16963_compbranch6505935_result\;
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when \$17018_W36575938\ =>
                \$v7407\ := work.Int.ge(\$17018_w36575938_arg\(0 to 15), \$17018_w36575938_arg\(32 to 47));
                if \$v7407\(0) = '1' then
                  \$17018_w36575938_result\ := \$17018_w36575938_arg\(16 to 31);
                  \$17012_sp\ := \$17018_w36575938_result\;
                  result6468 := work.Int.add(work.Int.add(\$13911\(0 to 15), X"000" & X"3"), eclat_resize(\$15851_argument1\,16)) & \$17001\(64 to 95) & \$17012_sp\ & \$17001\(32 to 63) & \$13911\(96 to 103) & \$13911\(104 to 119) & \$13911\(120 to 121);
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                else
                  \$v7406\ := \$ram_lock\;
                  if \$v7406\(0) = '1' then
                    state_var7460 := Q_WAIT7405;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17018_w36575938_arg\(16 to 31)));
                    \$ram_write\ <= eclat_resize(work.Int.add(eclat_resize(\$17018_w36575938_arg\(48 to 78),16), 
                                                              work.Int.mul(
                                                              X"000" & X"2", \$17018_w36575938_arg\(0 to 15))),31) & eclat_true; \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET7404;
                  end if;
                end if;
              when \$17048_W16565937\ =>
                \$v7420\ := work.Int.ge(\$17048_w16565937_arg\(0 to 15), \$17048_w16565937_arg\(32 to 47));
                if \$v7420\(0) = '1' then
                  \$17048_w16565937_result\ := eclat_unit;
                  \$17010\ := \$17048_w16565937_result\;
                  \$v7410\ := \$ram_lock\;
                  if \$v7410\(0) = '1' then
                    state_var7460 := Q_WAIT7409;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17009_sp\));
                    \$ram_write\ <= \$17001\(64 to 95); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET7408;
                  end if;
                else
                  \$v7419\ := \$ram_lock\;
                  if \$v7419\(0) = '1' then
                    state_var7460 := Q_WAIT7418;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            work.Int.add(
                                                            eclat_resize(\$17048_w16565937_arg\(48 to 78),16), 
                                                            work.Int.sub(
                                                            work.Int.mul(
                                                            X"000" & X"2", \$17048_w16565937_arg\(0 to 15)), X"000" & X"1")), X"000" & X"1")));
                    \$ram_write\ <= work.Int.lor(work.Int.lsl(eclat_resize("11111001",31), X"000000" & X"18"), 
                                                 work.Int.lsl(eclat_resize(
                                                              work.Int.mul(
                                                              X"000" & X"2", \$17048_w16565937_arg\(0 to 15)),31), X"0000000" & X"2")) & eclat_true; \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET7417;
                  end if;
                end if;
              when \$17105_W06555936\ =>
                \$v7427\ := work.Int.ge(\$17105_w06555936_arg\(0 to 15), \$17105_w06555936_arg\(48 to 63));
                if \$v7427\(0) = '1' then
                  \$17105_w06555936_result\ := \$17105_w06555936_arg\(16 to 31);
                  \$17009_sp\ := \$17105_w06555936_result\;
                  \$17048_w16565937_id\ := "000010111000";
                  \$17048_w16565937_arg\ := X"000" & X"1" & \$13911\(0 to 15) & eclat_resize(\$15851_argument1\,16) & \$17001\(64 to 95);
                  state_var7460 := \$17048_W16565937\;
                else
                  \$v7426\ := \$ram_lock\;
                  if \$v7426\(0) = '1' then
                    state_var7460 := Q_WAIT7425;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$17105_w06555936_arg\(16 to 31), X"000" & X"1")));
                    state_var7460 := PAUSE_GET7424;
                  end if;
                end if;
              when PAUSE_GET6474 =>
                \$18545\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6473\ := \$ram_lock\;
                if \$v6473\(0) = '1' then
                  state_var7460 := Q_WAIT6472;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$13920_loop666_arg\(16 to 31), \$13920_loop666_arg\(0 to 15))));
                  \$ram_write\ <= \$18545\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6471;
                end if;
              when PAUSE_GET6490 =>
                \$18464_hd\ := \$ram_value\;
                release(\$ram_lock\);
                \$18468\ := work.Print.print_string(clk,of_string("bloc "));
                \$18469\ := work.Int.print(clk,eclat_resize(\$18443\(0 to 30),16));
                \$18470\ := work.Print.print_string(clk,of_string(" of size "));
                \$18471\ := work.Int.print(clk,work.Int.add(eclat_resize(
                                                            work.Int.lsr(
                                                            \$18464_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$18472\ := work.Print.print_string(clk,of_string(" from "));
                \$18473\ := work.Int.print(clk,eclat_resize(\$18443\(0 to 30),16));
                \$18474\ := work.Print.print_string(clk,of_string(" to "));
                \$18475\ := work.Int.print(clk,\$13921_loop665_arg\(16 to 31));
                \$18476\ := work.Print.print_newline(clk,eclat_unit);
                \$v6489\ := \$ram_lock\;
                if \$v6489\(0) = '1' then
                  state_var7460 := Q_WAIT6488;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13921_loop665_arg\(16 to 31)));
                  \$ram_write\ <= \$18464_hd\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6487;
                end if;
              when PAUSE_GET6494 =>
                \$18459_w\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6493\ := eclat_if(work.Bool.lnot(""&\$18459_w\(31)) & 
                            eclat_if(work.Int.le(\$13921_loop665_arg\(48 to 63), eclat_resize(\$18459_w\(0 to 30),16)) & 
                            work.Int.lt(eclat_resize(\$18459_w\(0 to 30),16), 
                                        work.Int.add(\$13921_loop665_arg\(48 to 63), X"1770")) & eclat_false) & eclat_false);
                if \$v6493\(0) = '1' then
                  \$18447\ := \$18459_w\ & \$13921_loop665_arg\(16 to 31);
                  \$v6480\ := \$ram_lock\;
                  if \$v6480\(0) = '1' then
                    state_var7460 := Q_WAIT6479;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            \$13921_loop665_arg\(64 to 79), \$13921_loop665_arg\(0 to 15))));
                    \$ram_write\ <= \$18447\(0 to 31); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET6478;
                  end if;
                else
                  \$v6492\ := \$ram_lock\;
                  if \$v6492\(0) = '1' then
                    state_var7460 := Q_WAIT6491;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18443\(0 to 30),16)));
                    state_var7460 := PAUSE_GET6490;
                  end if;
                end if;
              when PAUSE_GET6498 =>
                \$18443\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6497\ := work.Bool.lnot(eclat_if(work.Bool.lnot(""&\$18443\(31)) & 
                                           eclat_if(work.Int.le(\$13921_loop665_arg\(32 to 47), eclat_resize(\$18443\(0 to 30),16)) & 
                                           work.Int.lt(eclat_resize(\$18443\(0 to 30),16), 
                                                       work.Int.add(\$13921_loop665_arg\(32 to 47), X"1770")) & eclat_false) & eclat_false));
                if \$v6497\(0) = '1' then
                  \$18447\ := \$18443\ & \$13921_loop665_arg\(16 to 31);
                  \$v6480\ := \$ram_lock\;
                  if \$v6480\(0) = '1' then
                    state_var7460 := Q_WAIT6479;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            \$13921_loop665_arg\(64 to 79), \$13921_loop665_arg\(0 to 15))));
                    \$ram_write\ <= \$18447\(0 to 31); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET6478;
                  end if;
                else
                  \$v6496\ := \$ram_lock\;
                  if \$v6496\(0) = '1' then
                    state_var7460 := Q_WAIT6495;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18443\(0 to 30),16), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6494;
                  end if;
                end if;
              when PAUSE_GET6715 =>
                \$17337\ := \$ram_value\;
                release(\$ram_lock\);
                \$13924_apply638_result\ := eclat_resize(\$17337\(0 to 30),16) & \$13924_apply638_arg\(60 to 91) & \$17333_sp\ & \$13924_apply638_arg\(60 to 91) & \$13924_apply638_arg\(3 to 10) & \$13924_apply638_arg\(150 to 165) & \$13924_apply638_arg\(108 to 109);
                result6468 := \$13924_apply638_result\;
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6740 =>
                \$17368_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$17327\ := \$17368_v\ & work.Int.sub(\$17324\(32 to 47), X"000" & X"1");
                \$v6739\ := ""&\$13924_apply638_arg\(11);
                if \$v6739\(0) = '1' then
                  \$17330_sp\ := work.Int.add(work.Int.sub(\$17327\(32 to 47), \$13924_apply638_arg\(12 to 27)), \$13924_apply638_arg\(28 to 43));
                  \$v6729\ := ""&\$13924_apply638_arg\(2);
                  if \$v6729\(0) = '1' then
                    \$v6728\ := \$ram_lock\;
                    if \$v6728\(0) = '1' then
                      state_var7460 := Q_WAIT6727;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(\$17330_sp\));
                      \$ram_write\ <= \$17327\(0 to 31); \$ram_write_request\ <= '1';
                      state_var7460 := PAUSE_SET6726;
                    end if;
                  else
                    \$17331_sp\ := \$17330_sp\;
                    \$v6725\ := ""&\$13924_apply638_arg\(1);
                    if \$v6725\(0) = '1' then
                      \$v6724\ := \$ram_lock\;
                      if \$v6724\(0) = '1' then
                        state_var7460 := Q_WAIT6723;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr_write\ <= to_integer(unsigned(\$17331_sp\));
                        \$ram_write\ <= \$17324\(0 to 31); \$ram_write_request\ <= '1';
                        state_var7460 := PAUSE_SET6722;
                      end if;
                    else
                      \$17332_sp\ := \$17331_sp\;
                      \$v6721\ := ""&\$13924_apply638_arg\(0);
                      if \$v6721\(0) = '1' then
                        \$v6720\ := \$ram_lock\;
                        if \$v6720\(0) = '1' then
                          state_var7460 := Q_WAIT6719;
                        else
                          acquire(\$ram_lock\);
                          \$ram_ptr_write\ <= to_integer(unsigned(\$17332_sp\));
                          \$ram_write\ <= \$17321\(0 to 31); \$ram_write_request\ <= '1';
                          state_var7460 := PAUSE_SET6718;
                        end if;
                      else
                        \$17333_sp\ := \$17332_sp\;
                        \$v6717\ := \$ram_lock\;
                        if \$v6717\(0) = '1' then
                          state_var7460 := Q_WAIT6716;
                        else
                          acquire(\$ram_lock\);
                          \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                            work.Int.add(
                                                            eclat_resize(\$13924_apply638_arg\(60 to 90),16), X"000" & X"0"), X"000" & X"1")));
                          state_var7460 := PAUSE_GET6715;
                        end if;
                      end if;
                    end if;
                  end if;
                else
                  \$v6738\ := \$ram_lock\;
                  if \$v6738\(0) = '1' then
                    state_var7460 := Q_WAIT6737;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17327\(32 to 47)));
                    \$ram_write\ <= eclat_resize(\$13924_apply638_arg\(142 to 149),31) & eclat_true; \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET6736;
                  end if;
                end if;
              when PAUSE_GET6744 =>
                \$17371_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$17324\ := \$17371_v\ & work.Int.sub(\$17321\(32 to 47), X"000" & X"1");
                \$v6743\ := ""&\$13924_apply638_arg\(2);
                if \$v6743\(0) = '1' then
                  \$v6742\ := \$ram_lock\;
                  if \$v6742\(0) = '1' then
                    state_var7460 := Q_WAIT6741;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$17324\(32 to 47), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6740;
                  end if;
                else
                  \$17327\ := "000"& X"000000" & X"1" & eclat_true & \$17324\(32 to 47);
                  \$v6739\ := ""&\$13924_apply638_arg\(11);
                  if \$v6739\(0) = '1' then
                    \$17330_sp\ := work.Int.add(work.Int.sub(\$17327\(32 to 47), \$13924_apply638_arg\(12 to 27)), \$13924_apply638_arg\(28 to 43));
                    \$v6729\ := ""&\$13924_apply638_arg\(2);
                    if \$v6729\(0) = '1' then
                      \$v6728\ := \$ram_lock\;
                      if \$v6728\(0) = '1' then
                        state_var7460 := Q_WAIT6727;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr_write\ <= to_integer(unsigned(\$17330_sp\));
                        \$ram_write\ <= \$17327\(0 to 31); \$ram_write_request\ <= '1';
                        state_var7460 := PAUSE_SET6726;
                      end if;
                    else
                      \$17331_sp\ := \$17330_sp\;
                      \$v6725\ := ""&\$13924_apply638_arg\(1);
                      if \$v6725\(0) = '1' then
                        \$v6724\ := \$ram_lock\;
                        if \$v6724\(0) = '1' then
                          state_var7460 := Q_WAIT6723;
                        else
                          acquire(\$ram_lock\);
                          \$ram_ptr_write\ <= to_integer(unsigned(\$17331_sp\));
                          \$ram_write\ <= \$17324\(0 to 31); \$ram_write_request\ <= '1';
                          state_var7460 := PAUSE_SET6722;
                        end if;
                      else
                        \$17332_sp\ := \$17331_sp\;
                        \$v6721\ := ""&\$13924_apply638_arg\(0);
                        if \$v6721\(0) = '1' then
                          \$v6720\ := \$ram_lock\;
                          if \$v6720\(0) = '1' then
                            state_var7460 := Q_WAIT6719;
                          else
                            acquire(\$ram_lock\);
                            \$ram_ptr_write\ <= to_integer(unsigned(\$17332_sp\));
                            \$ram_write\ <= \$17321\(0 to 31); \$ram_write_request\ <= '1';
                            state_var7460 := PAUSE_SET6718;
                          end if;
                        else
                          \$17333_sp\ := \$17332_sp\;
                          \$v6717\ := \$ram_lock\;
                          if \$v6717\(0) = '1' then
                            state_var7460 := Q_WAIT6716;
                          else
                            acquire(\$ram_lock\);
                            \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                              work.Int.add(
                                                              eclat_resize(\$13924_apply638_arg\(60 to 90),16), X"000" & X"0"), X"000" & X"1")));
                            state_var7460 := PAUSE_GET6715;
                          end if;
                        end if;
                      end if;
                    end if;
                  else
                    \$v6738\ := \$ram_lock\;
                    if \$v6738\(0) = '1' then
                      state_var7460 := Q_WAIT6737;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(\$17327\(32 to 47)));
                      \$ram_write\ <= eclat_resize(\$13924_apply638_arg\(142 to 149),31) & eclat_true; \$ram_write_request\ <= '1';
                      state_var7460 := PAUSE_SET6736;
                    end if;
                  end if;
                end if;
              when PAUSE_GET6748 =>
                \$17374_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$17321\ := \$17374_v\ & work.Int.sub(\$13924_apply638_arg\(92 to 107), X"000" & X"1");
                \$v6747\ := ""&\$13924_apply638_arg\(1);
                if \$v6747\(0) = '1' then
                  \$v6746\ := \$ram_lock\;
                  if \$v6746\(0) = '1' then
                    state_var7460 := Q_WAIT6745;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$17321\(32 to 47), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6744;
                  end if;
                else
                  \$17324\ := "000"& X"000000" & X"1" & eclat_true & \$17321\(32 to 47);
                  \$v6743\ := ""&\$13924_apply638_arg\(2);
                  if \$v6743\(0) = '1' then
                    \$v6742\ := \$ram_lock\;
                    if \$v6742\(0) = '1' then
                      state_var7460 := Q_WAIT6741;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(
                                                        \$17324\(32 to 47), X"000" & X"1")));
                      state_var7460 := PAUSE_GET6740;
                    end if;
                  else
                    \$17327\ := "000"& X"000000" & X"1" & eclat_true & \$17324\(32 to 47);
                    \$v6739\ := ""&\$13924_apply638_arg\(11);
                    if \$v6739\(0) = '1' then
                      \$17330_sp\ := work.Int.add(work.Int.sub(\$17327\(32 to 47), \$13924_apply638_arg\(12 to 27)), \$13924_apply638_arg\(28 to 43));
                      \$v6729\ := ""&\$13924_apply638_arg\(2);
                      if \$v6729\(0) = '1' then
                        \$v6728\ := \$ram_lock\;
                        if \$v6728\(0) = '1' then
                          state_var7460 := Q_WAIT6727;
                        else
                          acquire(\$ram_lock\);
                          \$ram_ptr_write\ <= to_integer(unsigned(\$17330_sp\));
                          \$ram_write\ <= \$17327\(0 to 31); \$ram_write_request\ <= '1';
                          state_var7460 := PAUSE_SET6726;
                        end if;
                      else
                        \$17331_sp\ := \$17330_sp\;
                        \$v6725\ := ""&\$13924_apply638_arg\(1);
                        if \$v6725\(0) = '1' then
                          \$v6724\ := \$ram_lock\;
                          if \$v6724\(0) = '1' then
                            state_var7460 := Q_WAIT6723;
                          else
                            acquire(\$ram_lock\);
                            \$ram_ptr_write\ <= to_integer(unsigned(\$17331_sp\));
                            \$ram_write\ <= \$17324\(0 to 31); \$ram_write_request\ <= '1';
                            state_var7460 := PAUSE_SET6722;
                          end if;
                        else
                          \$17332_sp\ := \$17331_sp\;
                          \$v6721\ := ""&\$13924_apply638_arg\(0);
                          if \$v6721\(0) = '1' then
                            \$v6720\ := \$ram_lock\;
                            if \$v6720\(0) = '1' then
                              state_var7460 := Q_WAIT6719;
                            else
                              acquire(\$ram_lock\);
                              \$ram_ptr_write\ <= to_integer(unsigned(\$17332_sp\));
                              \$ram_write\ <= \$17321\(0 to 31); \$ram_write_request\ <= '1';
                              state_var7460 := PAUSE_SET6718;
                            end if;
                          else
                            \$17333_sp\ := \$17332_sp\;
                            \$v6717\ := \$ram_lock\;
                            if \$v6717\(0) = '1' then
                              state_var7460 := Q_WAIT6716;
                            else
                              acquire(\$ram_lock\);
                              \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                                work.Int.add(
                                                                eclat_resize(\$13924_apply638_arg\(60 to 90),16), X"000" & X"0"), X"000" & X"1")));
                              state_var7460 := PAUSE_GET6715;
                            end if;
                          end if;
                        end if;
                      end if;
                    else
                      \$v6738\ := \$ram_lock\;
                      if \$v6738\(0) = '1' then
                        state_var7460 := Q_WAIT6737;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr_write\ <= to_integer(unsigned(\$17327\(32 to 47)));
                        \$ram_write\ <= eclat_resize(\$13924_apply638_arg\(142 to 149),31) & eclat_true; \$ram_write_request\ <= '1';
                        state_var7460 := PAUSE_SET6736;
                      end if;
                    end if;
                  end if;
                end if;
              when PAUSE_GET6756 =>
                \$17239_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6755\ := \$ram_lock\;
                if \$v6755\(0) = '1' then
                  state_var7460 := Q_WAIT6754;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$17232\(64 to 94),16), X"000" & X"2"), X"000" & X"1")));
                  \$ram_write\ <= \$17239_v\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6753;
                end if;
              when PAUSE_GET6763 =>
                \$17250_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6762\ := \$ram_lock\;
                if \$v6762\(0) = '1' then
                  state_var7460 := Q_WAIT6761;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$17232\(64 to 94),16), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= \$17250_v\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6760;
                end if;
              when PAUSE_GET6771 =>
                \$17207_arg\ := \$code_value\;
                release(\$code_lock\);
                \$13927_branch_if648_result\ := work.Int.add(work.Int.add(
                                                             \$13927_branch_if648_arg\(1 to 16), X"000" & X"1"), eclat_resize(\$17207_arg\,16)) & \$13927_branch_if648_arg\(17 to 48) & \$13927_branch_if648_arg\(49 to 64) & \$13927_branch_if648_arg\(65 to 120) & \$13927_branch_if648_arg\(121 to 122);
                result6468 := \$13927_branch_if648_result\;
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6778 =>
                \$17183\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6777\ := \$ram_lock\;
                if \$v6777\(0) = '1' then
                  state_var7460 := Q_WAIT6776;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.sub(
                                                          work.Int.sub(
                                                          work.Int.sub(
                                                          \$13928_w652_arg\(16 to 31), \$13928_w652_arg\(32 to 47)), \$13928_w652_arg\(48 to 63)), \$13928_w652_arg\(0 to 15))));
                  \$ram_write\ <= \$17183\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6775;
                end if;
              when PAUSE_GET6782 =>
                \$13967_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$13967_v\ & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6785 =>
                \$13972_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$13972_v\ & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6788 =>
                \$13977_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$13977_v\ & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6791 =>
                \$13982_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$13982_v\ & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6794 =>
                \$13987_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$13987_v\ & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6797 =>
                \$13992_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$13992_v\ & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6800 =>
                \$13997_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$13997_v\ & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6803 =>
                \$14002_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$14002_v\ & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6812 =>
                \$14016_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$14016_v\ & 
                work.Int.add(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6818 =>
                \$14025_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$14025_v\ & 
                work.Int.add(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6824 =>
                \$14034_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$14034_v\ & 
                work.Int.add(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6830 =>
                \$14043_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$14043_v\ & 
                work.Int.add(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6836 =>
                \$14052_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$14052_v\ & 
                work.Int.add(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6842 =>
                \$14061_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$14061_v\ & 
                work.Int.add(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6848 =>
                \$14070_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$14070_v\ & 
                work.Int.add(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6854 =>
                \$14081\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$14081\ & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6857 =>
                \$14092\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$14092\ & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6860 =>
                \$14103\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$14103\ & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6863 =>
                \$14114\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$14114\ & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6866 =>
                \$14126\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$14126\ & 
                work.Int.add(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6872 =>
                \$14139\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$14139\ & 
                work.Int.add(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6878 =>
                \$14152\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$14152\ & 
                work.Int.add(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6884 =>
                \$14165\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$14165\ & 
                work.Int.add(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6890 =>
                \$14185_next_env\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$13911\(16 to 47) & \$14181_sp\ & \$14185_next_env\ & 
                work.Int.add(\$13911\(96 to 103), work.Int.sub(eclat_resize(eclat_resize(
                                                               work.Int.lsr(
                                                               eclat_resize(eclat_resize(\$14177_hd\(0 to 30),16),31), X"0000000" & X"2"),16),8), "00000010")) & \$13911\(104 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6896 =>
                \$14221\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6895\ := \$ram_lock\;
                if \$v6895\(0) = '1' then
                  state_var7460 := Q_WAIT6894;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$14207_loop_push6495899_arg\(0 to 15)));
                  \$ram_write\ <= \$14221\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6893;
                end if;
              when PAUSE_GET6900 =>
                \$14177_hd\ := \$ram_value\;
                release(\$ram_lock\);
                \$14207_loop_push6495899_id\ := "000000111000";
                \$14207_loop_push6495899_arg\ := \$13911\(48 to 63) & "00000000" & \$13911\(64 to 95) & eclat_resize(eclat_resize(
                work.Int.lsr(eclat_resize(eclat_resize(\$14177_hd\(0 to 30),16),31), X"0000000" & X"2"),16),8);
                state_var7460 := \$14207_LOOP_PUSH6495899\;
              when PAUSE_GET6915 =>
                \$14285_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$14285_v\ & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6918 =>
                \$14300_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$14300_v\ & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6921 =>
                \$14315_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$14315_v\ & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6924 =>
                \$14330_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$14330_v\ & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6930 =>
                \$14338_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6929\ := \$ram_lock\;
                if \$v6929\(0) = '1' then
                  state_var7460 := Q_WAIT6928;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$13911\(16 to 46),16), X"000" & X"0"), X"000" & X"1")));
                  \$ram_write\ <= \$14338_v\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6927;
                end if;
              when PAUSE_GET6936 =>
                \$14351_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6935\ := \$ram_lock\;
                if \$v6935\(0) = '1' then
                  state_var7460 := Q_WAIT6934;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$13911\(16 to 46),16), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= \$14351_v\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6933;
                end if;
              when PAUSE_GET6942 =>
                \$14364_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6941\ := \$ram_lock\;
                if \$v6941\(0) = '1' then
                  state_var7460 := Q_WAIT6940;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$13911\(16 to 46),16), X"000" & X"2"), X"000" & X"1")));
                  \$ram_write\ <= \$14364_v\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6939;
                end if;
              when PAUSE_GET6948 =>
                \$14377_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6947\ := \$ram_lock\;
                if \$v6947\(0) = '1' then
                  state_var7460 := Q_WAIT6946;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$13911\(16 to 46),16), X"000" & X"3"), X"000" & X"1")));
                  \$ram_write\ <= \$14377_v\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6945;
                end if;
              when PAUSE_GET6951 =>
                \$14393_hd\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & eclat_resize(eclat_resize(
                work.Int.lsr(eclat_resize(eclat_resize(\$14393_hd\(0 to 30),16),31), X"0000000" & X"2"),16),31) & eclat_true & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6954 =>
                \$14413_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$14413_v\ & 
                work.Int.sub(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6957 =>
                \$14406_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6956\ := \$ram_lock\;
                if \$v6956\(0) = '1' then
                  state_var7460 := Q_WAIT6955;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13911\(16 to 46),16), eclat_resize(\$14406_v\(0 to 30),16)), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6954;
                end if;
              when PAUSE_GET6963 =>
                \$14424_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6962\ := \$ram_lock\;
                if \$v6962\(0) = '1' then
                  state_var7460 := Q_WAIT6961;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$13911\(16 to 46),16), eclat_resize(\$14423_v\(0 to 30),16)), X"000" & X"1")));
                  \$ram_write\ <= \$14424_v\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6960;
                end if;
              when PAUSE_GET6966 =>
                \$14423_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6965\ := \$ram_lock\;
                if \$v6965\(0) = '1' then
                  state_var7460 := Q_WAIT6964;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6963;
                end if;
              when PAUSE_GET6969 =>
                \$14453_next_acc\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$14453_next_acc\ & 
                work.Int.sub(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6972 =>
                \$14446_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6971\ := \$ram_lock\;
                if \$v6971\(0) = '1' then
                  state_var7460 := Q_WAIT6970;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13911\(16 to 46),16), eclat_resize(\$14446_v\(0 to 30),16)), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6969;
                end if;
              when PAUSE_GET6978 =>
                \$14464_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6977\ := \$ram_lock\;
                if \$v6977\(0) = '1' then
                  state_var7460 := Q_WAIT6976;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$13911\(16 to 46),16), eclat_resize(\$14463_v\(0 to 30),16)), X"000" & X"1")));
                  \$ram_write\ <= \$14464_v\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6975;
                end if;
              when PAUSE_GET6981 =>
                \$14463_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6980\ := \$ram_lock\;
                if \$v6980\(0) = '1' then
                  state_var7460 := Q_WAIT6979;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6978;
                end if;
              when PAUSE_GET6984 =>
                \$14493_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$13911\(16 to 47) & 
                work.Int.sub(work.Int.sub(work.Int.sub(\$13911\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"2") & \$13911\(64 to 95) & \$13911\(96 to 103) & eclat_resize(\$14493_v\(0 to 30),16) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6987 =>
                \$14517_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := eclat_resize(\$14508_v\(0 to 30),16) & \$13911\(16 to 47) & 
                work.Int.sub(work.Int.sub(work.Int.sub(work.Int.sub(\$13911\(104 to 119), X"000" & X"1"), X"000" & X"1"), X"000" & X"1"), X"000" & X"1") & \$14516_v\ & eclat_resize(\$14517_v\(0 to 30),8) & eclat_resize(\$14512_v\(0 to 30),16) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET6990 =>
                \$14516_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6989\ := \$ram_lock\;
                if \$v6989\(0) = '1' then
                  state_var7460 := Q_WAIT6988;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$13911\(104 to 119), X"000" & X"1"), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6987;
                end if;
              when PAUSE_GET6993 =>
                \$14512_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6992\ := \$ram_lock\;
                if \$v6992\(0) = '1' then
                  state_var7460 := Q_WAIT6991;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$13911\(104 to 119), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6990;
                end if;
              when PAUSE_GET6996 =>
                \$14508_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v6995\ := \$ram_lock\;
                if \$v6995\(0) = '1' then
                  state_var7460 := Q_WAIT6994;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$13911\(104 to 119), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6993;
                end if;
              when PAUSE_GET7018 =>
                \$14578_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7017\ := \$14564_binop_int6435900_arg\(0 to 31);
                case \$v7017\ is
                when X"0000000" & X"0" =>
                  \$14582_res\ := work.Int.add(\$14564_binop_int6435900_arg\(48 to 78), \$14578_v\(0 to 30));
                  \$14564_binop_int6435900_result\ := work.Int.add(\$14564_binop_int6435900_arg\(32 to 47), X"000" & X"1") & \$14582_res\ & eclat_true & 
                  work.Int.sub(\$14564_binop_int6435900_arg\(80 to 95), X"000" & X"1") & \$14564_binop_int6435900_arg\(96 to 151) & \$14564_binop_int6435900_arg\(152 to 153);
                  result6468 := \$14564_binop_int6435900_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"1" =>
                  \$14582_res\ := work.Int.sub(\$14564_binop_int6435900_arg\(48 to 78), \$14578_v\(0 to 30));
                  \$14564_binop_int6435900_result\ := work.Int.add(\$14564_binop_int6435900_arg\(32 to 47), X"000" & X"1") & \$14582_res\ & eclat_true & 
                  work.Int.sub(\$14564_binop_int6435900_arg\(80 to 95), X"000" & X"1") & \$14564_binop_int6435900_arg\(96 to 151) & \$14564_binop_int6435900_arg\(152 to 153);
                  result6468 := \$14564_binop_int6435900_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"2" =>
                  \$14582_res\ := work.Int.mul(\$14564_binop_int6435900_arg\(48 to 78), \$14578_v\(0 to 30));
                  \$14564_binop_int6435900_result\ := work.Int.add(\$14564_binop_int6435900_arg\(32 to 47), X"000" & X"1") & \$14582_res\ & eclat_true & 
                  work.Int.sub(\$14564_binop_int6435900_arg\(80 to 95), X"000" & X"1") & \$14564_binop_int6435900_arg\(96 to 151) & \$14564_binop_int6435900_arg\(152 to 153);
                  result6468 := \$14564_binop_int6435900_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"3" =>
                  \$v7013\ := work.Int.eq(\$14578_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v7013\(0) = '1' then
                    \$14582_res\ := "000"& X"000000" & X"0";
                    \$14564_binop_int6435900_result\ := work.Int.add(
                                                        \$14564_binop_int6435900_arg\(32 to 47), X"000" & X"1") & \$14582_res\ & eclat_true & 
                    work.Int.sub(\$14564_binop_int6435900_arg\(80 to 95), X"000" & X"1") & \$14564_binop_int6435900_arg\(96 to 151) & \$14564_binop_int6435900_arg\(152 to 153);
                    result6468 := \$14564_binop_int6435900_result\;
                    rdy6469 := eclat_true;
                    state_var7460 := IDLE6470;
                  else
                    \$14589_modulo6685895_id\ := "000001000100";
                    \$14589_modulo6685895_arg\ := work.Int.absv(\$14564_binop_int6435900_arg\(48 to 78)) & 
                    work.Int.absv(\$14578_v\(0 to 30));
                    state_var7460 := \$14589_MODULO6685895\;
                  end if;
                when X"0000000" & X"4" =>
                  \$v7016\ := work.Int.eq(\$14578_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v7016\(0) = '1' then
                    \$14582_res\ := "000"& X"000000" & X"0";
                    \$14564_binop_int6435900_result\ := work.Int.add(
                                                        \$14564_binop_int6435900_arg\(32 to 47), X"000" & X"1") & \$14582_res\ & eclat_true & 
                    work.Int.sub(\$14564_binop_int6435900_arg\(80 to 95), X"000" & X"1") & \$14564_binop_int6435900_arg\(96 to 151) & \$14564_binop_int6435900_arg\(152 to 153);
                    result6468 := \$14564_binop_int6435900_result\;
                    rdy6469 := eclat_true;
                    state_var7460 := IDLE6470;
                  else
                    \$14613_modulo6685896_id\ := "000001000110";
                    \$14613_modulo6685896_arg\ := work.Int.absv(\$14564_binop_int6435900_arg\(48 to 78)) & 
                    work.Int.absv(\$14578_v\(0 to 30));
                    state_var7460 := \$14613_MODULO6685896\;
                  end if;
                when X"0000000" & X"5" =>
                  \$14582_res\ := work.Int.land(\$14564_binop_int6435900_arg\(48 to 78), \$14578_v\(0 to 30));
                  \$14564_binop_int6435900_result\ := work.Int.add(\$14564_binop_int6435900_arg\(32 to 47), X"000" & X"1") & \$14582_res\ & eclat_true & 
                  work.Int.sub(\$14564_binop_int6435900_arg\(80 to 95), X"000" & X"1") & \$14564_binop_int6435900_arg\(96 to 151) & \$14564_binop_int6435900_arg\(152 to 153);
                  result6468 := \$14564_binop_int6435900_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"6" =>
                  \$14582_res\ := work.Int.lor(\$14564_binop_int6435900_arg\(48 to 78), \$14578_v\(0 to 30));
                  \$14564_binop_int6435900_result\ := work.Int.add(\$14564_binop_int6435900_arg\(32 to 47), X"000" & X"1") & \$14582_res\ & eclat_true & 
                  work.Int.sub(\$14564_binop_int6435900_arg\(80 to 95), X"000" & X"1") & \$14564_binop_int6435900_arg\(96 to 151) & \$14564_binop_int6435900_arg\(152 to 153);
                  result6468 := \$14564_binop_int6435900_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"7" =>
                  \$14582_res\ := work.Int.lxor(\$14564_binop_int6435900_arg\(48 to 78), \$14578_v\(0 to 30));
                  \$14564_binop_int6435900_result\ := work.Int.add(\$14564_binop_int6435900_arg\(32 to 47), X"000" & X"1") & \$14582_res\ & eclat_true & 
                  work.Int.sub(\$14564_binop_int6435900_arg\(80 to 95), X"000" & X"1") & \$14564_binop_int6435900_arg\(96 to 151) & \$14564_binop_int6435900_arg\(152 to 153);
                  result6468 := \$14564_binop_int6435900_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"8" =>
                  \$14582_res\ := work.Int.lsl(\$14564_binop_int6435900_arg\(48 to 78), \$14578_v\(0 to 30));
                  \$14564_binop_int6435900_result\ := work.Int.add(\$14564_binop_int6435900_arg\(32 to 47), X"000" & X"1") & \$14582_res\ & eclat_true & 
                  work.Int.sub(\$14564_binop_int6435900_arg\(80 to 95), X"000" & X"1") & \$14564_binop_int6435900_arg\(96 to 151) & \$14564_binop_int6435900_arg\(152 to 153);
                  result6468 := \$14564_binop_int6435900_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"9" =>
                  \$14582_res\ := work.Int.lsr(\$14564_binop_int6435900_arg\(48 to 78), \$14578_v\(0 to 30));
                  \$14564_binop_int6435900_result\ := work.Int.add(\$14564_binop_int6435900_arg\(32 to 47), X"000" & X"1") & \$14582_res\ & eclat_true & 
                  work.Int.sub(\$14564_binop_int6435900_arg\(80 to 95), X"000" & X"1") & \$14564_binop_int6435900_arg\(96 to 151) & \$14564_binop_int6435900_arg\(152 to 153);
                  result6468 := \$14564_binop_int6435900_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"a" =>
                  \$14582_res\ := work.Int.asr(\$14564_binop_int6435900_arg\(48 to 78), \$14578_v\(0 to 30));
                  \$14564_binop_int6435900_result\ := work.Int.add(\$14564_binop_int6435900_arg\(32 to 47), X"000" & X"1") & \$14582_res\ & eclat_true & 
                  work.Int.sub(\$14564_binop_int6435900_arg\(80 to 95), X"000" & X"1") & \$14564_binop_int6435900_arg\(96 to 151) & \$14564_binop_int6435900_arg\(152 to 153);
                  result6468 := \$14564_binop_int6435900_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"b" =>
                  \$14582_res\ := eclat_if(work.Int.lt(\$14564_binop_int6435900_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$14578_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.gt(\$14564_binop_int6435900_arg\(48 to 78), \$14578_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$14578_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"0" & 
                                  eclat_if(work.Int.lt(\$14564_binop_int6435900_arg\(48 to 78), \$14578_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$14564_binop_int6435900_result\ := work.Int.add(\$14564_binop_int6435900_arg\(32 to 47), X"000" & X"1") & \$14582_res\ & eclat_true & 
                  work.Int.sub(\$14564_binop_int6435900_arg\(80 to 95), X"000" & X"1") & \$14564_binop_int6435900_arg\(96 to 151) & \$14564_binop_int6435900_arg\(152 to 153);
                  result6468 := \$14564_binop_int6435900_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"c" =>
                  \$14582_res\ := eclat_if(work.Int.lt(\$14564_binop_int6435900_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$14578_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.le(\$14564_binop_int6435900_arg\(48 to 78), \$14578_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"1") & 
                                  eclat_if(work.Int.lt(\$14578_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & 
                                  eclat_if(work.Int.ge(\$14564_binop_int6435900_arg\(48 to 78), \$14578_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$14564_binop_int6435900_result\ := work.Int.add(\$14564_binop_int6435900_arg\(32 to 47), X"000" & X"1") & \$14582_res\ & eclat_true & 
                  work.Int.sub(\$14564_binop_int6435900_arg\(80 to 95), X"000" & X"1") & \$14564_binop_int6435900_arg\(96 to 151) & \$14564_binop_int6435900_arg\(152 to 153);
                  result6468 := \$14564_binop_int6435900_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when others =>
                  \$14582_res\ := "000"& X"000000" & X"0";
                  \$14564_binop_int6435900_result\ := work.Int.add(\$14564_binop_int6435900_arg\(32 to 47), X"000" & X"1") & \$14582_res\ & eclat_true & 
                  work.Int.sub(\$14564_binop_int6435900_arg\(80 to 95), X"000" & X"1") & \$14564_binop_int6435900_arg\(96 to 151) & \$14564_binop_int6435900_arg\(152 to 153);
                  result6468 := \$14564_binop_int6435900_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                end case;
              when PAUSE_GET7028 =>
                \$14658_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7027\ := \$14644_binop_int6435901_arg\(0 to 31);
                case \$v7027\ is
                when X"0000000" & X"0" =>
                  \$14662_res\ := work.Int.add(\$14644_binop_int6435901_arg\(48 to 78), \$14658_v\(0 to 30));
                  \$14644_binop_int6435901_result\ := work.Int.add(\$14644_binop_int6435901_arg\(32 to 47), X"000" & X"1") & \$14662_res\ & eclat_true & 
                  work.Int.sub(\$14644_binop_int6435901_arg\(80 to 95), X"000" & X"1") & \$14644_binop_int6435901_arg\(96 to 151) & \$14644_binop_int6435901_arg\(152 to 153);
                  result6468 := \$14644_binop_int6435901_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"1" =>
                  \$14662_res\ := work.Int.sub(\$14644_binop_int6435901_arg\(48 to 78), \$14658_v\(0 to 30));
                  \$14644_binop_int6435901_result\ := work.Int.add(\$14644_binop_int6435901_arg\(32 to 47), X"000" & X"1") & \$14662_res\ & eclat_true & 
                  work.Int.sub(\$14644_binop_int6435901_arg\(80 to 95), X"000" & X"1") & \$14644_binop_int6435901_arg\(96 to 151) & \$14644_binop_int6435901_arg\(152 to 153);
                  result6468 := \$14644_binop_int6435901_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"2" =>
                  \$14662_res\ := work.Int.mul(\$14644_binop_int6435901_arg\(48 to 78), \$14658_v\(0 to 30));
                  \$14644_binop_int6435901_result\ := work.Int.add(\$14644_binop_int6435901_arg\(32 to 47), X"000" & X"1") & \$14662_res\ & eclat_true & 
                  work.Int.sub(\$14644_binop_int6435901_arg\(80 to 95), X"000" & X"1") & \$14644_binop_int6435901_arg\(96 to 151) & \$14644_binop_int6435901_arg\(152 to 153);
                  result6468 := \$14644_binop_int6435901_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"3" =>
                  \$v7023\ := work.Int.eq(\$14658_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v7023\(0) = '1' then
                    \$14662_res\ := "000"& X"000000" & X"0";
                    \$14644_binop_int6435901_result\ := work.Int.add(
                                                        \$14644_binop_int6435901_arg\(32 to 47), X"000" & X"1") & \$14662_res\ & eclat_true & 
                    work.Int.sub(\$14644_binop_int6435901_arg\(80 to 95), X"000" & X"1") & \$14644_binop_int6435901_arg\(96 to 151) & \$14644_binop_int6435901_arg\(152 to 153);
                    result6468 := \$14644_binop_int6435901_result\;
                    rdy6469 := eclat_true;
                    state_var7460 := IDLE6470;
                  else
                    \$14669_modulo6685895_id\ := "000001001001";
                    \$14669_modulo6685895_arg\ := work.Int.absv(\$14644_binop_int6435901_arg\(48 to 78)) & 
                    work.Int.absv(\$14658_v\(0 to 30));
                    state_var7460 := \$14669_MODULO6685895\;
                  end if;
                when X"0000000" & X"4" =>
                  \$v7026\ := work.Int.eq(\$14658_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v7026\(0) = '1' then
                    \$14662_res\ := "000"& X"000000" & X"0";
                    \$14644_binop_int6435901_result\ := work.Int.add(
                                                        \$14644_binop_int6435901_arg\(32 to 47), X"000" & X"1") & \$14662_res\ & eclat_true & 
                    work.Int.sub(\$14644_binop_int6435901_arg\(80 to 95), X"000" & X"1") & \$14644_binop_int6435901_arg\(96 to 151) & \$14644_binop_int6435901_arg\(152 to 153);
                    result6468 := \$14644_binop_int6435901_result\;
                    rdy6469 := eclat_true;
                    state_var7460 := IDLE6470;
                  else
                    \$14693_modulo6685896_id\ := "000001001011";
                    \$14693_modulo6685896_arg\ := work.Int.absv(\$14644_binop_int6435901_arg\(48 to 78)) & 
                    work.Int.absv(\$14658_v\(0 to 30));
                    state_var7460 := \$14693_MODULO6685896\;
                  end if;
                when X"0000000" & X"5" =>
                  \$14662_res\ := work.Int.land(\$14644_binop_int6435901_arg\(48 to 78), \$14658_v\(0 to 30));
                  \$14644_binop_int6435901_result\ := work.Int.add(\$14644_binop_int6435901_arg\(32 to 47), X"000" & X"1") & \$14662_res\ & eclat_true & 
                  work.Int.sub(\$14644_binop_int6435901_arg\(80 to 95), X"000" & X"1") & \$14644_binop_int6435901_arg\(96 to 151) & \$14644_binop_int6435901_arg\(152 to 153);
                  result6468 := \$14644_binop_int6435901_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"6" =>
                  \$14662_res\ := work.Int.lor(\$14644_binop_int6435901_arg\(48 to 78), \$14658_v\(0 to 30));
                  \$14644_binop_int6435901_result\ := work.Int.add(\$14644_binop_int6435901_arg\(32 to 47), X"000" & X"1") & \$14662_res\ & eclat_true & 
                  work.Int.sub(\$14644_binop_int6435901_arg\(80 to 95), X"000" & X"1") & \$14644_binop_int6435901_arg\(96 to 151) & \$14644_binop_int6435901_arg\(152 to 153);
                  result6468 := \$14644_binop_int6435901_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"7" =>
                  \$14662_res\ := work.Int.lxor(\$14644_binop_int6435901_arg\(48 to 78), \$14658_v\(0 to 30));
                  \$14644_binop_int6435901_result\ := work.Int.add(\$14644_binop_int6435901_arg\(32 to 47), X"000" & X"1") & \$14662_res\ & eclat_true & 
                  work.Int.sub(\$14644_binop_int6435901_arg\(80 to 95), X"000" & X"1") & \$14644_binop_int6435901_arg\(96 to 151) & \$14644_binop_int6435901_arg\(152 to 153);
                  result6468 := \$14644_binop_int6435901_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"8" =>
                  \$14662_res\ := work.Int.lsl(\$14644_binop_int6435901_arg\(48 to 78), \$14658_v\(0 to 30));
                  \$14644_binop_int6435901_result\ := work.Int.add(\$14644_binop_int6435901_arg\(32 to 47), X"000" & X"1") & \$14662_res\ & eclat_true & 
                  work.Int.sub(\$14644_binop_int6435901_arg\(80 to 95), X"000" & X"1") & \$14644_binop_int6435901_arg\(96 to 151) & \$14644_binop_int6435901_arg\(152 to 153);
                  result6468 := \$14644_binop_int6435901_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"9" =>
                  \$14662_res\ := work.Int.lsr(\$14644_binop_int6435901_arg\(48 to 78), \$14658_v\(0 to 30));
                  \$14644_binop_int6435901_result\ := work.Int.add(\$14644_binop_int6435901_arg\(32 to 47), X"000" & X"1") & \$14662_res\ & eclat_true & 
                  work.Int.sub(\$14644_binop_int6435901_arg\(80 to 95), X"000" & X"1") & \$14644_binop_int6435901_arg\(96 to 151) & \$14644_binop_int6435901_arg\(152 to 153);
                  result6468 := \$14644_binop_int6435901_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"a" =>
                  \$14662_res\ := work.Int.asr(\$14644_binop_int6435901_arg\(48 to 78), \$14658_v\(0 to 30));
                  \$14644_binop_int6435901_result\ := work.Int.add(\$14644_binop_int6435901_arg\(32 to 47), X"000" & X"1") & \$14662_res\ & eclat_true & 
                  work.Int.sub(\$14644_binop_int6435901_arg\(80 to 95), X"000" & X"1") & \$14644_binop_int6435901_arg\(96 to 151) & \$14644_binop_int6435901_arg\(152 to 153);
                  result6468 := \$14644_binop_int6435901_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"b" =>
                  \$14662_res\ := eclat_if(work.Int.lt(\$14644_binop_int6435901_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$14658_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.gt(\$14644_binop_int6435901_arg\(48 to 78), \$14658_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$14658_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"0" & 
                                  eclat_if(work.Int.lt(\$14644_binop_int6435901_arg\(48 to 78), \$14658_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$14644_binop_int6435901_result\ := work.Int.add(\$14644_binop_int6435901_arg\(32 to 47), X"000" & X"1") & \$14662_res\ & eclat_true & 
                  work.Int.sub(\$14644_binop_int6435901_arg\(80 to 95), X"000" & X"1") & \$14644_binop_int6435901_arg\(96 to 151) & \$14644_binop_int6435901_arg\(152 to 153);
                  result6468 := \$14644_binop_int6435901_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"c" =>
                  \$14662_res\ := eclat_if(work.Int.lt(\$14644_binop_int6435901_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$14658_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.le(\$14644_binop_int6435901_arg\(48 to 78), \$14658_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"1") & 
                                  eclat_if(work.Int.lt(\$14658_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & 
                                  eclat_if(work.Int.ge(\$14644_binop_int6435901_arg\(48 to 78), \$14658_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$14644_binop_int6435901_result\ := work.Int.add(\$14644_binop_int6435901_arg\(32 to 47), X"000" & X"1") & \$14662_res\ & eclat_true & 
                  work.Int.sub(\$14644_binop_int6435901_arg\(80 to 95), X"000" & X"1") & \$14644_binop_int6435901_arg\(96 to 151) & \$14644_binop_int6435901_arg\(152 to 153);
                  result6468 := \$14644_binop_int6435901_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when others =>
                  \$14662_res\ := "000"& X"000000" & X"0";
                  \$14644_binop_int6435901_result\ := work.Int.add(\$14644_binop_int6435901_arg\(32 to 47), X"000" & X"1") & \$14662_res\ & eclat_true & 
                  work.Int.sub(\$14644_binop_int6435901_arg\(80 to 95), X"000" & X"1") & \$14644_binop_int6435901_arg\(96 to 151) & \$14644_binop_int6435901_arg\(152 to 153);
                  result6468 := \$14644_binop_int6435901_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                end case;
              when PAUSE_GET7038 =>
                \$14738_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7037\ := \$14724_binop_int6435902_arg\(0 to 31);
                case \$v7037\ is
                when X"0000000" & X"0" =>
                  \$14742_res\ := work.Int.add(\$14724_binop_int6435902_arg\(48 to 78), \$14738_v\(0 to 30));
                  \$14724_binop_int6435902_result\ := work.Int.add(\$14724_binop_int6435902_arg\(32 to 47), X"000" & X"1") & \$14742_res\ & eclat_true & 
                  work.Int.sub(\$14724_binop_int6435902_arg\(80 to 95), X"000" & X"1") & \$14724_binop_int6435902_arg\(96 to 151) & \$14724_binop_int6435902_arg\(152 to 153);
                  result6468 := \$14724_binop_int6435902_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"1" =>
                  \$14742_res\ := work.Int.sub(\$14724_binop_int6435902_arg\(48 to 78), \$14738_v\(0 to 30));
                  \$14724_binop_int6435902_result\ := work.Int.add(\$14724_binop_int6435902_arg\(32 to 47), X"000" & X"1") & \$14742_res\ & eclat_true & 
                  work.Int.sub(\$14724_binop_int6435902_arg\(80 to 95), X"000" & X"1") & \$14724_binop_int6435902_arg\(96 to 151) & \$14724_binop_int6435902_arg\(152 to 153);
                  result6468 := \$14724_binop_int6435902_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"2" =>
                  \$14742_res\ := work.Int.mul(\$14724_binop_int6435902_arg\(48 to 78), \$14738_v\(0 to 30));
                  \$14724_binop_int6435902_result\ := work.Int.add(\$14724_binop_int6435902_arg\(32 to 47), X"000" & X"1") & \$14742_res\ & eclat_true & 
                  work.Int.sub(\$14724_binop_int6435902_arg\(80 to 95), X"000" & X"1") & \$14724_binop_int6435902_arg\(96 to 151) & \$14724_binop_int6435902_arg\(152 to 153);
                  result6468 := \$14724_binop_int6435902_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"3" =>
                  \$v7033\ := work.Int.eq(\$14738_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v7033\(0) = '1' then
                    \$14742_res\ := "000"& X"000000" & X"0";
                    \$14724_binop_int6435902_result\ := work.Int.add(
                                                        \$14724_binop_int6435902_arg\(32 to 47), X"000" & X"1") & \$14742_res\ & eclat_true & 
                    work.Int.sub(\$14724_binop_int6435902_arg\(80 to 95), X"000" & X"1") & \$14724_binop_int6435902_arg\(96 to 151) & \$14724_binop_int6435902_arg\(152 to 153);
                    result6468 := \$14724_binop_int6435902_result\;
                    rdy6469 := eclat_true;
                    state_var7460 := IDLE6470;
                  else
                    \$14749_modulo6685895_id\ := "000001001110";
                    \$14749_modulo6685895_arg\ := work.Int.absv(\$14724_binop_int6435902_arg\(48 to 78)) & 
                    work.Int.absv(\$14738_v\(0 to 30));
                    state_var7460 := \$14749_MODULO6685895\;
                  end if;
                when X"0000000" & X"4" =>
                  \$v7036\ := work.Int.eq(\$14738_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v7036\(0) = '1' then
                    \$14742_res\ := "000"& X"000000" & X"0";
                    \$14724_binop_int6435902_result\ := work.Int.add(
                                                        \$14724_binop_int6435902_arg\(32 to 47), X"000" & X"1") & \$14742_res\ & eclat_true & 
                    work.Int.sub(\$14724_binop_int6435902_arg\(80 to 95), X"000" & X"1") & \$14724_binop_int6435902_arg\(96 to 151) & \$14724_binop_int6435902_arg\(152 to 153);
                    result6468 := \$14724_binop_int6435902_result\;
                    rdy6469 := eclat_true;
                    state_var7460 := IDLE6470;
                  else
                    \$14773_modulo6685896_id\ := "000001010000";
                    \$14773_modulo6685896_arg\ := work.Int.absv(\$14724_binop_int6435902_arg\(48 to 78)) & 
                    work.Int.absv(\$14738_v\(0 to 30));
                    state_var7460 := \$14773_MODULO6685896\;
                  end if;
                when X"0000000" & X"5" =>
                  \$14742_res\ := work.Int.land(\$14724_binop_int6435902_arg\(48 to 78), \$14738_v\(0 to 30));
                  \$14724_binop_int6435902_result\ := work.Int.add(\$14724_binop_int6435902_arg\(32 to 47), X"000" & X"1") & \$14742_res\ & eclat_true & 
                  work.Int.sub(\$14724_binop_int6435902_arg\(80 to 95), X"000" & X"1") & \$14724_binop_int6435902_arg\(96 to 151) & \$14724_binop_int6435902_arg\(152 to 153);
                  result6468 := \$14724_binop_int6435902_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"6" =>
                  \$14742_res\ := work.Int.lor(\$14724_binop_int6435902_arg\(48 to 78), \$14738_v\(0 to 30));
                  \$14724_binop_int6435902_result\ := work.Int.add(\$14724_binop_int6435902_arg\(32 to 47), X"000" & X"1") & \$14742_res\ & eclat_true & 
                  work.Int.sub(\$14724_binop_int6435902_arg\(80 to 95), X"000" & X"1") & \$14724_binop_int6435902_arg\(96 to 151) & \$14724_binop_int6435902_arg\(152 to 153);
                  result6468 := \$14724_binop_int6435902_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"7" =>
                  \$14742_res\ := work.Int.lxor(\$14724_binop_int6435902_arg\(48 to 78), \$14738_v\(0 to 30));
                  \$14724_binop_int6435902_result\ := work.Int.add(\$14724_binop_int6435902_arg\(32 to 47), X"000" & X"1") & \$14742_res\ & eclat_true & 
                  work.Int.sub(\$14724_binop_int6435902_arg\(80 to 95), X"000" & X"1") & \$14724_binop_int6435902_arg\(96 to 151) & \$14724_binop_int6435902_arg\(152 to 153);
                  result6468 := \$14724_binop_int6435902_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"8" =>
                  \$14742_res\ := work.Int.lsl(\$14724_binop_int6435902_arg\(48 to 78), \$14738_v\(0 to 30));
                  \$14724_binop_int6435902_result\ := work.Int.add(\$14724_binop_int6435902_arg\(32 to 47), X"000" & X"1") & \$14742_res\ & eclat_true & 
                  work.Int.sub(\$14724_binop_int6435902_arg\(80 to 95), X"000" & X"1") & \$14724_binop_int6435902_arg\(96 to 151) & \$14724_binop_int6435902_arg\(152 to 153);
                  result6468 := \$14724_binop_int6435902_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"9" =>
                  \$14742_res\ := work.Int.lsr(\$14724_binop_int6435902_arg\(48 to 78), \$14738_v\(0 to 30));
                  \$14724_binop_int6435902_result\ := work.Int.add(\$14724_binop_int6435902_arg\(32 to 47), X"000" & X"1") & \$14742_res\ & eclat_true & 
                  work.Int.sub(\$14724_binop_int6435902_arg\(80 to 95), X"000" & X"1") & \$14724_binop_int6435902_arg\(96 to 151) & \$14724_binop_int6435902_arg\(152 to 153);
                  result6468 := \$14724_binop_int6435902_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"a" =>
                  \$14742_res\ := work.Int.asr(\$14724_binop_int6435902_arg\(48 to 78), \$14738_v\(0 to 30));
                  \$14724_binop_int6435902_result\ := work.Int.add(\$14724_binop_int6435902_arg\(32 to 47), X"000" & X"1") & \$14742_res\ & eclat_true & 
                  work.Int.sub(\$14724_binop_int6435902_arg\(80 to 95), X"000" & X"1") & \$14724_binop_int6435902_arg\(96 to 151) & \$14724_binop_int6435902_arg\(152 to 153);
                  result6468 := \$14724_binop_int6435902_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"b" =>
                  \$14742_res\ := eclat_if(work.Int.lt(\$14724_binop_int6435902_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$14738_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.gt(\$14724_binop_int6435902_arg\(48 to 78), \$14738_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$14738_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"0" & 
                                  eclat_if(work.Int.lt(\$14724_binop_int6435902_arg\(48 to 78), \$14738_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$14724_binop_int6435902_result\ := work.Int.add(\$14724_binop_int6435902_arg\(32 to 47), X"000" & X"1") & \$14742_res\ & eclat_true & 
                  work.Int.sub(\$14724_binop_int6435902_arg\(80 to 95), X"000" & X"1") & \$14724_binop_int6435902_arg\(96 to 151) & \$14724_binop_int6435902_arg\(152 to 153);
                  result6468 := \$14724_binop_int6435902_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"c" =>
                  \$14742_res\ := eclat_if(work.Int.lt(\$14724_binop_int6435902_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$14738_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.le(\$14724_binop_int6435902_arg\(48 to 78), \$14738_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"1") & 
                                  eclat_if(work.Int.lt(\$14738_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & 
                                  eclat_if(work.Int.ge(\$14724_binop_int6435902_arg\(48 to 78), \$14738_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$14724_binop_int6435902_result\ := work.Int.add(\$14724_binop_int6435902_arg\(32 to 47), X"000" & X"1") & \$14742_res\ & eclat_true & 
                  work.Int.sub(\$14724_binop_int6435902_arg\(80 to 95), X"000" & X"1") & \$14724_binop_int6435902_arg\(96 to 151) & \$14724_binop_int6435902_arg\(152 to 153);
                  result6468 := \$14724_binop_int6435902_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when others =>
                  \$14742_res\ := "000"& X"000000" & X"0";
                  \$14724_binop_int6435902_result\ := work.Int.add(\$14724_binop_int6435902_arg\(32 to 47), X"000" & X"1") & \$14742_res\ & eclat_true & 
                  work.Int.sub(\$14724_binop_int6435902_arg\(80 to 95), X"000" & X"1") & \$14724_binop_int6435902_arg\(96 to 151) & \$14724_binop_int6435902_arg\(152 to 153);
                  result6468 := \$14724_binop_int6435902_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                end case;
              when PAUSE_GET7048 =>
                \$14818_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7047\ := \$14804_binop_int6435903_arg\(0 to 31);
                case \$v7047\ is
                when X"0000000" & X"0" =>
                  \$14822_res\ := work.Int.add(\$14804_binop_int6435903_arg\(48 to 78), \$14818_v\(0 to 30));
                  \$14804_binop_int6435903_result\ := work.Int.add(\$14804_binop_int6435903_arg\(32 to 47), X"000" & X"1") & \$14822_res\ & eclat_true & 
                  work.Int.sub(\$14804_binop_int6435903_arg\(80 to 95), X"000" & X"1") & \$14804_binop_int6435903_arg\(96 to 151) & \$14804_binop_int6435903_arg\(152 to 153);
                  result6468 := \$14804_binop_int6435903_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"1" =>
                  \$14822_res\ := work.Int.sub(\$14804_binop_int6435903_arg\(48 to 78), \$14818_v\(0 to 30));
                  \$14804_binop_int6435903_result\ := work.Int.add(\$14804_binop_int6435903_arg\(32 to 47), X"000" & X"1") & \$14822_res\ & eclat_true & 
                  work.Int.sub(\$14804_binop_int6435903_arg\(80 to 95), X"000" & X"1") & \$14804_binop_int6435903_arg\(96 to 151) & \$14804_binop_int6435903_arg\(152 to 153);
                  result6468 := \$14804_binop_int6435903_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"2" =>
                  \$14822_res\ := work.Int.mul(\$14804_binop_int6435903_arg\(48 to 78), \$14818_v\(0 to 30));
                  \$14804_binop_int6435903_result\ := work.Int.add(\$14804_binop_int6435903_arg\(32 to 47), X"000" & X"1") & \$14822_res\ & eclat_true & 
                  work.Int.sub(\$14804_binop_int6435903_arg\(80 to 95), X"000" & X"1") & \$14804_binop_int6435903_arg\(96 to 151) & \$14804_binop_int6435903_arg\(152 to 153);
                  result6468 := \$14804_binop_int6435903_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"3" =>
                  \$v7043\ := work.Int.eq(\$14818_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v7043\(0) = '1' then
                    \$14822_res\ := "000"& X"000000" & X"0";
                    \$14804_binop_int6435903_result\ := work.Int.add(
                                                        \$14804_binop_int6435903_arg\(32 to 47), X"000" & X"1") & \$14822_res\ & eclat_true & 
                    work.Int.sub(\$14804_binop_int6435903_arg\(80 to 95), X"000" & X"1") & \$14804_binop_int6435903_arg\(96 to 151) & \$14804_binop_int6435903_arg\(152 to 153);
                    result6468 := \$14804_binop_int6435903_result\;
                    rdy6469 := eclat_true;
                    state_var7460 := IDLE6470;
                  else
                    \$14829_modulo6685895_id\ := "000001010011";
                    \$14829_modulo6685895_arg\ := work.Int.absv(\$14804_binop_int6435903_arg\(48 to 78)) & 
                    work.Int.absv(\$14818_v\(0 to 30));
                    state_var7460 := \$14829_MODULO6685895\;
                  end if;
                when X"0000000" & X"4" =>
                  \$v7046\ := work.Int.eq(\$14818_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v7046\(0) = '1' then
                    \$14822_res\ := "000"& X"000000" & X"0";
                    \$14804_binop_int6435903_result\ := work.Int.add(
                                                        \$14804_binop_int6435903_arg\(32 to 47), X"000" & X"1") & \$14822_res\ & eclat_true & 
                    work.Int.sub(\$14804_binop_int6435903_arg\(80 to 95), X"000" & X"1") & \$14804_binop_int6435903_arg\(96 to 151) & \$14804_binop_int6435903_arg\(152 to 153);
                    result6468 := \$14804_binop_int6435903_result\;
                    rdy6469 := eclat_true;
                    state_var7460 := IDLE6470;
                  else
                    \$14853_modulo6685896_id\ := "000001010101";
                    \$14853_modulo6685896_arg\ := work.Int.absv(\$14804_binop_int6435903_arg\(48 to 78)) & 
                    work.Int.absv(\$14818_v\(0 to 30));
                    state_var7460 := \$14853_MODULO6685896\;
                  end if;
                when X"0000000" & X"5" =>
                  \$14822_res\ := work.Int.land(\$14804_binop_int6435903_arg\(48 to 78), \$14818_v\(0 to 30));
                  \$14804_binop_int6435903_result\ := work.Int.add(\$14804_binop_int6435903_arg\(32 to 47), X"000" & X"1") & \$14822_res\ & eclat_true & 
                  work.Int.sub(\$14804_binop_int6435903_arg\(80 to 95), X"000" & X"1") & \$14804_binop_int6435903_arg\(96 to 151) & \$14804_binop_int6435903_arg\(152 to 153);
                  result6468 := \$14804_binop_int6435903_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"6" =>
                  \$14822_res\ := work.Int.lor(\$14804_binop_int6435903_arg\(48 to 78), \$14818_v\(0 to 30));
                  \$14804_binop_int6435903_result\ := work.Int.add(\$14804_binop_int6435903_arg\(32 to 47), X"000" & X"1") & \$14822_res\ & eclat_true & 
                  work.Int.sub(\$14804_binop_int6435903_arg\(80 to 95), X"000" & X"1") & \$14804_binop_int6435903_arg\(96 to 151) & \$14804_binop_int6435903_arg\(152 to 153);
                  result6468 := \$14804_binop_int6435903_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"7" =>
                  \$14822_res\ := work.Int.lxor(\$14804_binop_int6435903_arg\(48 to 78), \$14818_v\(0 to 30));
                  \$14804_binop_int6435903_result\ := work.Int.add(\$14804_binop_int6435903_arg\(32 to 47), X"000" & X"1") & \$14822_res\ & eclat_true & 
                  work.Int.sub(\$14804_binop_int6435903_arg\(80 to 95), X"000" & X"1") & \$14804_binop_int6435903_arg\(96 to 151) & \$14804_binop_int6435903_arg\(152 to 153);
                  result6468 := \$14804_binop_int6435903_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"8" =>
                  \$14822_res\ := work.Int.lsl(\$14804_binop_int6435903_arg\(48 to 78), \$14818_v\(0 to 30));
                  \$14804_binop_int6435903_result\ := work.Int.add(\$14804_binop_int6435903_arg\(32 to 47), X"000" & X"1") & \$14822_res\ & eclat_true & 
                  work.Int.sub(\$14804_binop_int6435903_arg\(80 to 95), X"000" & X"1") & \$14804_binop_int6435903_arg\(96 to 151) & \$14804_binop_int6435903_arg\(152 to 153);
                  result6468 := \$14804_binop_int6435903_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"9" =>
                  \$14822_res\ := work.Int.lsr(\$14804_binop_int6435903_arg\(48 to 78), \$14818_v\(0 to 30));
                  \$14804_binop_int6435903_result\ := work.Int.add(\$14804_binop_int6435903_arg\(32 to 47), X"000" & X"1") & \$14822_res\ & eclat_true & 
                  work.Int.sub(\$14804_binop_int6435903_arg\(80 to 95), X"000" & X"1") & \$14804_binop_int6435903_arg\(96 to 151) & \$14804_binop_int6435903_arg\(152 to 153);
                  result6468 := \$14804_binop_int6435903_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"a" =>
                  \$14822_res\ := work.Int.asr(\$14804_binop_int6435903_arg\(48 to 78), \$14818_v\(0 to 30));
                  \$14804_binop_int6435903_result\ := work.Int.add(\$14804_binop_int6435903_arg\(32 to 47), X"000" & X"1") & \$14822_res\ & eclat_true & 
                  work.Int.sub(\$14804_binop_int6435903_arg\(80 to 95), X"000" & X"1") & \$14804_binop_int6435903_arg\(96 to 151) & \$14804_binop_int6435903_arg\(152 to 153);
                  result6468 := \$14804_binop_int6435903_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"b" =>
                  \$14822_res\ := eclat_if(work.Int.lt(\$14804_binop_int6435903_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$14818_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.gt(\$14804_binop_int6435903_arg\(48 to 78), \$14818_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$14818_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"0" & 
                                  eclat_if(work.Int.lt(\$14804_binop_int6435903_arg\(48 to 78), \$14818_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$14804_binop_int6435903_result\ := work.Int.add(\$14804_binop_int6435903_arg\(32 to 47), X"000" & X"1") & \$14822_res\ & eclat_true & 
                  work.Int.sub(\$14804_binop_int6435903_arg\(80 to 95), X"000" & X"1") & \$14804_binop_int6435903_arg\(96 to 151) & \$14804_binop_int6435903_arg\(152 to 153);
                  result6468 := \$14804_binop_int6435903_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"c" =>
                  \$14822_res\ := eclat_if(work.Int.lt(\$14804_binop_int6435903_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$14818_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.le(\$14804_binop_int6435903_arg\(48 to 78), \$14818_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"1") & 
                                  eclat_if(work.Int.lt(\$14818_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & 
                                  eclat_if(work.Int.ge(\$14804_binop_int6435903_arg\(48 to 78), \$14818_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$14804_binop_int6435903_result\ := work.Int.add(\$14804_binop_int6435903_arg\(32 to 47), X"000" & X"1") & \$14822_res\ & eclat_true & 
                  work.Int.sub(\$14804_binop_int6435903_arg\(80 to 95), X"000" & X"1") & \$14804_binop_int6435903_arg\(96 to 151) & \$14804_binop_int6435903_arg\(152 to 153);
                  result6468 := \$14804_binop_int6435903_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when others =>
                  \$14822_res\ := "000"& X"000000" & X"0";
                  \$14804_binop_int6435903_result\ := work.Int.add(\$14804_binop_int6435903_arg\(32 to 47), X"000" & X"1") & \$14822_res\ & eclat_true & 
                  work.Int.sub(\$14804_binop_int6435903_arg\(80 to 95), X"000" & X"1") & \$14804_binop_int6435903_arg\(96 to 151) & \$14804_binop_int6435903_arg\(152 to 153);
                  result6468 := \$14804_binop_int6435903_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                end case;
              when PAUSE_GET7058 =>
                \$14898_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7057\ := \$14884_binop_int6435904_arg\(0 to 31);
                case \$v7057\ is
                when X"0000000" & X"0" =>
                  \$14902_res\ := work.Int.add(\$14884_binop_int6435904_arg\(48 to 78), \$14898_v\(0 to 30));
                  \$14884_binop_int6435904_result\ := work.Int.add(\$14884_binop_int6435904_arg\(32 to 47), X"000" & X"1") & \$14902_res\ & eclat_true & 
                  work.Int.sub(\$14884_binop_int6435904_arg\(80 to 95), X"000" & X"1") & \$14884_binop_int6435904_arg\(96 to 151) & \$14884_binop_int6435904_arg\(152 to 153);
                  result6468 := \$14884_binop_int6435904_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"1" =>
                  \$14902_res\ := work.Int.sub(\$14884_binop_int6435904_arg\(48 to 78), \$14898_v\(0 to 30));
                  \$14884_binop_int6435904_result\ := work.Int.add(\$14884_binop_int6435904_arg\(32 to 47), X"000" & X"1") & \$14902_res\ & eclat_true & 
                  work.Int.sub(\$14884_binop_int6435904_arg\(80 to 95), X"000" & X"1") & \$14884_binop_int6435904_arg\(96 to 151) & \$14884_binop_int6435904_arg\(152 to 153);
                  result6468 := \$14884_binop_int6435904_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"2" =>
                  \$14902_res\ := work.Int.mul(\$14884_binop_int6435904_arg\(48 to 78), \$14898_v\(0 to 30));
                  \$14884_binop_int6435904_result\ := work.Int.add(\$14884_binop_int6435904_arg\(32 to 47), X"000" & X"1") & \$14902_res\ & eclat_true & 
                  work.Int.sub(\$14884_binop_int6435904_arg\(80 to 95), X"000" & X"1") & \$14884_binop_int6435904_arg\(96 to 151) & \$14884_binop_int6435904_arg\(152 to 153);
                  result6468 := \$14884_binop_int6435904_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"3" =>
                  \$v7053\ := work.Int.eq(\$14898_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v7053\(0) = '1' then
                    \$14902_res\ := "000"& X"000000" & X"0";
                    \$14884_binop_int6435904_result\ := work.Int.add(
                                                        \$14884_binop_int6435904_arg\(32 to 47), X"000" & X"1") & \$14902_res\ & eclat_true & 
                    work.Int.sub(\$14884_binop_int6435904_arg\(80 to 95), X"000" & X"1") & \$14884_binop_int6435904_arg\(96 to 151) & \$14884_binop_int6435904_arg\(152 to 153);
                    result6468 := \$14884_binop_int6435904_result\;
                    rdy6469 := eclat_true;
                    state_var7460 := IDLE6470;
                  else
                    \$14909_modulo6685895_id\ := "000001011000";
                    \$14909_modulo6685895_arg\ := work.Int.absv(\$14884_binop_int6435904_arg\(48 to 78)) & 
                    work.Int.absv(\$14898_v\(0 to 30));
                    state_var7460 := \$14909_MODULO6685895\;
                  end if;
                when X"0000000" & X"4" =>
                  \$v7056\ := work.Int.eq(\$14898_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v7056\(0) = '1' then
                    \$14902_res\ := "000"& X"000000" & X"0";
                    \$14884_binop_int6435904_result\ := work.Int.add(
                                                        \$14884_binop_int6435904_arg\(32 to 47), X"000" & X"1") & \$14902_res\ & eclat_true & 
                    work.Int.sub(\$14884_binop_int6435904_arg\(80 to 95), X"000" & X"1") & \$14884_binop_int6435904_arg\(96 to 151) & \$14884_binop_int6435904_arg\(152 to 153);
                    result6468 := \$14884_binop_int6435904_result\;
                    rdy6469 := eclat_true;
                    state_var7460 := IDLE6470;
                  else
                    \$14933_modulo6685896_id\ := "000001011010";
                    \$14933_modulo6685896_arg\ := work.Int.absv(\$14884_binop_int6435904_arg\(48 to 78)) & 
                    work.Int.absv(\$14898_v\(0 to 30));
                    state_var7460 := \$14933_MODULO6685896\;
                  end if;
                when X"0000000" & X"5" =>
                  \$14902_res\ := work.Int.land(\$14884_binop_int6435904_arg\(48 to 78), \$14898_v\(0 to 30));
                  \$14884_binop_int6435904_result\ := work.Int.add(\$14884_binop_int6435904_arg\(32 to 47), X"000" & X"1") & \$14902_res\ & eclat_true & 
                  work.Int.sub(\$14884_binop_int6435904_arg\(80 to 95), X"000" & X"1") & \$14884_binop_int6435904_arg\(96 to 151) & \$14884_binop_int6435904_arg\(152 to 153);
                  result6468 := \$14884_binop_int6435904_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"6" =>
                  \$14902_res\ := work.Int.lor(\$14884_binop_int6435904_arg\(48 to 78), \$14898_v\(0 to 30));
                  \$14884_binop_int6435904_result\ := work.Int.add(\$14884_binop_int6435904_arg\(32 to 47), X"000" & X"1") & \$14902_res\ & eclat_true & 
                  work.Int.sub(\$14884_binop_int6435904_arg\(80 to 95), X"000" & X"1") & \$14884_binop_int6435904_arg\(96 to 151) & \$14884_binop_int6435904_arg\(152 to 153);
                  result6468 := \$14884_binop_int6435904_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"7" =>
                  \$14902_res\ := work.Int.lxor(\$14884_binop_int6435904_arg\(48 to 78), \$14898_v\(0 to 30));
                  \$14884_binop_int6435904_result\ := work.Int.add(\$14884_binop_int6435904_arg\(32 to 47), X"000" & X"1") & \$14902_res\ & eclat_true & 
                  work.Int.sub(\$14884_binop_int6435904_arg\(80 to 95), X"000" & X"1") & \$14884_binop_int6435904_arg\(96 to 151) & \$14884_binop_int6435904_arg\(152 to 153);
                  result6468 := \$14884_binop_int6435904_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"8" =>
                  \$14902_res\ := work.Int.lsl(\$14884_binop_int6435904_arg\(48 to 78), \$14898_v\(0 to 30));
                  \$14884_binop_int6435904_result\ := work.Int.add(\$14884_binop_int6435904_arg\(32 to 47), X"000" & X"1") & \$14902_res\ & eclat_true & 
                  work.Int.sub(\$14884_binop_int6435904_arg\(80 to 95), X"000" & X"1") & \$14884_binop_int6435904_arg\(96 to 151) & \$14884_binop_int6435904_arg\(152 to 153);
                  result6468 := \$14884_binop_int6435904_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"9" =>
                  \$14902_res\ := work.Int.lsr(\$14884_binop_int6435904_arg\(48 to 78), \$14898_v\(0 to 30));
                  \$14884_binop_int6435904_result\ := work.Int.add(\$14884_binop_int6435904_arg\(32 to 47), X"000" & X"1") & \$14902_res\ & eclat_true & 
                  work.Int.sub(\$14884_binop_int6435904_arg\(80 to 95), X"000" & X"1") & \$14884_binop_int6435904_arg\(96 to 151) & \$14884_binop_int6435904_arg\(152 to 153);
                  result6468 := \$14884_binop_int6435904_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"a" =>
                  \$14902_res\ := work.Int.asr(\$14884_binop_int6435904_arg\(48 to 78), \$14898_v\(0 to 30));
                  \$14884_binop_int6435904_result\ := work.Int.add(\$14884_binop_int6435904_arg\(32 to 47), X"000" & X"1") & \$14902_res\ & eclat_true & 
                  work.Int.sub(\$14884_binop_int6435904_arg\(80 to 95), X"000" & X"1") & \$14884_binop_int6435904_arg\(96 to 151) & \$14884_binop_int6435904_arg\(152 to 153);
                  result6468 := \$14884_binop_int6435904_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"b" =>
                  \$14902_res\ := eclat_if(work.Int.lt(\$14884_binop_int6435904_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$14898_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.gt(\$14884_binop_int6435904_arg\(48 to 78), \$14898_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$14898_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"0" & 
                                  eclat_if(work.Int.lt(\$14884_binop_int6435904_arg\(48 to 78), \$14898_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$14884_binop_int6435904_result\ := work.Int.add(\$14884_binop_int6435904_arg\(32 to 47), X"000" & X"1") & \$14902_res\ & eclat_true & 
                  work.Int.sub(\$14884_binop_int6435904_arg\(80 to 95), X"000" & X"1") & \$14884_binop_int6435904_arg\(96 to 151) & \$14884_binop_int6435904_arg\(152 to 153);
                  result6468 := \$14884_binop_int6435904_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"c" =>
                  \$14902_res\ := eclat_if(work.Int.lt(\$14884_binop_int6435904_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$14898_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.le(\$14884_binop_int6435904_arg\(48 to 78), \$14898_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"1") & 
                                  eclat_if(work.Int.lt(\$14898_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & 
                                  eclat_if(work.Int.ge(\$14884_binop_int6435904_arg\(48 to 78), \$14898_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$14884_binop_int6435904_result\ := work.Int.add(\$14884_binop_int6435904_arg\(32 to 47), X"000" & X"1") & \$14902_res\ & eclat_true & 
                  work.Int.sub(\$14884_binop_int6435904_arg\(80 to 95), X"000" & X"1") & \$14884_binop_int6435904_arg\(96 to 151) & \$14884_binop_int6435904_arg\(152 to 153);
                  result6468 := \$14884_binop_int6435904_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when others =>
                  \$14902_res\ := "000"& X"000000" & X"0";
                  \$14884_binop_int6435904_result\ := work.Int.add(\$14884_binop_int6435904_arg\(32 to 47), X"000" & X"1") & \$14902_res\ & eclat_true & 
                  work.Int.sub(\$14884_binop_int6435904_arg\(80 to 95), X"000" & X"1") & \$14884_binop_int6435904_arg\(96 to 151) & \$14884_binop_int6435904_arg\(152 to 153);
                  result6468 := \$14884_binop_int6435904_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                end case;
              when PAUSE_GET7068 =>
                \$14978_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7067\ := \$14964_binop_int6435905_arg\(0 to 31);
                case \$v7067\ is
                when X"0000000" & X"0" =>
                  \$14982_res\ := work.Int.add(\$14964_binop_int6435905_arg\(48 to 78), \$14978_v\(0 to 30));
                  \$14964_binop_int6435905_result\ := work.Int.add(\$14964_binop_int6435905_arg\(32 to 47), X"000" & X"1") & \$14982_res\ & eclat_true & 
                  work.Int.sub(\$14964_binop_int6435905_arg\(80 to 95), X"000" & X"1") & \$14964_binop_int6435905_arg\(96 to 151) & \$14964_binop_int6435905_arg\(152 to 153);
                  result6468 := \$14964_binop_int6435905_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"1" =>
                  \$14982_res\ := work.Int.sub(\$14964_binop_int6435905_arg\(48 to 78), \$14978_v\(0 to 30));
                  \$14964_binop_int6435905_result\ := work.Int.add(\$14964_binop_int6435905_arg\(32 to 47), X"000" & X"1") & \$14982_res\ & eclat_true & 
                  work.Int.sub(\$14964_binop_int6435905_arg\(80 to 95), X"000" & X"1") & \$14964_binop_int6435905_arg\(96 to 151) & \$14964_binop_int6435905_arg\(152 to 153);
                  result6468 := \$14964_binop_int6435905_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"2" =>
                  \$14982_res\ := work.Int.mul(\$14964_binop_int6435905_arg\(48 to 78), \$14978_v\(0 to 30));
                  \$14964_binop_int6435905_result\ := work.Int.add(\$14964_binop_int6435905_arg\(32 to 47), X"000" & X"1") & \$14982_res\ & eclat_true & 
                  work.Int.sub(\$14964_binop_int6435905_arg\(80 to 95), X"000" & X"1") & \$14964_binop_int6435905_arg\(96 to 151) & \$14964_binop_int6435905_arg\(152 to 153);
                  result6468 := \$14964_binop_int6435905_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"3" =>
                  \$v7063\ := work.Int.eq(\$14978_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v7063\(0) = '1' then
                    \$14982_res\ := "000"& X"000000" & X"0";
                    \$14964_binop_int6435905_result\ := work.Int.add(
                                                        \$14964_binop_int6435905_arg\(32 to 47), X"000" & X"1") & \$14982_res\ & eclat_true & 
                    work.Int.sub(\$14964_binop_int6435905_arg\(80 to 95), X"000" & X"1") & \$14964_binop_int6435905_arg\(96 to 151) & \$14964_binop_int6435905_arg\(152 to 153);
                    result6468 := \$14964_binop_int6435905_result\;
                    rdy6469 := eclat_true;
                    state_var7460 := IDLE6470;
                  else
                    \$14989_modulo6685895_id\ := "000001011101";
                    \$14989_modulo6685895_arg\ := work.Int.absv(\$14964_binop_int6435905_arg\(48 to 78)) & 
                    work.Int.absv(\$14978_v\(0 to 30));
                    state_var7460 := \$14989_MODULO6685895\;
                  end if;
                when X"0000000" & X"4" =>
                  \$v7066\ := work.Int.eq(\$14978_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v7066\(0) = '1' then
                    \$14982_res\ := "000"& X"000000" & X"0";
                    \$14964_binop_int6435905_result\ := work.Int.add(
                                                        \$14964_binop_int6435905_arg\(32 to 47), X"000" & X"1") & \$14982_res\ & eclat_true & 
                    work.Int.sub(\$14964_binop_int6435905_arg\(80 to 95), X"000" & X"1") & \$14964_binop_int6435905_arg\(96 to 151) & \$14964_binop_int6435905_arg\(152 to 153);
                    result6468 := \$14964_binop_int6435905_result\;
                    rdy6469 := eclat_true;
                    state_var7460 := IDLE6470;
                  else
                    \$15013_modulo6685896_id\ := "000001011111";
                    \$15013_modulo6685896_arg\ := work.Int.absv(\$14964_binop_int6435905_arg\(48 to 78)) & 
                    work.Int.absv(\$14978_v\(0 to 30));
                    state_var7460 := \$15013_MODULO6685896\;
                  end if;
                when X"0000000" & X"5" =>
                  \$14982_res\ := work.Int.land(\$14964_binop_int6435905_arg\(48 to 78), \$14978_v\(0 to 30));
                  \$14964_binop_int6435905_result\ := work.Int.add(\$14964_binop_int6435905_arg\(32 to 47), X"000" & X"1") & \$14982_res\ & eclat_true & 
                  work.Int.sub(\$14964_binop_int6435905_arg\(80 to 95), X"000" & X"1") & \$14964_binop_int6435905_arg\(96 to 151) & \$14964_binop_int6435905_arg\(152 to 153);
                  result6468 := \$14964_binop_int6435905_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"6" =>
                  \$14982_res\ := work.Int.lor(\$14964_binop_int6435905_arg\(48 to 78), \$14978_v\(0 to 30));
                  \$14964_binop_int6435905_result\ := work.Int.add(\$14964_binop_int6435905_arg\(32 to 47), X"000" & X"1") & \$14982_res\ & eclat_true & 
                  work.Int.sub(\$14964_binop_int6435905_arg\(80 to 95), X"000" & X"1") & \$14964_binop_int6435905_arg\(96 to 151) & \$14964_binop_int6435905_arg\(152 to 153);
                  result6468 := \$14964_binop_int6435905_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"7" =>
                  \$14982_res\ := work.Int.lxor(\$14964_binop_int6435905_arg\(48 to 78), \$14978_v\(0 to 30));
                  \$14964_binop_int6435905_result\ := work.Int.add(\$14964_binop_int6435905_arg\(32 to 47), X"000" & X"1") & \$14982_res\ & eclat_true & 
                  work.Int.sub(\$14964_binop_int6435905_arg\(80 to 95), X"000" & X"1") & \$14964_binop_int6435905_arg\(96 to 151) & \$14964_binop_int6435905_arg\(152 to 153);
                  result6468 := \$14964_binop_int6435905_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"8" =>
                  \$14982_res\ := work.Int.lsl(\$14964_binop_int6435905_arg\(48 to 78), \$14978_v\(0 to 30));
                  \$14964_binop_int6435905_result\ := work.Int.add(\$14964_binop_int6435905_arg\(32 to 47), X"000" & X"1") & \$14982_res\ & eclat_true & 
                  work.Int.sub(\$14964_binop_int6435905_arg\(80 to 95), X"000" & X"1") & \$14964_binop_int6435905_arg\(96 to 151) & \$14964_binop_int6435905_arg\(152 to 153);
                  result6468 := \$14964_binop_int6435905_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"9" =>
                  \$14982_res\ := work.Int.lsr(\$14964_binop_int6435905_arg\(48 to 78), \$14978_v\(0 to 30));
                  \$14964_binop_int6435905_result\ := work.Int.add(\$14964_binop_int6435905_arg\(32 to 47), X"000" & X"1") & \$14982_res\ & eclat_true & 
                  work.Int.sub(\$14964_binop_int6435905_arg\(80 to 95), X"000" & X"1") & \$14964_binop_int6435905_arg\(96 to 151) & \$14964_binop_int6435905_arg\(152 to 153);
                  result6468 := \$14964_binop_int6435905_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"a" =>
                  \$14982_res\ := work.Int.asr(\$14964_binop_int6435905_arg\(48 to 78), \$14978_v\(0 to 30));
                  \$14964_binop_int6435905_result\ := work.Int.add(\$14964_binop_int6435905_arg\(32 to 47), X"000" & X"1") & \$14982_res\ & eclat_true & 
                  work.Int.sub(\$14964_binop_int6435905_arg\(80 to 95), X"000" & X"1") & \$14964_binop_int6435905_arg\(96 to 151) & \$14964_binop_int6435905_arg\(152 to 153);
                  result6468 := \$14964_binop_int6435905_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"b" =>
                  \$14982_res\ := eclat_if(work.Int.lt(\$14964_binop_int6435905_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$14978_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.gt(\$14964_binop_int6435905_arg\(48 to 78), \$14978_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$14978_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"0" & 
                                  eclat_if(work.Int.lt(\$14964_binop_int6435905_arg\(48 to 78), \$14978_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$14964_binop_int6435905_result\ := work.Int.add(\$14964_binop_int6435905_arg\(32 to 47), X"000" & X"1") & \$14982_res\ & eclat_true & 
                  work.Int.sub(\$14964_binop_int6435905_arg\(80 to 95), X"000" & X"1") & \$14964_binop_int6435905_arg\(96 to 151) & \$14964_binop_int6435905_arg\(152 to 153);
                  result6468 := \$14964_binop_int6435905_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"c" =>
                  \$14982_res\ := eclat_if(work.Int.lt(\$14964_binop_int6435905_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$14978_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.le(\$14964_binop_int6435905_arg\(48 to 78), \$14978_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"1") & 
                                  eclat_if(work.Int.lt(\$14978_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & 
                                  eclat_if(work.Int.ge(\$14964_binop_int6435905_arg\(48 to 78), \$14978_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$14964_binop_int6435905_result\ := work.Int.add(\$14964_binop_int6435905_arg\(32 to 47), X"000" & X"1") & \$14982_res\ & eclat_true & 
                  work.Int.sub(\$14964_binop_int6435905_arg\(80 to 95), X"000" & X"1") & \$14964_binop_int6435905_arg\(96 to 151) & \$14964_binop_int6435905_arg\(152 to 153);
                  result6468 := \$14964_binop_int6435905_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when others =>
                  \$14982_res\ := "000"& X"000000" & X"0";
                  \$14964_binop_int6435905_result\ := work.Int.add(\$14964_binop_int6435905_arg\(32 to 47), X"000" & X"1") & \$14982_res\ & eclat_true & 
                  work.Int.sub(\$14964_binop_int6435905_arg\(80 to 95), X"000" & X"1") & \$14964_binop_int6435905_arg\(96 to 151) & \$14964_binop_int6435905_arg\(152 to 153);
                  result6468 := \$14964_binop_int6435905_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                end case;
              when PAUSE_GET7078 =>
                \$15058_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7077\ := \$15044_binop_int6435906_arg\(0 to 31);
                case \$v7077\ is
                when X"0000000" & X"0" =>
                  \$15062_res\ := work.Int.add(\$15044_binop_int6435906_arg\(48 to 78), \$15058_v\(0 to 30));
                  \$15044_binop_int6435906_result\ := work.Int.add(\$15044_binop_int6435906_arg\(32 to 47), X"000" & X"1") & \$15062_res\ & eclat_true & 
                  work.Int.sub(\$15044_binop_int6435906_arg\(80 to 95), X"000" & X"1") & \$15044_binop_int6435906_arg\(96 to 151) & \$15044_binop_int6435906_arg\(152 to 153);
                  result6468 := \$15044_binop_int6435906_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"1" =>
                  \$15062_res\ := work.Int.sub(\$15044_binop_int6435906_arg\(48 to 78), \$15058_v\(0 to 30));
                  \$15044_binop_int6435906_result\ := work.Int.add(\$15044_binop_int6435906_arg\(32 to 47), X"000" & X"1") & \$15062_res\ & eclat_true & 
                  work.Int.sub(\$15044_binop_int6435906_arg\(80 to 95), X"000" & X"1") & \$15044_binop_int6435906_arg\(96 to 151) & \$15044_binop_int6435906_arg\(152 to 153);
                  result6468 := \$15044_binop_int6435906_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"2" =>
                  \$15062_res\ := work.Int.mul(\$15044_binop_int6435906_arg\(48 to 78), \$15058_v\(0 to 30));
                  \$15044_binop_int6435906_result\ := work.Int.add(\$15044_binop_int6435906_arg\(32 to 47), X"000" & X"1") & \$15062_res\ & eclat_true & 
                  work.Int.sub(\$15044_binop_int6435906_arg\(80 to 95), X"000" & X"1") & \$15044_binop_int6435906_arg\(96 to 151) & \$15044_binop_int6435906_arg\(152 to 153);
                  result6468 := \$15044_binop_int6435906_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"3" =>
                  \$v7073\ := work.Int.eq(\$15058_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v7073\(0) = '1' then
                    \$15062_res\ := "000"& X"000000" & X"0";
                    \$15044_binop_int6435906_result\ := work.Int.add(
                                                        \$15044_binop_int6435906_arg\(32 to 47), X"000" & X"1") & \$15062_res\ & eclat_true & 
                    work.Int.sub(\$15044_binop_int6435906_arg\(80 to 95), X"000" & X"1") & \$15044_binop_int6435906_arg\(96 to 151) & \$15044_binop_int6435906_arg\(152 to 153);
                    result6468 := \$15044_binop_int6435906_result\;
                    rdy6469 := eclat_true;
                    state_var7460 := IDLE6470;
                  else
                    \$15069_modulo6685895_id\ := "000001100010";
                    \$15069_modulo6685895_arg\ := work.Int.absv(\$15044_binop_int6435906_arg\(48 to 78)) & 
                    work.Int.absv(\$15058_v\(0 to 30));
                    state_var7460 := \$15069_MODULO6685895\;
                  end if;
                when X"0000000" & X"4" =>
                  \$v7076\ := work.Int.eq(\$15058_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v7076\(0) = '1' then
                    \$15062_res\ := "000"& X"000000" & X"0";
                    \$15044_binop_int6435906_result\ := work.Int.add(
                                                        \$15044_binop_int6435906_arg\(32 to 47), X"000" & X"1") & \$15062_res\ & eclat_true & 
                    work.Int.sub(\$15044_binop_int6435906_arg\(80 to 95), X"000" & X"1") & \$15044_binop_int6435906_arg\(96 to 151) & \$15044_binop_int6435906_arg\(152 to 153);
                    result6468 := \$15044_binop_int6435906_result\;
                    rdy6469 := eclat_true;
                    state_var7460 := IDLE6470;
                  else
                    \$15093_modulo6685896_id\ := "000001100100";
                    \$15093_modulo6685896_arg\ := work.Int.absv(\$15044_binop_int6435906_arg\(48 to 78)) & 
                    work.Int.absv(\$15058_v\(0 to 30));
                    state_var7460 := \$15093_MODULO6685896\;
                  end if;
                when X"0000000" & X"5" =>
                  \$15062_res\ := work.Int.land(\$15044_binop_int6435906_arg\(48 to 78), \$15058_v\(0 to 30));
                  \$15044_binop_int6435906_result\ := work.Int.add(\$15044_binop_int6435906_arg\(32 to 47), X"000" & X"1") & \$15062_res\ & eclat_true & 
                  work.Int.sub(\$15044_binop_int6435906_arg\(80 to 95), X"000" & X"1") & \$15044_binop_int6435906_arg\(96 to 151) & \$15044_binop_int6435906_arg\(152 to 153);
                  result6468 := \$15044_binop_int6435906_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"6" =>
                  \$15062_res\ := work.Int.lor(\$15044_binop_int6435906_arg\(48 to 78), \$15058_v\(0 to 30));
                  \$15044_binop_int6435906_result\ := work.Int.add(\$15044_binop_int6435906_arg\(32 to 47), X"000" & X"1") & \$15062_res\ & eclat_true & 
                  work.Int.sub(\$15044_binop_int6435906_arg\(80 to 95), X"000" & X"1") & \$15044_binop_int6435906_arg\(96 to 151) & \$15044_binop_int6435906_arg\(152 to 153);
                  result6468 := \$15044_binop_int6435906_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"7" =>
                  \$15062_res\ := work.Int.lxor(\$15044_binop_int6435906_arg\(48 to 78), \$15058_v\(0 to 30));
                  \$15044_binop_int6435906_result\ := work.Int.add(\$15044_binop_int6435906_arg\(32 to 47), X"000" & X"1") & \$15062_res\ & eclat_true & 
                  work.Int.sub(\$15044_binop_int6435906_arg\(80 to 95), X"000" & X"1") & \$15044_binop_int6435906_arg\(96 to 151) & \$15044_binop_int6435906_arg\(152 to 153);
                  result6468 := \$15044_binop_int6435906_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"8" =>
                  \$15062_res\ := work.Int.lsl(\$15044_binop_int6435906_arg\(48 to 78), \$15058_v\(0 to 30));
                  \$15044_binop_int6435906_result\ := work.Int.add(\$15044_binop_int6435906_arg\(32 to 47), X"000" & X"1") & \$15062_res\ & eclat_true & 
                  work.Int.sub(\$15044_binop_int6435906_arg\(80 to 95), X"000" & X"1") & \$15044_binop_int6435906_arg\(96 to 151) & \$15044_binop_int6435906_arg\(152 to 153);
                  result6468 := \$15044_binop_int6435906_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"9" =>
                  \$15062_res\ := work.Int.lsr(\$15044_binop_int6435906_arg\(48 to 78), \$15058_v\(0 to 30));
                  \$15044_binop_int6435906_result\ := work.Int.add(\$15044_binop_int6435906_arg\(32 to 47), X"000" & X"1") & \$15062_res\ & eclat_true & 
                  work.Int.sub(\$15044_binop_int6435906_arg\(80 to 95), X"000" & X"1") & \$15044_binop_int6435906_arg\(96 to 151) & \$15044_binop_int6435906_arg\(152 to 153);
                  result6468 := \$15044_binop_int6435906_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"a" =>
                  \$15062_res\ := work.Int.asr(\$15044_binop_int6435906_arg\(48 to 78), \$15058_v\(0 to 30));
                  \$15044_binop_int6435906_result\ := work.Int.add(\$15044_binop_int6435906_arg\(32 to 47), X"000" & X"1") & \$15062_res\ & eclat_true & 
                  work.Int.sub(\$15044_binop_int6435906_arg\(80 to 95), X"000" & X"1") & \$15044_binop_int6435906_arg\(96 to 151) & \$15044_binop_int6435906_arg\(152 to 153);
                  result6468 := \$15044_binop_int6435906_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"b" =>
                  \$15062_res\ := eclat_if(work.Int.lt(\$15044_binop_int6435906_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$15058_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.gt(\$15044_binop_int6435906_arg\(48 to 78), \$15058_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$15058_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"0" & 
                                  eclat_if(work.Int.lt(\$15044_binop_int6435906_arg\(48 to 78), \$15058_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$15044_binop_int6435906_result\ := work.Int.add(\$15044_binop_int6435906_arg\(32 to 47), X"000" & X"1") & \$15062_res\ & eclat_true & 
                  work.Int.sub(\$15044_binop_int6435906_arg\(80 to 95), X"000" & X"1") & \$15044_binop_int6435906_arg\(96 to 151) & \$15044_binop_int6435906_arg\(152 to 153);
                  result6468 := \$15044_binop_int6435906_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"c" =>
                  \$15062_res\ := eclat_if(work.Int.lt(\$15044_binop_int6435906_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$15058_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.le(\$15044_binop_int6435906_arg\(48 to 78), \$15058_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"1") & 
                                  eclat_if(work.Int.lt(\$15058_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & 
                                  eclat_if(work.Int.ge(\$15044_binop_int6435906_arg\(48 to 78), \$15058_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$15044_binop_int6435906_result\ := work.Int.add(\$15044_binop_int6435906_arg\(32 to 47), X"000" & X"1") & \$15062_res\ & eclat_true & 
                  work.Int.sub(\$15044_binop_int6435906_arg\(80 to 95), X"000" & X"1") & \$15044_binop_int6435906_arg\(96 to 151) & \$15044_binop_int6435906_arg\(152 to 153);
                  result6468 := \$15044_binop_int6435906_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when others =>
                  \$15062_res\ := "000"& X"000000" & X"0";
                  \$15044_binop_int6435906_result\ := work.Int.add(\$15044_binop_int6435906_arg\(32 to 47), X"000" & X"1") & \$15062_res\ & eclat_true & 
                  work.Int.sub(\$15044_binop_int6435906_arg\(80 to 95), X"000" & X"1") & \$15044_binop_int6435906_arg\(96 to 151) & \$15044_binop_int6435906_arg\(152 to 153);
                  result6468 := \$15044_binop_int6435906_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                end case;
              when PAUSE_GET7088 =>
                \$15138_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7087\ := \$15124_binop_int6435907_arg\(0 to 31);
                case \$v7087\ is
                when X"0000000" & X"0" =>
                  \$15142_res\ := work.Int.add(\$15124_binop_int6435907_arg\(48 to 78), \$15138_v\(0 to 30));
                  \$15124_binop_int6435907_result\ := work.Int.add(\$15124_binop_int6435907_arg\(32 to 47), X"000" & X"1") & \$15142_res\ & eclat_true & 
                  work.Int.sub(\$15124_binop_int6435907_arg\(80 to 95), X"000" & X"1") & \$15124_binop_int6435907_arg\(96 to 151) & \$15124_binop_int6435907_arg\(152 to 153);
                  result6468 := \$15124_binop_int6435907_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"1" =>
                  \$15142_res\ := work.Int.sub(\$15124_binop_int6435907_arg\(48 to 78), \$15138_v\(0 to 30));
                  \$15124_binop_int6435907_result\ := work.Int.add(\$15124_binop_int6435907_arg\(32 to 47), X"000" & X"1") & \$15142_res\ & eclat_true & 
                  work.Int.sub(\$15124_binop_int6435907_arg\(80 to 95), X"000" & X"1") & \$15124_binop_int6435907_arg\(96 to 151) & \$15124_binop_int6435907_arg\(152 to 153);
                  result6468 := \$15124_binop_int6435907_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"2" =>
                  \$15142_res\ := work.Int.mul(\$15124_binop_int6435907_arg\(48 to 78), \$15138_v\(0 to 30));
                  \$15124_binop_int6435907_result\ := work.Int.add(\$15124_binop_int6435907_arg\(32 to 47), X"000" & X"1") & \$15142_res\ & eclat_true & 
                  work.Int.sub(\$15124_binop_int6435907_arg\(80 to 95), X"000" & X"1") & \$15124_binop_int6435907_arg\(96 to 151) & \$15124_binop_int6435907_arg\(152 to 153);
                  result6468 := \$15124_binop_int6435907_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"3" =>
                  \$v7083\ := work.Int.eq(\$15138_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v7083\(0) = '1' then
                    \$15142_res\ := "000"& X"000000" & X"0";
                    \$15124_binop_int6435907_result\ := work.Int.add(
                                                        \$15124_binop_int6435907_arg\(32 to 47), X"000" & X"1") & \$15142_res\ & eclat_true & 
                    work.Int.sub(\$15124_binop_int6435907_arg\(80 to 95), X"000" & X"1") & \$15124_binop_int6435907_arg\(96 to 151) & \$15124_binop_int6435907_arg\(152 to 153);
                    result6468 := \$15124_binop_int6435907_result\;
                    rdy6469 := eclat_true;
                    state_var7460 := IDLE6470;
                  else
                    \$15149_modulo6685895_id\ := "000001100111";
                    \$15149_modulo6685895_arg\ := work.Int.absv(\$15124_binop_int6435907_arg\(48 to 78)) & 
                    work.Int.absv(\$15138_v\(0 to 30));
                    state_var7460 := \$15149_MODULO6685895\;
                  end if;
                when X"0000000" & X"4" =>
                  \$v7086\ := work.Int.eq(\$15138_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v7086\(0) = '1' then
                    \$15142_res\ := "000"& X"000000" & X"0";
                    \$15124_binop_int6435907_result\ := work.Int.add(
                                                        \$15124_binop_int6435907_arg\(32 to 47), X"000" & X"1") & \$15142_res\ & eclat_true & 
                    work.Int.sub(\$15124_binop_int6435907_arg\(80 to 95), X"000" & X"1") & \$15124_binop_int6435907_arg\(96 to 151) & \$15124_binop_int6435907_arg\(152 to 153);
                    result6468 := \$15124_binop_int6435907_result\;
                    rdy6469 := eclat_true;
                    state_var7460 := IDLE6470;
                  else
                    \$15173_modulo6685896_id\ := "000001101001";
                    \$15173_modulo6685896_arg\ := work.Int.absv(\$15124_binop_int6435907_arg\(48 to 78)) & 
                    work.Int.absv(\$15138_v\(0 to 30));
                    state_var7460 := \$15173_MODULO6685896\;
                  end if;
                when X"0000000" & X"5" =>
                  \$15142_res\ := work.Int.land(\$15124_binop_int6435907_arg\(48 to 78), \$15138_v\(0 to 30));
                  \$15124_binop_int6435907_result\ := work.Int.add(\$15124_binop_int6435907_arg\(32 to 47), X"000" & X"1") & \$15142_res\ & eclat_true & 
                  work.Int.sub(\$15124_binop_int6435907_arg\(80 to 95), X"000" & X"1") & \$15124_binop_int6435907_arg\(96 to 151) & \$15124_binop_int6435907_arg\(152 to 153);
                  result6468 := \$15124_binop_int6435907_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"6" =>
                  \$15142_res\ := work.Int.lor(\$15124_binop_int6435907_arg\(48 to 78), \$15138_v\(0 to 30));
                  \$15124_binop_int6435907_result\ := work.Int.add(\$15124_binop_int6435907_arg\(32 to 47), X"000" & X"1") & \$15142_res\ & eclat_true & 
                  work.Int.sub(\$15124_binop_int6435907_arg\(80 to 95), X"000" & X"1") & \$15124_binop_int6435907_arg\(96 to 151) & \$15124_binop_int6435907_arg\(152 to 153);
                  result6468 := \$15124_binop_int6435907_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"7" =>
                  \$15142_res\ := work.Int.lxor(\$15124_binop_int6435907_arg\(48 to 78), \$15138_v\(0 to 30));
                  \$15124_binop_int6435907_result\ := work.Int.add(\$15124_binop_int6435907_arg\(32 to 47), X"000" & X"1") & \$15142_res\ & eclat_true & 
                  work.Int.sub(\$15124_binop_int6435907_arg\(80 to 95), X"000" & X"1") & \$15124_binop_int6435907_arg\(96 to 151) & \$15124_binop_int6435907_arg\(152 to 153);
                  result6468 := \$15124_binop_int6435907_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"8" =>
                  \$15142_res\ := work.Int.lsl(\$15124_binop_int6435907_arg\(48 to 78), \$15138_v\(0 to 30));
                  \$15124_binop_int6435907_result\ := work.Int.add(\$15124_binop_int6435907_arg\(32 to 47), X"000" & X"1") & \$15142_res\ & eclat_true & 
                  work.Int.sub(\$15124_binop_int6435907_arg\(80 to 95), X"000" & X"1") & \$15124_binop_int6435907_arg\(96 to 151) & \$15124_binop_int6435907_arg\(152 to 153);
                  result6468 := \$15124_binop_int6435907_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"9" =>
                  \$15142_res\ := work.Int.lsr(\$15124_binop_int6435907_arg\(48 to 78), \$15138_v\(0 to 30));
                  \$15124_binop_int6435907_result\ := work.Int.add(\$15124_binop_int6435907_arg\(32 to 47), X"000" & X"1") & \$15142_res\ & eclat_true & 
                  work.Int.sub(\$15124_binop_int6435907_arg\(80 to 95), X"000" & X"1") & \$15124_binop_int6435907_arg\(96 to 151) & \$15124_binop_int6435907_arg\(152 to 153);
                  result6468 := \$15124_binop_int6435907_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"a" =>
                  \$15142_res\ := work.Int.asr(\$15124_binop_int6435907_arg\(48 to 78), \$15138_v\(0 to 30));
                  \$15124_binop_int6435907_result\ := work.Int.add(\$15124_binop_int6435907_arg\(32 to 47), X"000" & X"1") & \$15142_res\ & eclat_true & 
                  work.Int.sub(\$15124_binop_int6435907_arg\(80 to 95), X"000" & X"1") & \$15124_binop_int6435907_arg\(96 to 151) & \$15124_binop_int6435907_arg\(152 to 153);
                  result6468 := \$15124_binop_int6435907_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"b" =>
                  \$15142_res\ := eclat_if(work.Int.lt(\$15124_binop_int6435907_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$15138_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.gt(\$15124_binop_int6435907_arg\(48 to 78), \$15138_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$15138_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"0" & 
                                  eclat_if(work.Int.lt(\$15124_binop_int6435907_arg\(48 to 78), \$15138_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$15124_binop_int6435907_result\ := work.Int.add(\$15124_binop_int6435907_arg\(32 to 47), X"000" & X"1") & \$15142_res\ & eclat_true & 
                  work.Int.sub(\$15124_binop_int6435907_arg\(80 to 95), X"000" & X"1") & \$15124_binop_int6435907_arg\(96 to 151) & \$15124_binop_int6435907_arg\(152 to 153);
                  result6468 := \$15124_binop_int6435907_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"c" =>
                  \$15142_res\ := eclat_if(work.Int.lt(\$15124_binop_int6435907_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$15138_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.le(\$15124_binop_int6435907_arg\(48 to 78), \$15138_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"1") & 
                                  eclat_if(work.Int.lt(\$15138_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & 
                                  eclat_if(work.Int.ge(\$15124_binop_int6435907_arg\(48 to 78), \$15138_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$15124_binop_int6435907_result\ := work.Int.add(\$15124_binop_int6435907_arg\(32 to 47), X"000" & X"1") & \$15142_res\ & eclat_true & 
                  work.Int.sub(\$15124_binop_int6435907_arg\(80 to 95), X"000" & X"1") & \$15124_binop_int6435907_arg\(96 to 151) & \$15124_binop_int6435907_arg\(152 to 153);
                  result6468 := \$15124_binop_int6435907_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when others =>
                  \$15142_res\ := "000"& X"000000" & X"0";
                  \$15124_binop_int6435907_result\ := work.Int.add(\$15124_binop_int6435907_arg\(32 to 47), X"000" & X"1") & \$15142_res\ & eclat_true & 
                  work.Int.sub(\$15124_binop_int6435907_arg\(80 to 95), X"000" & X"1") & \$15124_binop_int6435907_arg\(96 to 151) & \$15124_binop_int6435907_arg\(152 to 153);
                  result6468 := \$15124_binop_int6435907_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                end case;
              when PAUSE_GET7098 =>
                \$15218_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7097\ := \$15204_binop_int6435908_arg\(0 to 31);
                case \$v7097\ is
                when X"0000000" & X"0" =>
                  \$15222_res\ := work.Int.add(\$15204_binop_int6435908_arg\(48 to 78), \$15218_v\(0 to 30));
                  \$15204_binop_int6435908_result\ := work.Int.add(\$15204_binop_int6435908_arg\(32 to 47), X"000" & X"1") & \$15222_res\ & eclat_true & 
                  work.Int.sub(\$15204_binop_int6435908_arg\(80 to 95), X"000" & X"1") & \$15204_binop_int6435908_arg\(96 to 151) & \$15204_binop_int6435908_arg\(152 to 153);
                  result6468 := \$15204_binop_int6435908_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"1" =>
                  \$15222_res\ := work.Int.sub(\$15204_binop_int6435908_arg\(48 to 78), \$15218_v\(0 to 30));
                  \$15204_binop_int6435908_result\ := work.Int.add(\$15204_binop_int6435908_arg\(32 to 47), X"000" & X"1") & \$15222_res\ & eclat_true & 
                  work.Int.sub(\$15204_binop_int6435908_arg\(80 to 95), X"000" & X"1") & \$15204_binop_int6435908_arg\(96 to 151) & \$15204_binop_int6435908_arg\(152 to 153);
                  result6468 := \$15204_binop_int6435908_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"2" =>
                  \$15222_res\ := work.Int.mul(\$15204_binop_int6435908_arg\(48 to 78), \$15218_v\(0 to 30));
                  \$15204_binop_int6435908_result\ := work.Int.add(\$15204_binop_int6435908_arg\(32 to 47), X"000" & X"1") & \$15222_res\ & eclat_true & 
                  work.Int.sub(\$15204_binop_int6435908_arg\(80 to 95), X"000" & X"1") & \$15204_binop_int6435908_arg\(96 to 151) & \$15204_binop_int6435908_arg\(152 to 153);
                  result6468 := \$15204_binop_int6435908_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"3" =>
                  \$v7093\ := work.Int.eq(\$15218_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v7093\(0) = '1' then
                    \$15222_res\ := "000"& X"000000" & X"0";
                    \$15204_binop_int6435908_result\ := work.Int.add(
                                                        \$15204_binop_int6435908_arg\(32 to 47), X"000" & X"1") & \$15222_res\ & eclat_true & 
                    work.Int.sub(\$15204_binop_int6435908_arg\(80 to 95), X"000" & X"1") & \$15204_binop_int6435908_arg\(96 to 151) & \$15204_binop_int6435908_arg\(152 to 153);
                    result6468 := \$15204_binop_int6435908_result\;
                    rdy6469 := eclat_true;
                    state_var7460 := IDLE6470;
                  else
                    \$15229_modulo6685895_id\ := "000001101100";
                    \$15229_modulo6685895_arg\ := work.Int.absv(\$15204_binop_int6435908_arg\(48 to 78)) & 
                    work.Int.absv(\$15218_v\(0 to 30));
                    state_var7460 := \$15229_MODULO6685895\;
                  end if;
                when X"0000000" & X"4" =>
                  \$v7096\ := work.Int.eq(\$15218_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v7096\(0) = '1' then
                    \$15222_res\ := "000"& X"000000" & X"0";
                    \$15204_binop_int6435908_result\ := work.Int.add(
                                                        \$15204_binop_int6435908_arg\(32 to 47), X"000" & X"1") & \$15222_res\ & eclat_true & 
                    work.Int.sub(\$15204_binop_int6435908_arg\(80 to 95), X"000" & X"1") & \$15204_binop_int6435908_arg\(96 to 151) & \$15204_binop_int6435908_arg\(152 to 153);
                    result6468 := \$15204_binop_int6435908_result\;
                    rdy6469 := eclat_true;
                    state_var7460 := IDLE6470;
                  else
                    \$15253_modulo6685896_id\ := "000001101110";
                    \$15253_modulo6685896_arg\ := work.Int.absv(\$15204_binop_int6435908_arg\(48 to 78)) & 
                    work.Int.absv(\$15218_v\(0 to 30));
                    state_var7460 := \$15253_MODULO6685896\;
                  end if;
                when X"0000000" & X"5" =>
                  \$15222_res\ := work.Int.land(\$15204_binop_int6435908_arg\(48 to 78), \$15218_v\(0 to 30));
                  \$15204_binop_int6435908_result\ := work.Int.add(\$15204_binop_int6435908_arg\(32 to 47), X"000" & X"1") & \$15222_res\ & eclat_true & 
                  work.Int.sub(\$15204_binop_int6435908_arg\(80 to 95), X"000" & X"1") & \$15204_binop_int6435908_arg\(96 to 151) & \$15204_binop_int6435908_arg\(152 to 153);
                  result6468 := \$15204_binop_int6435908_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"6" =>
                  \$15222_res\ := work.Int.lor(\$15204_binop_int6435908_arg\(48 to 78), \$15218_v\(0 to 30));
                  \$15204_binop_int6435908_result\ := work.Int.add(\$15204_binop_int6435908_arg\(32 to 47), X"000" & X"1") & \$15222_res\ & eclat_true & 
                  work.Int.sub(\$15204_binop_int6435908_arg\(80 to 95), X"000" & X"1") & \$15204_binop_int6435908_arg\(96 to 151) & \$15204_binop_int6435908_arg\(152 to 153);
                  result6468 := \$15204_binop_int6435908_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"7" =>
                  \$15222_res\ := work.Int.lxor(\$15204_binop_int6435908_arg\(48 to 78), \$15218_v\(0 to 30));
                  \$15204_binop_int6435908_result\ := work.Int.add(\$15204_binop_int6435908_arg\(32 to 47), X"000" & X"1") & \$15222_res\ & eclat_true & 
                  work.Int.sub(\$15204_binop_int6435908_arg\(80 to 95), X"000" & X"1") & \$15204_binop_int6435908_arg\(96 to 151) & \$15204_binop_int6435908_arg\(152 to 153);
                  result6468 := \$15204_binop_int6435908_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"8" =>
                  \$15222_res\ := work.Int.lsl(\$15204_binop_int6435908_arg\(48 to 78), \$15218_v\(0 to 30));
                  \$15204_binop_int6435908_result\ := work.Int.add(\$15204_binop_int6435908_arg\(32 to 47), X"000" & X"1") & \$15222_res\ & eclat_true & 
                  work.Int.sub(\$15204_binop_int6435908_arg\(80 to 95), X"000" & X"1") & \$15204_binop_int6435908_arg\(96 to 151) & \$15204_binop_int6435908_arg\(152 to 153);
                  result6468 := \$15204_binop_int6435908_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"9" =>
                  \$15222_res\ := work.Int.lsr(\$15204_binop_int6435908_arg\(48 to 78), \$15218_v\(0 to 30));
                  \$15204_binop_int6435908_result\ := work.Int.add(\$15204_binop_int6435908_arg\(32 to 47), X"000" & X"1") & \$15222_res\ & eclat_true & 
                  work.Int.sub(\$15204_binop_int6435908_arg\(80 to 95), X"000" & X"1") & \$15204_binop_int6435908_arg\(96 to 151) & \$15204_binop_int6435908_arg\(152 to 153);
                  result6468 := \$15204_binop_int6435908_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"a" =>
                  \$15222_res\ := work.Int.asr(\$15204_binop_int6435908_arg\(48 to 78), \$15218_v\(0 to 30));
                  \$15204_binop_int6435908_result\ := work.Int.add(\$15204_binop_int6435908_arg\(32 to 47), X"000" & X"1") & \$15222_res\ & eclat_true & 
                  work.Int.sub(\$15204_binop_int6435908_arg\(80 to 95), X"000" & X"1") & \$15204_binop_int6435908_arg\(96 to 151) & \$15204_binop_int6435908_arg\(152 to 153);
                  result6468 := \$15204_binop_int6435908_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"b" =>
                  \$15222_res\ := eclat_if(work.Int.lt(\$15204_binop_int6435908_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$15218_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.gt(\$15204_binop_int6435908_arg\(48 to 78), \$15218_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$15218_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"0" & 
                                  eclat_if(work.Int.lt(\$15204_binop_int6435908_arg\(48 to 78), \$15218_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$15204_binop_int6435908_result\ := work.Int.add(\$15204_binop_int6435908_arg\(32 to 47), X"000" & X"1") & \$15222_res\ & eclat_true & 
                  work.Int.sub(\$15204_binop_int6435908_arg\(80 to 95), X"000" & X"1") & \$15204_binop_int6435908_arg\(96 to 151) & \$15204_binop_int6435908_arg\(152 to 153);
                  result6468 := \$15204_binop_int6435908_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"c" =>
                  \$15222_res\ := eclat_if(work.Int.lt(\$15204_binop_int6435908_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$15218_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.le(\$15204_binop_int6435908_arg\(48 to 78), \$15218_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"1") & 
                                  eclat_if(work.Int.lt(\$15218_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & 
                                  eclat_if(work.Int.ge(\$15204_binop_int6435908_arg\(48 to 78), \$15218_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$15204_binop_int6435908_result\ := work.Int.add(\$15204_binop_int6435908_arg\(32 to 47), X"000" & X"1") & \$15222_res\ & eclat_true & 
                  work.Int.sub(\$15204_binop_int6435908_arg\(80 to 95), X"000" & X"1") & \$15204_binop_int6435908_arg\(96 to 151) & \$15204_binop_int6435908_arg\(152 to 153);
                  result6468 := \$15204_binop_int6435908_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when others =>
                  \$15222_res\ := "000"& X"000000" & X"0";
                  \$15204_binop_int6435908_result\ := work.Int.add(\$15204_binop_int6435908_arg\(32 to 47), X"000" & X"1") & \$15222_res\ & eclat_true & 
                  work.Int.sub(\$15204_binop_int6435908_arg\(80 to 95), X"000" & X"1") & \$15204_binop_int6435908_arg\(96 to 151) & \$15204_binop_int6435908_arg\(152 to 153);
                  result6468 := \$15204_binop_int6435908_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                end case;
              when PAUSE_GET7108 =>
                \$15298_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7107\ := \$15284_binop_int6435909_arg\(0 to 31);
                case \$v7107\ is
                when X"0000000" & X"0" =>
                  \$15302_res\ := work.Int.add(\$15284_binop_int6435909_arg\(48 to 78), \$15298_v\(0 to 30));
                  \$15284_binop_int6435909_result\ := work.Int.add(\$15284_binop_int6435909_arg\(32 to 47), X"000" & X"1") & \$15302_res\ & eclat_true & 
                  work.Int.sub(\$15284_binop_int6435909_arg\(80 to 95), X"000" & X"1") & \$15284_binop_int6435909_arg\(96 to 151) & \$15284_binop_int6435909_arg\(152 to 153);
                  result6468 := \$15284_binop_int6435909_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"1" =>
                  \$15302_res\ := work.Int.sub(\$15284_binop_int6435909_arg\(48 to 78), \$15298_v\(0 to 30));
                  \$15284_binop_int6435909_result\ := work.Int.add(\$15284_binop_int6435909_arg\(32 to 47), X"000" & X"1") & \$15302_res\ & eclat_true & 
                  work.Int.sub(\$15284_binop_int6435909_arg\(80 to 95), X"000" & X"1") & \$15284_binop_int6435909_arg\(96 to 151) & \$15284_binop_int6435909_arg\(152 to 153);
                  result6468 := \$15284_binop_int6435909_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"2" =>
                  \$15302_res\ := work.Int.mul(\$15284_binop_int6435909_arg\(48 to 78), \$15298_v\(0 to 30));
                  \$15284_binop_int6435909_result\ := work.Int.add(\$15284_binop_int6435909_arg\(32 to 47), X"000" & X"1") & \$15302_res\ & eclat_true & 
                  work.Int.sub(\$15284_binop_int6435909_arg\(80 to 95), X"000" & X"1") & \$15284_binop_int6435909_arg\(96 to 151) & \$15284_binop_int6435909_arg\(152 to 153);
                  result6468 := \$15284_binop_int6435909_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"3" =>
                  \$v7103\ := work.Int.eq(\$15298_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v7103\(0) = '1' then
                    \$15302_res\ := "000"& X"000000" & X"0";
                    \$15284_binop_int6435909_result\ := work.Int.add(
                                                        \$15284_binop_int6435909_arg\(32 to 47), X"000" & X"1") & \$15302_res\ & eclat_true & 
                    work.Int.sub(\$15284_binop_int6435909_arg\(80 to 95), X"000" & X"1") & \$15284_binop_int6435909_arg\(96 to 151) & \$15284_binop_int6435909_arg\(152 to 153);
                    result6468 := \$15284_binop_int6435909_result\;
                    rdy6469 := eclat_true;
                    state_var7460 := IDLE6470;
                  else
                    \$15309_modulo6685895_id\ := "000001110001";
                    \$15309_modulo6685895_arg\ := work.Int.absv(\$15284_binop_int6435909_arg\(48 to 78)) & 
                    work.Int.absv(\$15298_v\(0 to 30));
                    state_var7460 := \$15309_MODULO6685895\;
                  end if;
                when X"0000000" & X"4" =>
                  \$v7106\ := work.Int.eq(\$15298_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v7106\(0) = '1' then
                    \$15302_res\ := "000"& X"000000" & X"0";
                    \$15284_binop_int6435909_result\ := work.Int.add(
                                                        \$15284_binop_int6435909_arg\(32 to 47), X"000" & X"1") & \$15302_res\ & eclat_true & 
                    work.Int.sub(\$15284_binop_int6435909_arg\(80 to 95), X"000" & X"1") & \$15284_binop_int6435909_arg\(96 to 151) & \$15284_binop_int6435909_arg\(152 to 153);
                    result6468 := \$15284_binop_int6435909_result\;
                    rdy6469 := eclat_true;
                    state_var7460 := IDLE6470;
                  else
                    \$15333_modulo6685896_id\ := "000001110011";
                    \$15333_modulo6685896_arg\ := work.Int.absv(\$15284_binop_int6435909_arg\(48 to 78)) & 
                    work.Int.absv(\$15298_v\(0 to 30));
                    state_var7460 := \$15333_MODULO6685896\;
                  end if;
                when X"0000000" & X"5" =>
                  \$15302_res\ := work.Int.land(\$15284_binop_int6435909_arg\(48 to 78), \$15298_v\(0 to 30));
                  \$15284_binop_int6435909_result\ := work.Int.add(\$15284_binop_int6435909_arg\(32 to 47), X"000" & X"1") & \$15302_res\ & eclat_true & 
                  work.Int.sub(\$15284_binop_int6435909_arg\(80 to 95), X"000" & X"1") & \$15284_binop_int6435909_arg\(96 to 151) & \$15284_binop_int6435909_arg\(152 to 153);
                  result6468 := \$15284_binop_int6435909_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"6" =>
                  \$15302_res\ := work.Int.lor(\$15284_binop_int6435909_arg\(48 to 78), \$15298_v\(0 to 30));
                  \$15284_binop_int6435909_result\ := work.Int.add(\$15284_binop_int6435909_arg\(32 to 47), X"000" & X"1") & \$15302_res\ & eclat_true & 
                  work.Int.sub(\$15284_binop_int6435909_arg\(80 to 95), X"000" & X"1") & \$15284_binop_int6435909_arg\(96 to 151) & \$15284_binop_int6435909_arg\(152 to 153);
                  result6468 := \$15284_binop_int6435909_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"7" =>
                  \$15302_res\ := work.Int.lxor(\$15284_binop_int6435909_arg\(48 to 78), \$15298_v\(0 to 30));
                  \$15284_binop_int6435909_result\ := work.Int.add(\$15284_binop_int6435909_arg\(32 to 47), X"000" & X"1") & \$15302_res\ & eclat_true & 
                  work.Int.sub(\$15284_binop_int6435909_arg\(80 to 95), X"000" & X"1") & \$15284_binop_int6435909_arg\(96 to 151) & \$15284_binop_int6435909_arg\(152 to 153);
                  result6468 := \$15284_binop_int6435909_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"8" =>
                  \$15302_res\ := work.Int.lsl(\$15284_binop_int6435909_arg\(48 to 78), \$15298_v\(0 to 30));
                  \$15284_binop_int6435909_result\ := work.Int.add(\$15284_binop_int6435909_arg\(32 to 47), X"000" & X"1") & \$15302_res\ & eclat_true & 
                  work.Int.sub(\$15284_binop_int6435909_arg\(80 to 95), X"000" & X"1") & \$15284_binop_int6435909_arg\(96 to 151) & \$15284_binop_int6435909_arg\(152 to 153);
                  result6468 := \$15284_binop_int6435909_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"9" =>
                  \$15302_res\ := work.Int.lsr(\$15284_binop_int6435909_arg\(48 to 78), \$15298_v\(0 to 30));
                  \$15284_binop_int6435909_result\ := work.Int.add(\$15284_binop_int6435909_arg\(32 to 47), X"000" & X"1") & \$15302_res\ & eclat_true & 
                  work.Int.sub(\$15284_binop_int6435909_arg\(80 to 95), X"000" & X"1") & \$15284_binop_int6435909_arg\(96 to 151) & \$15284_binop_int6435909_arg\(152 to 153);
                  result6468 := \$15284_binop_int6435909_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"a" =>
                  \$15302_res\ := work.Int.asr(\$15284_binop_int6435909_arg\(48 to 78), \$15298_v\(0 to 30));
                  \$15284_binop_int6435909_result\ := work.Int.add(\$15284_binop_int6435909_arg\(32 to 47), X"000" & X"1") & \$15302_res\ & eclat_true & 
                  work.Int.sub(\$15284_binop_int6435909_arg\(80 to 95), X"000" & X"1") & \$15284_binop_int6435909_arg\(96 to 151) & \$15284_binop_int6435909_arg\(152 to 153);
                  result6468 := \$15284_binop_int6435909_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"b" =>
                  \$15302_res\ := eclat_if(work.Int.lt(\$15284_binop_int6435909_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$15298_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.gt(\$15284_binop_int6435909_arg\(48 to 78), \$15298_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$15298_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"0" & 
                                  eclat_if(work.Int.lt(\$15284_binop_int6435909_arg\(48 to 78), \$15298_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$15284_binop_int6435909_result\ := work.Int.add(\$15284_binop_int6435909_arg\(32 to 47), X"000" & X"1") & \$15302_res\ & eclat_true & 
                  work.Int.sub(\$15284_binop_int6435909_arg\(80 to 95), X"000" & X"1") & \$15284_binop_int6435909_arg\(96 to 151) & \$15284_binop_int6435909_arg\(152 to 153);
                  result6468 := \$15284_binop_int6435909_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"c" =>
                  \$15302_res\ := eclat_if(work.Int.lt(\$15284_binop_int6435909_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$15298_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.le(\$15284_binop_int6435909_arg\(48 to 78), \$15298_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"1") & 
                                  eclat_if(work.Int.lt(\$15298_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & 
                                  eclat_if(work.Int.ge(\$15284_binop_int6435909_arg\(48 to 78), \$15298_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$15284_binop_int6435909_result\ := work.Int.add(\$15284_binop_int6435909_arg\(32 to 47), X"000" & X"1") & \$15302_res\ & eclat_true & 
                  work.Int.sub(\$15284_binop_int6435909_arg\(80 to 95), X"000" & X"1") & \$15284_binop_int6435909_arg\(96 to 151) & \$15284_binop_int6435909_arg\(152 to 153);
                  result6468 := \$15284_binop_int6435909_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when others =>
                  \$15302_res\ := "000"& X"000000" & X"0";
                  \$15284_binop_int6435909_result\ := work.Int.add(\$15284_binop_int6435909_arg\(32 to 47), X"000" & X"1") & \$15302_res\ & eclat_true & 
                  work.Int.sub(\$15284_binop_int6435909_arg\(80 to 95), X"000" & X"1") & \$15284_binop_int6435909_arg\(96 to 151) & \$15284_binop_int6435909_arg\(152 to 153);
                  result6468 := \$15284_binop_int6435909_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                end case;
              when PAUSE_GET7118 =>
                \$15378_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7117\ := \$15364_binop_int6435910_arg\(0 to 31);
                case \$v7117\ is
                when X"0000000" & X"0" =>
                  \$15382_res\ := work.Int.add(\$15364_binop_int6435910_arg\(48 to 78), \$15378_v\(0 to 30));
                  \$15364_binop_int6435910_result\ := work.Int.add(\$15364_binop_int6435910_arg\(32 to 47), X"000" & X"1") & \$15382_res\ & eclat_true & 
                  work.Int.sub(\$15364_binop_int6435910_arg\(80 to 95), X"000" & X"1") & \$15364_binop_int6435910_arg\(96 to 151) & \$15364_binop_int6435910_arg\(152 to 153);
                  result6468 := \$15364_binop_int6435910_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"1" =>
                  \$15382_res\ := work.Int.sub(\$15364_binop_int6435910_arg\(48 to 78), \$15378_v\(0 to 30));
                  \$15364_binop_int6435910_result\ := work.Int.add(\$15364_binop_int6435910_arg\(32 to 47), X"000" & X"1") & \$15382_res\ & eclat_true & 
                  work.Int.sub(\$15364_binop_int6435910_arg\(80 to 95), X"000" & X"1") & \$15364_binop_int6435910_arg\(96 to 151) & \$15364_binop_int6435910_arg\(152 to 153);
                  result6468 := \$15364_binop_int6435910_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"2" =>
                  \$15382_res\ := work.Int.mul(\$15364_binop_int6435910_arg\(48 to 78), \$15378_v\(0 to 30));
                  \$15364_binop_int6435910_result\ := work.Int.add(\$15364_binop_int6435910_arg\(32 to 47), X"000" & X"1") & \$15382_res\ & eclat_true & 
                  work.Int.sub(\$15364_binop_int6435910_arg\(80 to 95), X"000" & X"1") & \$15364_binop_int6435910_arg\(96 to 151) & \$15364_binop_int6435910_arg\(152 to 153);
                  result6468 := \$15364_binop_int6435910_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"3" =>
                  \$v7113\ := work.Int.eq(\$15378_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v7113\(0) = '1' then
                    \$15382_res\ := "000"& X"000000" & X"0";
                    \$15364_binop_int6435910_result\ := work.Int.add(
                                                        \$15364_binop_int6435910_arg\(32 to 47), X"000" & X"1") & \$15382_res\ & eclat_true & 
                    work.Int.sub(\$15364_binop_int6435910_arg\(80 to 95), X"000" & X"1") & \$15364_binop_int6435910_arg\(96 to 151) & \$15364_binop_int6435910_arg\(152 to 153);
                    result6468 := \$15364_binop_int6435910_result\;
                    rdy6469 := eclat_true;
                    state_var7460 := IDLE6470;
                  else
                    \$15389_modulo6685895_id\ := "000001110110";
                    \$15389_modulo6685895_arg\ := work.Int.absv(\$15364_binop_int6435910_arg\(48 to 78)) & 
                    work.Int.absv(\$15378_v\(0 to 30));
                    state_var7460 := \$15389_MODULO6685895\;
                  end if;
                when X"0000000" & X"4" =>
                  \$v7116\ := work.Int.eq(\$15378_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v7116\(0) = '1' then
                    \$15382_res\ := "000"& X"000000" & X"0";
                    \$15364_binop_int6435910_result\ := work.Int.add(
                                                        \$15364_binop_int6435910_arg\(32 to 47), X"000" & X"1") & \$15382_res\ & eclat_true & 
                    work.Int.sub(\$15364_binop_int6435910_arg\(80 to 95), X"000" & X"1") & \$15364_binop_int6435910_arg\(96 to 151) & \$15364_binop_int6435910_arg\(152 to 153);
                    result6468 := \$15364_binop_int6435910_result\;
                    rdy6469 := eclat_true;
                    state_var7460 := IDLE6470;
                  else
                    \$15413_modulo6685896_id\ := "000001111000";
                    \$15413_modulo6685896_arg\ := work.Int.absv(\$15364_binop_int6435910_arg\(48 to 78)) & 
                    work.Int.absv(\$15378_v\(0 to 30));
                    state_var7460 := \$15413_MODULO6685896\;
                  end if;
                when X"0000000" & X"5" =>
                  \$15382_res\ := work.Int.land(\$15364_binop_int6435910_arg\(48 to 78), \$15378_v\(0 to 30));
                  \$15364_binop_int6435910_result\ := work.Int.add(\$15364_binop_int6435910_arg\(32 to 47), X"000" & X"1") & \$15382_res\ & eclat_true & 
                  work.Int.sub(\$15364_binop_int6435910_arg\(80 to 95), X"000" & X"1") & \$15364_binop_int6435910_arg\(96 to 151) & \$15364_binop_int6435910_arg\(152 to 153);
                  result6468 := \$15364_binop_int6435910_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"6" =>
                  \$15382_res\ := work.Int.lor(\$15364_binop_int6435910_arg\(48 to 78), \$15378_v\(0 to 30));
                  \$15364_binop_int6435910_result\ := work.Int.add(\$15364_binop_int6435910_arg\(32 to 47), X"000" & X"1") & \$15382_res\ & eclat_true & 
                  work.Int.sub(\$15364_binop_int6435910_arg\(80 to 95), X"000" & X"1") & \$15364_binop_int6435910_arg\(96 to 151) & \$15364_binop_int6435910_arg\(152 to 153);
                  result6468 := \$15364_binop_int6435910_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"7" =>
                  \$15382_res\ := work.Int.lxor(\$15364_binop_int6435910_arg\(48 to 78), \$15378_v\(0 to 30));
                  \$15364_binop_int6435910_result\ := work.Int.add(\$15364_binop_int6435910_arg\(32 to 47), X"000" & X"1") & \$15382_res\ & eclat_true & 
                  work.Int.sub(\$15364_binop_int6435910_arg\(80 to 95), X"000" & X"1") & \$15364_binop_int6435910_arg\(96 to 151) & \$15364_binop_int6435910_arg\(152 to 153);
                  result6468 := \$15364_binop_int6435910_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"8" =>
                  \$15382_res\ := work.Int.lsl(\$15364_binop_int6435910_arg\(48 to 78), \$15378_v\(0 to 30));
                  \$15364_binop_int6435910_result\ := work.Int.add(\$15364_binop_int6435910_arg\(32 to 47), X"000" & X"1") & \$15382_res\ & eclat_true & 
                  work.Int.sub(\$15364_binop_int6435910_arg\(80 to 95), X"000" & X"1") & \$15364_binop_int6435910_arg\(96 to 151) & \$15364_binop_int6435910_arg\(152 to 153);
                  result6468 := \$15364_binop_int6435910_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"9" =>
                  \$15382_res\ := work.Int.lsr(\$15364_binop_int6435910_arg\(48 to 78), \$15378_v\(0 to 30));
                  \$15364_binop_int6435910_result\ := work.Int.add(\$15364_binop_int6435910_arg\(32 to 47), X"000" & X"1") & \$15382_res\ & eclat_true & 
                  work.Int.sub(\$15364_binop_int6435910_arg\(80 to 95), X"000" & X"1") & \$15364_binop_int6435910_arg\(96 to 151) & \$15364_binop_int6435910_arg\(152 to 153);
                  result6468 := \$15364_binop_int6435910_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"a" =>
                  \$15382_res\ := work.Int.asr(\$15364_binop_int6435910_arg\(48 to 78), \$15378_v\(0 to 30));
                  \$15364_binop_int6435910_result\ := work.Int.add(\$15364_binop_int6435910_arg\(32 to 47), X"000" & X"1") & \$15382_res\ & eclat_true & 
                  work.Int.sub(\$15364_binop_int6435910_arg\(80 to 95), X"000" & X"1") & \$15364_binop_int6435910_arg\(96 to 151) & \$15364_binop_int6435910_arg\(152 to 153);
                  result6468 := \$15364_binop_int6435910_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"b" =>
                  \$15382_res\ := eclat_if(work.Int.lt(\$15364_binop_int6435910_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$15378_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.gt(\$15364_binop_int6435910_arg\(48 to 78), \$15378_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$15378_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"0" & 
                                  eclat_if(work.Int.lt(\$15364_binop_int6435910_arg\(48 to 78), \$15378_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$15364_binop_int6435910_result\ := work.Int.add(\$15364_binop_int6435910_arg\(32 to 47), X"000" & X"1") & \$15382_res\ & eclat_true & 
                  work.Int.sub(\$15364_binop_int6435910_arg\(80 to 95), X"000" & X"1") & \$15364_binop_int6435910_arg\(96 to 151) & \$15364_binop_int6435910_arg\(152 to 153);
                  result6468 := \$15364_binop_int6435910_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"c" =>
                  \$15382_res\ := eclat_if(work.Int.lt(\$15364_binop_int6435910_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$15378_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.le(\$15364_binop_int6435910_arg\(48 to 78), \$15378_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"1") & 
                                  eclat_if(work.Int.lt(\$15378_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & 
                                  eclat_if(work.Int.ge(\$15364_binop_int6435910_arg\(48 to 78), \$15378_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$15364_binop_int6435910_result\ := work.Int.add(\$15364_binop_int6435910_arg\(32 to 47), X"000" & X"1") & \$15382_res\ & eclat_true & 
                  work.Int.sub(\$15364_binop_int6435910_arg\(80 to 95), X"000" & X"1") & \$15364_binop_int6435910_arg\(96 to 151) & \$15364_binop_int6435910_arg\(152 to 153);
                  result6468 := \$15364_binop_int6435910_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when others =>
                  \$15382_res\ := "000"& X"000000" & X"0";
                  \$15364_binop_int6435910_result\ := work.Int.add(\$15364_binop_int6435910_arg\(32 to 47), X"000" & X"1") & \$15382_res\ & eclat_true & 
                  work.Int.sub(\$15364_binop_int6435910_arg\(80 to 95), X"000" & X"1") & \$15364_binop_int6435910_arg\(96 to 151) & \$15364_binop_int6435910_arg\(152 to 153);
                  result6468 := \$15364_binop_int6435910_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                end case;
              when PAUSE_GET7128 =>
                \$15465_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7127\ := \$15451_binop_int6435912_arg\(0 to 31);
                case \$v7127\ is
                when X"0000000" & X"0" =>
                  \$15469_res\ := work.Int.add(\$15451_binop_int6435912_arg\(48 to 78), \$15465_v\(0 to 30));
                  \$15451_binop_int6435912_result\ := work.Int.add(\$15451_binop_int6435912_arg\(32 to 47), X"000" & X"1") & \$15469_res\ & eclat_true & 
                  work.Int.sub(\$15451_binop_int6435912_arg\(80 to 95), X"000" & X"1") & \$15451_binop_int6435912_arg\(96 to 151) & \$15451_binop_int6435912_arg\(152 to 153);
                  result6468 := \$15451_binop_int6435912_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"1" =>
                  \$15469_res\ := work.Int.sub(\$15451_binop_int6435912_arg\(48 to 78), \$15465_v\(0 to 30));
                  \$15451_binop_int6435912_result\ := work.Int.add(\$15451_binop_int6435912_arg\(32 to 47), X"000" & X"1") & \$15469_res\ & eclat_true & 
                  work.Int.sub(\$15451_binop_int6435912_arg\(80 to 95), X"000" & X"1") & \$15451_binop_int6435912_arg\(96 to 151) & \$15451_binop_int6435912_arg\(152 to 153);
                  result6468 := \$15451_binop_int6435912_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"2" =>
                  \$15469_res\ := work.Int.mul(\$15451_binop_int6435912_arg\(48 to 78), \$15465_v\(0 to 30));
                  \$15451_binop_int6435912_result\ := work.Int.add(\$15451_binop_int6435912_arg\(32 to 47), X"000" & X"1") & \$15469_res\ & eclat_true & 
                  work.Int.sub(\$15451_binop_int6435912_arg\(80 to 95), X"000" & X"1") & \$15451_binop_int6435912_arg\(96 to 151) & \$15451_binop_int6435912_arg\(152 to 153);
                  result6468 := \$15451_binop_int6435912_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"3" =>
                  \$v7123\ := work.Int.eq(\$15465_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v7123\(0) = '1' then
                    \$15469_res\ := "000"& X"000000" & X"0";
                    \$15451_binop_int6435912_result\ := work.Int.add(
                                                        \$15451_binop_int6435912_arg\(32 to 47), X"000" & X"1") & \$15469_res\ & eclat_true & 
                    work.Int.sub(\$15451_binop_int6435912_arg\(80 to 95), X"000" & X"1") & \$15451_binop_int6435912_arg\(96 to 151) & \$15451_binop_int6435912_arg\(152 to 153);
                    result6468 := \$15451_binop_int6435912_result\;
                    rdy6469 := eclat_true;
                    state_var7460 := IDLE6470;
                  else
                    \$15476_modulo6685895_id\ := "000001111100";
                    \$15476_modulo6685895_arg\ := work.Int.absv(\$15451_binop_int6435912_arg\(48 to 78)) & 
                    work.Int.absv(\$15465_v\(0 to 30));
                    state_var7460 := \$15476_MODULO6685895\;
                  end if;
                when X"0000000" & X"4" =>
                  \$v7126\ := work.Int.eq(\$15465_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v7126\(0) = '1' then
                    \$15469_res\ := "000"& X"000000" & X"0";
                    \$15451_binop_int6435912_result\ := work.Int.add(
                                                        \$15451_binop_int6435912_arg\(32 to 47), X"000" & X"1") & \$15469_res\ & eclat_true & 
                    work.Int.sub(\$15451_binop_int6435912_arg\(80 to 95), X"000" & X"1") & \$15451_binop_int6435912_arg\(96 to 151) & \$15451_binop_int6435912_arg\(152 to 153);
                    result6468 := \$15451_binop_int6435912_result\;
                    rdy6469 := eclat_true;
                    state_var7460 := IDLE6470;
                  else
                    \$15500_modulo6685896_id\ := "000001111110";
                    \$15500_modulo6685896_arg\ := work.Int.absv(\$15451_binop_int6435912_arg\(48 to 78)) & 
                    work.Int.absv(\$15465_v\(0 to 30));
                    state_var7460 := \$15500_MODULO6685896\;
                  end if;
                when X"0000000" & X"5" =>
                  \$15469_res\ := work.Int.land(\$15451_binop_int6435912_arg\(48 to 78), \$15465_v\(0 to 30));
                  \$15451_binop_int6435912_result\ := work.Int.add(\$15451_binop_int6435912_arg\(32 to 47), X"000" & X"1") & \$15469_res\ & eclat_true & 
                  work.Int.sub(\$15451_binop_int6435912_arg\(80 to 95), X"000" & X"1") & \$15451_binop_int6435912_arg\(96 to 151) & \$15451_binop_int6435912_arg\(152 to 153);
                  result6468 := \$15451_binop_int6435912_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"6" =>
                  \$15469_res\ := work.Int.lor(\$15451_binop_int6435912_arg\(48 to 78), \$15465_v\(0 to 30));
                  \$15451_binop_int6435912_result\ := work.Int.add(\$15451_binop_int6435912_arg\(32 to 47), X"000" & X"1") & \$15469_res\ & eclat_true & 
                  work.Int.sub(\$15451_binop_int6435912_arg\(80 to 95), X"000" & X"1") & \$15451_binop_int6435912_arg\(96 to 151) & \$15451_binop_int6435912_arg\(152 to 153);
                  result6468 := \$15451_binop_int6435912_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"7" =>
                  \$15469_res\ := work.Int.lxor(\$15451_binop_int6435912_arg\(48 to 78), \$15465_v\(0 to 30));
                  \$15451_binop_int6435912_result\ := work.Int.add(\$15451_binop_int6435912_arg\(32 to 47), X"000" & X"1") & \$15469_res\ & eclat_true & 
                  work.Int.sub(\$15451_binop_int6435912_arg\(80 to 95), X"000" & X"1") & \$15451_binop_int6435912_arg\(96 to 151) & \$15451_binop_int6435912_arg\(152 to 153);
                  result6468 := \$15451_binop_int6435912_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"8" =>
                  \$15469_res\ := work.Int.lsl(\$15451_binop_int6435912_arg\(48 to 78), \$15465_v\(0 to 30));
                  \$15451_binop_int6435912_result\ := work.Int.add(\$15451_binop_int6435912_arg\(32 to 47), X"000" & X"1") & \$15469_res\ & eclat_true & 
                  work.Int.sub(\$15451_binop_int6435912_arg\(80 to 95), X"000" & X"1") & \$15451_binop_int6435912_arg\(96 to 151) & \$15451_binop_int6435912_arg\(152 to 153);
                  result6468 := \$15451_binop_int6435912_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"9" =>
                  \$15469_res\ := work.Int.lsr(\$15451_binop_int6435912_arg\(48 to 78), \$15465_v\(0 to 30));
                  \$15451_binop_int6435912_result\ := work.Int.add(\$15451_binop_int6435912_arg\(32 to 47), X"000" & X"1") & \$15469_res\ & eclat_true & 
                  work.Int.sub(\$15451_binop_int6435912_arg\(80 to 95), X"000" & X"1") & \$15451_binop_int6435912_arg\(96 to 151) & \$15451_binop_int6435912_arg\(152 to 153);
                  result6468 := \$15451_binop_int6435912_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"a" =>
                  \$15469_res\ := work.Int.asr(\$15451_binop_int6435912_arg\(48 to 78), \$15465_v\(0 to 30));
                  \$15451_binop_int6435912_result\ := work.Int.add(\$15451_binop_int6435912_arg\(32 to 47), X"000" & X"1") & \$15469_res\ & eclat_true & 
                  work.Int.sub(\$15451_binop_int6435912_arg\(80 to 95), X"000" & X"1") & \$15451_binop_int6435912_arg\(96 to 151) & \$15451_binop_int6435912_arg\(152 to 153);
                  result6468 := \$15451_binop_int6435912_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"b" =>
                  \$15469_res\ := eclat_if(work.Int.lt(\$15451_binop_int6435912_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$15465_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.gt(\$15451_binop_int6435912_arg\(48 to 78), \$15465_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$15465_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"0" & 
                                  eclat_if(work.Int.lt(\$15451_binop_int6435912_arg\(48 to 78), \$15465_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$15451_binop_int6435912_result\ := work.Int.add(\$15451_binop_int6435912_arg\(32 to 47), X"000" & X"1") & \$15469_res\ & eclat_true & 
                  work.Int.sub(\$15451_binop_int6435912_arg\(80 to 95), X"000" & X"1") & \$15451_binop_int6435912_arg\(96 to 151) & \$15451_binop_int6435912_arg\(152 to 153);
                  result6468 := \$15451_binop_int6435912_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"c" =>
                  \$15469_res\ := eclat_if(work.Int.lt(\$15451_binop_int6435912_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$15465_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.le(\$15451_binop_int6435912_arg\(48 to 78), \$15465_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"1") & 
                                  eclat_if(work.Int.lt(\$15465_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & 
                                  eclat_if(work.Int.ge(\$15451_binop_int6435912_arg\(48 to 78), \$15465_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$15451_binop_int6435912_result\ := work.Int.add(\$15451_binop_int6435912_arg\(32 to 47), X"000" & X"1") & \$15469_res\ & eclat_true & 
                  work.Int.sub(\$15451_binop_int6435912_arg\(80 to 95), X"000" & X"1") & \$15451_binop_int6435912_arg\(96 to 151) & \$15451_binop_int6435912_arg\(152 to 153);
                  result6468 := \$15451_binop_int6435912_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when others =>
                  \$15469_res\ := "000"& X"000000" & X"0";
                  \$15451_binop_int6435912_result\ := work.Int.add(\$15451_binop_int6435912_arg\(32 to 47), X"000" & X"1") & \$15469_res\ & eclat_true & 
                  work.Int.sub(\$15451_binop_int6435912_arg\(80 to 95), X"000" & X"1") & \$15451_binop_int6435912_arg\(96 to 151) & \$15451_binop_int6435912_arg\(152 to 153);
                  result6468 := \$15451_binop_int6435912_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                end case;
              when PAUSE_GET7138 =>
                \$15545_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7137\ := \$15531_binop_int6435913_arg\(0 to 31);
                case \$v7137\ is
                when X"0000000" & X"0" =>
                  \$15549_res\ := work.Int.add(\$15531_binop_int6435913_arg\(48 to 78), \$15545_v\(0 to 30));
                  \$15531_binop_int6435913_result\ := work.Int.add(\$15531_binop_int6435913_arg\(32 to 47), X"000" & X"1") & \$15549_res\ & eclat_true & 
                  work.Int.sub(\$15531_binop_int6435913_arg\(80 to 95), X"000" & X"1") & \$15531_binop_int6435913_arg\(96 to 151) & \$15531_binop_int6435913_arg\(152 to 153);
                  result6468 := \$15531_binop_int6435913_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"1" =>
                  \$15549_res\ := work.Int.sub(\$15531_binop_int6435913_arg\(48 to 78), \$15545_v\(0 to 30));
                  \$15531_binop_int6435913_result\ := work.Int.add(\$15531_binop_int6435913_arg\(32 to 47), X"000" & X"1") & \$15549_res\ & eclat_true & 
                  work.Int.sub(\$15531_binop_int6435913_arg\(80 to 95), X"000" & X"1") & \$15531_binop_int6435913_arg\(96 to 151) & \$15531_binop_int6435913_arg\(152 to 153);
                  result6468 := \$15531_binop_int6435913_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"2" =>
                  \$15549_res\ := work.Int.mul(\$15531_binop_int6435913_arg\(48 to 78), \$15545_v\(0 to 30));
                  \$15531_binop_int6435913_result\ := work.Int.add(\$15531_binop_int6435913_arg\(32 to 47), X"000" & X"1") & \$15549_res\ & eclat_true & 
                  work.Int.sub(\$15531_binop_int6435913_arg\(80 to 95), X"000" & X"1") & \$15531_binop_int6435913_arg\(96 to 151) & \$15531_binop_int6435913_arg\(152 to 153);
                  result6468 := \$15531_binop_int6435913_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"3" =>
                  \$v7133\ := work.Int.eq(\$15545_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v7133\(0) = '1' then
                    \$15549_res\ := "000"& X"000000" & X"0";
                    \$15531_binop_int6435913_result\ := work.Int.add(
                                                        \$15531_binop_int6435913_arg\(32 to 47), X"000" & X"1") & \$15549_res\ & eclat_true & 
                    work.Int.sub(\$15531_binop_int6435913_arg\(80 to 95), X"000" & X"1") & \$15531_binop_int6435913_arg\(96 to 151) & \$15531_binop_int6435913_arg\(152 to 153);
                    result6468 := \$15531_binop_int6435913_result\;
                    rdy6469 := eclat_true;
                    state_var7460 := IDLE6470;
                  else
                    \$15556_modulo6685895_id\ := "000010000001";
                    \$15556_modulo6685895_arg\ := work.Int.absv(\$15531_binop_int6435913_arg\(48 to 78)) & 
                    work.Int.absv(\$15545_v\(0 to 30));
                    state_var7460 := \$15556_MODULO6685895\;
                  end if;
                when X"0000000" & X"4" =>
                  \$v7136\ := work.Int.eq(\$15545_v\(0 to 30), "000"& X"000000" & X"0");
                  if \$v7136\(0) = '1' then
                    \$15549_res\ := "000"& X"000000" & X"0";
                    \$15531_binop_int6435913_result\ := work.Int.add(
                                                        \$15531_binop_int6435913_arg\(32 to 47), X"000" & X"1") & \$15549_res\ & eclat_true & 
                    work.Int.sub(\$15531_binop_int6435913_arg\(80 to 95), X"000" & X"1") & \$15531_binop_int6435913_arg\(96 to 151) & \$15531_binop_int6435913_arg\(152 to 153);
                    result6468 := \$15531_binop_int6435913_result\;
                    rdy6469 := eclat_true;
                    state_var7460 := IDLE6470;
                  else
                    \$15580_modulo6685896_id\ := "000010000011";
                    \$15580_modulo6685896_arg\ := work.Int.absv(\$15531_binop_int6435913_arg\(48 to 78)) & 
                    work.Int.absv(\$15545_v\(0 to 30));
                    state_var7460 := \$15580_MODULO6685896\;
                  end if;
                when X"0000000" & X"5" =>
                  \$15549_res\ := work.Int.land(\$15531_binop_int6435913_arg\(48 to 78), \$15545_v\(0 to 30));
                  \$15531_binop_int6435913_result\ := work.Int.add(\$15531_binop_int6435913_arg\(32 to 47), X"000" & X"1") & \$15549_res\ & eclat_true & 
                  work.Int.sub(\$15531_binop_int6435913_arg\(80 to 95), X"000" & X"1") & \$15531_binop_int6435913_arg\(96 to 151) & \$15531_binop_int6435913_arg\(152 to 153);
                  result6468 := \$15531_binop_int6435913_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"6" =>
                  \$15549_res\ := work.Int.lor(\$15531_binop_int6435913_arg\(48 to 78), \$15545_v\(0 to 30));
                  \$15531_binop_int6435913_result\ := work.Int.add(\$15531_binop_int6435913_arg\(32 to 47), X"000" & X"1") & \$15549_res\ & eclat_true & 
                  work.Int.sub(\$15531_binop_int6435913_arg\(80 to 95), X"000" & X"1") & \$15531_binop_int6435913_arg\(96 to 151) & \$15531_binop_int6435913_arg\(152 to 153);
                  result6468 := \$15531_binop_int6435913_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"7" =>
                  \$15549_res\ := work.Int.lxor(\$15531_binop_int6435913_arg\(48 to 78), \$15545_v\(0 to 30));
                  \$15531_binop_int6435913_result\ := work.Int.add(\$15531_binop_int6435913_arg\(32 to 47), X"000" & X"1") & \$15549_res\ & eclat_true & 
                  work.Int.sub(\$15531_binop_int6435913_arg\(80 to 95), X"000" & X"1") & \$15531_binop_int6435913_arg\(96 to 151) & \$15531_binop_int6435913_arg\(152 to 153);
                  result6468 := \$15531_binop_int6435913_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"8" =>
                  \$15549_res\ := work.Int.lsl(\$15531_binop_int6435913_arg\(48 to 78), \$15545_v\(0 to 30));
                  \$15531_binop_int6435913_result\ := work.Int.add(\$15531_binop_int6435913_arg\(32 to 47), X"000" & X"1") & \$15549_res\ & eclat_true & 
                  work.Int.sub(\$15531_binop_int6435913_arg\(80 to 95), X"000" & X"1") & \$15531_binop_int6435913_arg\(96 to 151) & \$15531_binop_int6435913_arg\(152 to 153);
                  result6468 := \$15531_binop_int6435913_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"9" =>
                  \$15549_res\ := work.Int.lsr(\$15531_binop_int6435913_arg\(48 to 78), \$15545_v\(0 to 30));
                  \$15531_binop_int6435913_result\ := work.Int.add(\$15531_binop_int6435913_arg\(32 to 47), X"000" & X"1") & \$15549_res\ & eclat_true & 
                  work.Int.sub(\$15531_binop_int6435913_arg\(80 to 95), X"000" & X"1") & \$15531_binop_int6435913_arg\(96 to 151) & \$15531_binop_int6435913_arg\(152 to 153);
                  result6468 := \$15531_binop_int6435913_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"a" =>
                  \$15549_res\ := work.Int.asr(\$15531_binop_int6435913_arg\(48 to 78), \$15545_v\(0 to 30));
                  \$15531_binop_int6435913_result\ := work.Int.add(\$15531_binop_int6435913_arg\(32 to 47), X"000" & X"1") & \$15549_res\ & eclat_true & 
                  work.Int.sub(\$15531_binop_int6435913_arg\(80 to 95), X"000" & X"1") & \$15531_binop_int6435913_arg\(96 to 151) & \$15531_binop_int6435913_arg\(152 to 153);
                  result6468 := \$15531_binop_int6435913_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"b" =>
                  \$15549_res\ := eclat_if(work.Int.lt(\$15531_binop_int6435913_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$15545_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.gt(\$15531_binop_int6435913_arg\(48 to 78), \$15545_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$15545_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"0" & 
                                  eclat_if(work.Int.lt(\$15531_binop_int6435913_arg\(48 to 78), \$15545_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$15531_binop_int6435913_result\ := work.Int.add(\$15531_binop_int6435913_arg\(32 to 47), X"000" & X"1") & \$15549_res\ & eclat_true & 
                  work.Int.sub(\$15531_binop_int6435913_arg\(80 to 95), X"000" & X"1") & \$15531_binop_int6435913_arg\(96 to 151) & \$15531_binop_int6435913_arg\(152 to 153);
                  result6468 := \$15531_binop_int6435913_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when X"0000000" & X"c" =>
                  \$15549_res\ := eclat_if(work.Int.lt(\$15531_binop_int6435913_arg\(48 to 78), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.lt(\$15545_v\(0 to 30), "000"& X"000000" & X"0") & 
                                  eclat_if(work.Int.le(\$15531_binop_int6435913_arg\(48 to 78), \$15545_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"1") & 
                                  eclat_if(work.Int.lt(\$15545_v\(0 to 30), "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & 
                                  eclat_if(work.Int.ge(\$15531_binop_int6435913_arg\(48 to 78), \$15545_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                  \$15531_binop_int6435913_result\ := work.Int.add(\$15531_binop_int6435913_arg\(32 to 47), X"000" & X"1") & \$15549_res\ & eclat_true & 
                  work.Int.sub(\$15531_binop_int6435913_arg\(80 to 95), X"000" & X"1") & \$15531_binop_int6435913_arg\(96 to 151) & \$15531_binop_int6435913_arg\(152 to 153);
                  result6468 := \$15531_binop_int6435913_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when others =>
                  \$15549_res\ := "000"& X"000000" & X"0";
                  \$15531_binop_int6435913_result\ := work.Int.add(\$15531_binop_int6435913_arg\(32 to 47), X"000" & X"1") & \$15549_res\ & eclat_true & 
                  work.Int.sub(\$15531_binop_int6435913_arg\(80 to 95), X"000" & X"1") & \$15531_binop_int6435913_arg\(96 to 151) & \$15531_binop_int6435913_arg\(152 to 153);
                  result6468 := \$15531_binop_int6435913_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                end case;
              when PAUSE_GET7142 =>
                \$15639_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$15648_compare6445897_id\ := "000010000111";
                \$15648_compare6445897_arg\ := \$15625_binop_compare6455916_arg\(0 to 31) & \$15625_binop_compare6455916_arg\(48 to 78) & \$15639_v\(0 to 30);
                state_var7460 := \$15648_COMPARE6445897\;
              when PAUSE_GET7146 =>
                \$15675_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$15684_compare6445897_id\ := "000010001001";
                \$15684_compare6445897_arg\ := \$15661_binop_compare6455917_arg\(0 to 31) & \$15661_binop_compare6455917_arg\(48 to 78) & \$15675_v\(0 to 30);
                state_var7460 := \$15684_COMPARE6445897\;
              when PAUSE_GET7150 =>
                \$15711_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$15720_compare6445897_id\ := "000010001011";
                \$15720_compare6445897_arg\ := \$15697_binop_compare6455918_arg\(0 to 31) & \$15697_binop_compare6455918_arg\(48 to 78) & \$15711_v\(0 to 30);
                state_var7460 := \$15720_COMPARE6445897\;
              when PAUSE_GET7154 =>
                \$15747_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$15756_compare6445897_id\ := "000010001101";
                \$15756_compare6445897_arg\ := \$15733_binop_compare6455919_arg\(0 to 31) & \$15733_binop_compare6455919_arg\(48 to 78) & \$15747_v\(0 to 30);
                state_var7460 := \$15756_COMPARE6445897\;
              when PAUSE_GET7158 =>
                \$15783_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$15792_compare6445897_id\ := "000010001111";
                \$15792_compare6445897_arg\ := \$15769_binop_compare6455920_arg\(0 to 31) & \$15769_binop_compare6455920_arg\(48 to 78) & \$15783_v\(0 to 30);
                state_var7460 := \$15792_COMPARE6445897\;
              when PAUSE_GET7162 =>
                \$15819_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$15828_compare6445897_id\ := "000010010001";
                \$15828_compare6445897_arg\ := \$15805_binop_compare6455921_arg\(0 to 31) & \$15805_binop_compare6455921_arg\(48 to 78) & \$15819_v\(0 to 30);
                state_var7460 := \$15828_COMPARE6445897\;
              when PAUSE_GET7165 =>
                \$15853_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$15853_v\ & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET7168 =>
                \$15861_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"2") & \$15861_v\ & 
                work.Int.add(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET7177 =>
                \$15883\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"2") & \$15883\ & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET7180 =>
                \$15897\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"2") & \$15897\ & 
                work.Int.add(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET7195 =>
                \$15932\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := eclat_resize(\$15932\(0 to 30),16) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(16 to 47) & 
                work.Int.sub(eclat_resize(\$15851_argument1\,8), "00000001") & \$13911\(104 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET7198 =>
                \$15961\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := eclat_resize(\$15961\(0 to 30),16) & \$13911\(16 to 47) & 
                work.Int.sub(\$13911\(48 to 63), eclat_resize(\$15851_argument1\,16)) & \$13911\(16 to 47) & 
                work.Int.sub(\$13911\(96 to 103), "00000001") & \$13911\(104 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET7201 =>
                \$15981_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := eclat_resize(\$15976_v\(0 to 30),16) & \$13911\(16 to 47) & 
                work.Int.sub(work.Int.sub(work.Int.sub(work.Int.sub(\$13911\(48 to 63), eclat_resize(\$15851_argument1\,16)), X"000" & X"1"), X"000" & X"1"), X"000" & X"1") & \$15980_v\ & eclat_resize(\$15981_v\(0 to 30),8) & \$13911\(104 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET7204 =>
                \$15980_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7203\ := \$ram_lock\;
                if \$v7203\(0) = '1' then
                  state_var7460 := Q_WAIT7202;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$13911\(48 to 63), eclat_resize(\$15851_argument1\,16)), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7201;
                end if;
              when PAUSE_GET7207 =>
                \$15976_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7206\ := \$ram_lock\;
                if \$v7206\(0) = '1' then
                  state_var7460 := Q_WAIT7205;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$13911\(48 to 63), eclat_resize(\$15851_argument1\,16)), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7204;
                end if;
              when PAUSE_GET7211 =>
                \$16042_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := eclat_resize(\$16037_v\(0 to 30),16) & \$16024\(64 to 95) & 
                work.Int.sub(work.Int.sub(work.Int.sub(\$16036_sp\, X"000" & X"1"), X"000" & X"1"), X"000" & X"1") & \$16041_v\ & eclat_resize(\$16042_v\(0 to 30),8) & \$13911\(104 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET7214 =>
                \$16041_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7213\ := \$ram_lock\;
                if \$v7213\(0) = '1' then
                  state_var7460 := Q_WAIT7212;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$16036_sp\, X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7211;
                end if;
              when PAUSE_GET7217 =>
                \$16037_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7216\ := \$ram_lock\;
                if \$v7216\(0) = '1' then
                  state_var7460 := Q_WAIT7215;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$16036_sp\, X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7214;
                end if;
              when PAUSE_GET7223 =>
                \$16074_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7222\ := \$ram_lock\;
                if \$v7222\(0) = '1' then
                  state_var7460 := Q_WAIT7221;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$16063_w6515922_arg\(32 to 62),16), eclat_resize(
                                                          work.Int.add(
                                                          \$16063_w6515922_arg\(0 to 7), "00000010"),16)), X"000" & X"1")));
                  \$ram_write\ <= \$16074_v\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7220;
                end if;
              when PAUSE_GET7237 =>
                \$16121_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"2") & \$16121_v\ & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET7240 =>
                \$16127_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"2") & \$16127_v\ & 
                work.Int.add(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET7252 =>
                \$16169_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"2") & \$16169_v\ & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET7258 =>
                \$16178_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7257\ := \$ram_lock\;
                if \$v7257\(0) = '1' then
                  state_var7460 := Q_WAIT7256;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$13911\(16 to 46),16), eclat_resize(\$15851_argument1\,16)), X"000" & X"1")));
                  \$ram_write\ <= \$16178_v\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7255;
                end if;
              when PAUSE_GET7261 =>
                \$16203\ := \$code_value\;
                release(\$code_lock\);
                result6468 := work.Int.add(work.Int.add(\$13911\(0 to 15), X"000" & X"2"), eclat_resize(\$16203\,16)) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET7264 =>
                \$16217_hd\ := \$ram_value\;
                release(\$ram_lock\);
                \$16202_ofs\ := work.Int.add(eclat_resize(\$15851_argument1\,16), 
                                             work.Int.lsr(eclat_resize(\$16217_hd\(0 to 30),16), X"000000" & X"18"));
                \$v7263\ := \$code_lock\;
                if \$v7263\(0) = '1' then
                  state_var7460 := Q_WAIT7262;
                else
                  acquire(\$code_lock\);
                  \$code_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                  \$13911\(0 to 15), X"000" & X"2"), \$16202_ofs\)));
                  state_var7460 := PAUSE_GET7261;
                end if;
              when PAUSE_GET7280 =>
                \$16284_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"2") & \$16272\(0 to 31) & 
                work.Int.sub(\$16272\(80 to 95), X"000" & X"1") & \$16284_v\ & \$16272\(128 to 135) & \$16272\(136 to 151) & \$16272\(152 to 153);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET7287 =>
                \$16313_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"2") & \$16301\(0 to 31) & 
                work.Int.sub(\$16301\(80 to 95), X"000" & X"1") & \$16313_v\ & \$16301\(128 to 135) & \$16301\(136 to 151) & \$16301\(152 to 153);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET7294 =>
                \$16299_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7293\ := \$ram_lock\;
                if \$v7293\(0) = '1' then
                  state_var7460 := Q_WAIT7292;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.sub(
                                                          \$13911\(48 to 63), X"000" & X"1")));
                  \$ram_write\ <= \$13911\(64 to 95); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7291;
                end if;
              when PAUSE_GET7297 =>
                \$16349_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"2") & \$16337\(0 to 31) & 
                work.Int.sub(\$16337\(80 to 95), X"000" & X"1") & \$16349_v\ & \$16337\(128 to 135) & \$16337\(136 to 151) & \$16337\(152 to 153);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET7304 =>
                \$16335_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7303\ := \$ram_lock\;
                if \$v7303\(0) = '1' then
                  state_var7460 := Q_WAIT7302;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.sub(
                                                          work.Int.sub(
                                                          \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= \$13911\(64 to 95); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7301;
                end if;
              when PAUSE_GET7307 =>
                \$16334_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7306\ := \$ram_lock\;
                if \$v7306\(0) = '1' then
                  state_var7460 := Q_WAIT7305;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7304;
                end if;
              when PAUSE_GET7310 =>
                \$16395_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"2") & \$16383\(0 to 31) & 
                work.Int.sub(\$16383\(80 to 95), X"000" & X"1") & \$16395_v\ & \$16383\(128 to 135) & \$16383\(136 to 151) & \$16383\(152 to 153);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET7317 =>
                \$16381_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7316\ := \$ram_lock\;
                if \$v7316\(0) = '1' then
                  state_var7460 := Q_WAIT7315;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.sub(
                                                          work.Int.sub(
                                                          work.Int.sub(
                                                          \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= \$13911\(64 to 95); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7314;
                end if;
              when PAUSE_GET7320 =>
                \$16380_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7319\ := \$ram_lock\;
                if \$v7319\(0) = '1' then
                  state_var7460 := Q_WAIT7318;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7317;
                end if;
              when PAUSE_GET7323 =>
                \$16379_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7322\ := \$ram_lock\;
                if \$v7322\(0) = '1' then
                  state_var7460 := Q_WAIT7321;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7320;
                end if;
              when PAUSE_GET7326 =>
                \$16453_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"2") & \$16441\(0 to 31) & 
                work.Int.sub(\$16441\(80 to 95), X"000" & X"1") & \$16453_v\ & \$16441\(128 to 135) & \$16441\(136 to 151) & \$16441\(152 to 153);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET7333 =>
                \$16439_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7332\ := \$ram_lock\;
                if \$v7332\(0) = '1' then
                  state_var7460 := Q_WAIT7331;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.sub(
                                                          work.Int.sub(
                                                          work.Int.sub(
                                                          work.Int.sub(
                                                          \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= \$13911\(64 to 95); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7330;
                end if;
              when PAUSE_GET7336 =>
                \$16438_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7335\ := \$ram_lock\;
                if \$v7335\(0) = '1' then
                  state_var7460 := Q_WAIT7334;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7333;
                end if;
              when PAUSE_GET7339 =>
                \$16437_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7338\ := \$ram_lock\;
                if \$v7338\(0) = '1' then
                  state_var7460 := Q_WAIT7337;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7336;
                end if;
              when PAUSE_GET7342 =>
                \$16436_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7341\ := \$ram_lock\;
                if \$v7341\(0) = '1' then
                  state_var7460 := Q_WAIT7340;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7339;
                end if;
              when PAUSE_GET7351 =>
                \$16527_f0\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7350\ := \$ram_lock\;
                if \$v7350\(0) = '1' then
                  state_var7460 := Q_WAIT7349;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$13911\(16 to 46),16), X"000" & X"0"), X"000" & X"1")));
                  \$ram_write\ <= work.Int.add(\$16527_f0\(0 to 30), \$15851_argument1\) & eclat_true; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7348;
                end if;
              when PAUSE_GET7356 =>
                \$16630\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := eclat_resize(\$16630\(0 to 30),16) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(16 to 47) & 
                work.Int.sub(work.Int.add(\$13911\(96 to 103), eclat_resize(\$15851_argument1\,8)), "00000001") & \$13911\(104 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET7362 =>
                \$16673_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7361\ := \$ram_lock\;
                if \$v7361\(0) = '1' then
                  state_var7460 := Q_WAIT7360;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$16662_fill6535928_arg\(48 to 78),16), \$16662_fill6535928_arg\(0 to 15)), X"000" & X"1")));
                  \$ram_write\ <= \$16673_v\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7359;
                end if;
              when PAUSE_GET7373 =>
                \$16713_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"3") & \$16713_v\ & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET7376 =>
                \$16709\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7375\ := \$ram_lock\;
                if \$v7375\(0) = '1' then
                  state_var7460 := Q_WAIT7374;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$16709\(0 to 30),16), eclat_resize(\$16624_argument2\,16)), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7373;
                end if;
              when PAUSE_GET7379 =>
                \$16729_v\ := \$ram_value\;
                release(\$ram_lock\);
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"3") & \$16729_v\ & 
                work.Int.add(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET7382 =>
                \$16725\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7381\ := \$ram_lock\;
                if \$v7381\(0) = '1' then
                  state_var7460 := Q_WAIT7380;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$16725\(0 to 30),16), eclat_resize(\$16624_argument2\,16)), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7379;
                end if;
              when PAUSE_GET7391 =>
                \$16763_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7390\ := \$ram_lock\;
                if \$v7390\(0) = '1' then
                  state_var7460 := Q_WAIT7389;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$16752_fill6545929_arg\(48 to 78),16), \$16752_fill6545929_arg\(0 to 15)), X"000" & X"1")));
                  \$ram_write\ <= \$16763_v\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7388;
                end if;
              when PAUSE_GET7414 =>
                \$17062\ := \$code_value\;
                release(\$code_lock\);
                \$v7413\ := \$ram_lock\;
                if \$v7413\(0) = '1' then
                  state_var7460 := Q_WAIT7412;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$17048_w16565937_arg\(48 to 78),16), 
                                                          work.Int.mul(
                                                          X"000" & X"2", \$17048_w16565937_arg\(0 to 15))), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(work.Int.add(work.Int.add(
                                                            \$17048_w16565937_arg\(16 to 31), X"000" & X"2"), eclat_resize(\$17062\,16)),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7411;
                end if;
              when PAUSE_GET7424 =>
                \$17117_v\ := \$ram_value\;
                release(\$ram_lock\);
                \$v7423\ := \$ram_lock\;
                if \$v7423\(0) = '1' then
                  state_var7460 := Q_WAIT7422;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$17105_w06555936_arg\(64 to 94),16), 
                                                          work.Int.sub(
                                                          work.Int.add(
                                                          \$17105_w06555936_arg\(0 to 15), 
                                                          work.Int.mul(
                                                          X"000" & X"2", \$17105_w06555936_arg\(32 to 47))), X"000" & X"1")), X"000" & X"1")));
                  \$ram_write\ <= \$17117_v\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7421;
                end if;
              when PAUSE_GET7435 =>
                \$17165\ := \$code_value\;
                release(\$code_lock\);
                \$17166\ := work.Int.print(clk,\$17165\);
                \$17167\ := work.Print.print_newline(clk,eclat_unit);
                result6468 := \$13911\(0 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_GET7439 =>
                \$16998_argument3\ := \$code_value\;
                release(\$code_lock\);
                \$v7438\ := eclat_resize(\$13965\,8);
                case \$v7438\ is
                when "00101100" =>
                  \$v7434\ := work.Int.gt(eclat_resize(\$16624_argument2\,16), X"000" & X"0");
                  if \$v7434\(0) = '1' then
                    \$v7433\ := \$ram_lock\;
                    if \$v7433\(0) = '1' then
                      state_var7460 := Q_WAIT7432;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                      \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                      state_var7460 := PAUSE_SET7431;
                    end if;
                  else
                    \$17000_sp\ := \$13911\(48 to 63);
                    \$13923_make_block579_id\ := "000010111010";
                    \$13923_make_block579_arg\ := \$17000_sp\ & \$13911\(16 to 47) & \$13911\(64 to 95) & "11110111" & 
                    work.Int.add(work.Int.sub(work.Int.mul(X"000" & X"2", eclat_resize(\$15851_argument1\,16)), X"000" & X"1"), eclat_resize(\$16624_argument2\,16));
                    state_var7460 := \$13923_MAKE_BLOCK579\;
                  end if;
                when others =>
                  \$17164\ := work.Print.print_string(clk,of_string("unknown opcode : "));
                  \$v7437\ := \$code_lock\;
                  if \$v7437\(0) = '1' then
                    state_var7460 := Q_WAIT7436;
                  else
                    acquire(\$code_lock\);
                    \$code_ptr\ <= to_integer(unsigned(\$13911\(0 to 15)));
                    state_var7460 := PAUSE_GET7435;
                  end if;
                end case;
              when PAUSE_GET7443 =>
                \$16624_argument2\ := \$code_value\;
                release(\$code_lock\);
                \$v7442\ := eclat_resize(\$13965\,8);
                case \$v7442\ is
                when "00100100" =>
                  \$13928_w652_id\ := "000010100110";
                  \$13928_w652_arg\ := X"000" & X"1" & \$13911\(48 to 63) & eclat_resize(\$15851_argument1\,16) & eclat_resize(\$16624_argument2\,16);
                  state_var7460 := \$13928_W652\;
                when "00101011" =>
                  \$v7372\ := work.Int.gt(eclat_resize(\$15851_argument1\,16), X"000" & X"0");
                  if \$v7372\(0) = '1' then
                    \$v7371\ := \$ram_lock\;
                    if \$v7371\(0) = '1' then
                      state_var7460 := Q_WAIT7370;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                      \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                      state_var7460 := PAUSE_SET7369;
                    end if;
                  else
                    \$16650_sp\ := \$13911\(48 to 63);
                    \$13923_make_block579_id\ := "000010101000";
                    \$13923_make_block579_arg\ := \$16650_sp\ & \$13911\(16 to 47) & \$13911\(64 to 95) & "11110111" & 
                    work.Int.add(eclat_resize(\$15851_argument1\,16), X"000" & X"1");
                    state_var7460 := \$13923_MAKE_BLOCK579\;
                  end if;
                when "00110111" =>
                  \$v7378\ := \$ram_lock\;
                  if \$v7378\(0) = '1' then
                    state_var7460 := Q_WAIT7377;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(X"3e80", eclat_resize(\$15851_argument1\,16))));
                    state_var7460 := PAUSE_GET7376;
                  end if;
                when "00111000" =>
                  \$v7387\ := \$ram_lock\;
                  if \$v7387\(0) = '1' then
                    state_var7460 := Q_WAIT7386;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET7385;
                  end if;
                when "00111110" =>
                  \$13923_make_block579_id\ := "000010101010";
                  \$13923_make_block579_arg\ := \$13911\(48 to 63) & \$13911\(16 to 47) & \$13911\(64 to 95) & eclat_resize(\$16624_argument2\,8) & eclat_resize(\$15851_argument1\,16);
                  state_var7460 := \$13923_MAKE_BLOCK579\;
                when "10000011" =>
                  \$16788_compbranch6505930_id\ := "000010101100";
                  \$16788_compbranch6505930_arg\ := X"0000000" & X"0" & \$15851_argument1\ & \$16624_argument2\ & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  state_var7460 := \$16788_COMPBRANCH6505930\;
                when "10000100" =>
                  \$16823_compbranch6505931_id\ := "000010101110";
                  \$16823_compbranch6505931_arg\ := X"0000000" & X"1" & \$15851_argument1\ & \$16624_argument2\ & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  state_var7460 := \$16823_COMPBRANCH6505931\;
                when "10000101" =>
                  \$16858_compbranch6505932_id\ := "000010110000";
                  \$16858_compbranch6505932_arg\ := X"0000000" & X"2" & \$15851_argument1\ & \$16624_argument2\ & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  state_var7460 := \$16858_COMPBRANCH6505932\;
                when "10000110" =>
                  \$16893_compbranch6505933_id\ := "000010110010";
                  \$16893_compbranch6505933_arg\ := X"0000000" & X"3" & \$15851_argument1\ & \$16624_argument2\ & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  state_var7460 := \$16893_COMPBRANCH6505933\;
                when "10000111" =>
                  \$16928_compbranch6505934_id\ := "000010110100";
                  \$16928_compbranch6505934_arg\ := X"0000000" & X"4" & \$15851_argument1\ & \$16624_argument2\ & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  state_var7460 := \$16928_COMPBRANCH6505934\;
                when "10001000" =>
                  \$16963_compbranch6505935_id\ := "000010110110";
                  \$16963_compbranch6505935_arg\ := X"0000000" & X"5" & \$15851_argument1\ & \$16624_argument2\ & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  state_var7460 := \$16963_COMPBRANCH6505935\;
                when others =>
                  \$v7441\ := \$code_lock\;
                  if \$v7441\(0) = '1' then
                    state_var7460 := Q_WAIT7440;
                  else
                    acquire(\$code_lock\);
                    \$code_ptr\ <= to_integer(unsigned(work.Int.add(\$13911\(0 to 15), X"000" & X"3")));
                    state_var7460 := PAUSE_GET7439;
                  end if;
                end case;
              when PAUSE_GET7447 =>
                \$15851_argument1\ := \$code_value\;
                release(\$code_lock\);
                \$v7446\ := eclat_resize(\$13965\,8);
                case \$v7446\ is
                when "00001000" =>
                  \$v7167\ := \$ram_lock\;
                  if \$v7167\(0) = '1' then
                    state_var7460 := Q_WAIT7166;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                   \$13911\(48 to 63), eclat_resize(\$15851_argument1\,16)), X"000" & X"1")));
                    state_var7460 := PAUSE_GET7165;
                  end if;
                when "00010010" =>
                  \$v7173\ := \$ram_lock\;
                  if \$v7173\(0) = '1' then
                    state_var7460 := Q_WAIT7172;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET7171;
                  end if;
                when "00010011" =>
                  result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"2") & \$13911\(16 to 47) & 
                  work.Int.sub(\$13911\(48 to 63), eclat_resize(\$15851_argument1\,16)) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when "00010100" =>
                  \$v7176\ := \$ram_lock\;
                  if \$v7176\(0) = '1' then
                    state_var7460 := Q_WAIT7175;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.sub(
                                                            work.Int.sub(
                                                            \$13911\(48 to 63), X"000" & X"1"), eclat_resize(\$15851_argument1\,16))));
                    \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET7174;
                  end if;
                when "00011001" =>
                  \$v7179\ := \$ram_lock\;
                  if \$v7179\(0) = '1' then
                    state_var7460 := Q_WAIT7178;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$13911\(64 to 94),16), 
                                                                   work.Int.sub(
                                                                   eclat_resize(\$15851_argument1\,16), X"000" & X"1")), X"000" & X"1")));
                    state_var7460 := PAUSE_GET7177;
                  end if;
                when "00011110" =>
                  \$v7185\ := \$ram_lock\;
                  if \$v7185\(0) = '1' then
                    state_var7460 := Q_WAIT7184;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET7183;
                  end if;
                when "00011111" =>
                  \$v7194\ := \$ram_lock\;
                  if \$v7194\(0) = '1' then
                    state_var7460 := Q_WAIT7193;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= eclat_resize(\$13911\(96 to 103),31) & eclat_true; \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET7192;
                  end if;
                when "00100000" =>
                  \$v7197\ := \$ram_lock\;
                  if \$v7197\(0) = '1' then
                    state_var7460 := Q_WAIT7196;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$13911\(16 to 46),16), X"000" & X"0"), X"000" & X"1")));
                    state_var7460 := PAUSE_GET7195;
                  end if;
                when "00100101" =>
                  \$13924_apply638_id\ := "000010010011";
                  \$13924_apply638_arg\ := eclat_true & eclat_false & eclat_false & \$13911\(96 to 103) & eclat_true & eclat_resize(\$15851_argument1\,16) & X"000" & X"1" & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(120 to 121) & \$13911\(64 to 95) & \$13911\(96 to 103) & \$13911\(104 to 119);
                  state_var7460 := \$13924_APPLY638\;
                when "00100110" =>
                  \$13924_apply638_id\ := "000010010100";
                  \$13924_apply638_arg\ := eclat_true & eclat_true & eclat_false & 
                  work.Int.add(\$13911\(96 to 103), "00000001") & eclat_true & eclat_resize(\$15851_argument1\,16) & X"000" & X"2" & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(120 to 121) & \$13911\(64 to 95) & \$13911\(96 to 103) & \$13911\(104 to 119);
                  state_var7460 := \$13924_APPLY638\;
                when "00100111" =>
                  \$13924_apply638_id\ := "000010010101";
                  \$13924_apply638_arg\ := eclat_true & eclat_true & eclat_true & 
                  work.Int.add(\$13911\(96 to 103), "00000010") & eclat_true & eclat_resize(\$15851_argument1\,16) & X"000" & X"3" & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(120 to 121) & \$13911\(64 to 95) & \$13911\(96 to 103) & \$13911\(104 to 119);
                  state_var7460 := \$13924_APPLY638\;
                when "00101000" =>
                  \$v7210\ := work.Int.gt(\$13911\(96 to 103), "00000000");
                  if \$v7210\(0) = '1' then
                    \$v7200\ := \$ram_lock\;
                    if \$v7200\(0) = '1' then
                      state_var7460 := Q_WAIT7199;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                        work.Int.add(
                                                        eclat_resize(\$13911\(16 to 46),16), X"000" & X"0"), X"000" & X"1")));
                      state_var7460 := PAUSE_GET7198;
                    end if;
                  else
                    \$v7209\ := \$ram_lock\;
                    if \$v7209\(0) = '1' then
                      state_var7460 := Q_WAIT7208;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(
                                                        work.Int.sub(
                                                        \$13911\(48 to 63), eclat_resize(\$15851_argument1\,16)), X"000" & X"1")));
                      state_var7460 := PAUSE_GET7207;
                    end if;
                  end if;
                when "00101010" =>
                  \$v7233\ := work.Int.ge(\$13911\(96 to 103), eclat_resize(\$15851_argument1\,8));
                  if \$v7233\(0) = '1' then
                    result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"2") & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 95) & 
                    work.Int.sub(\$13911\(96 to 103), eclat_resize(\$15851_argument1\,8)) & \$13911\(104 to 119) & \$13911\(120 to 121);
                    rdy6469 := eclat_true;
                    state_var7460 := IDLE6470;
                  else
                    \$13923_make_block579_id\ := "000010010111";
                    \$13923_make_block579_arg\ := \$13911\(48 to 63) & \$13911\(16 to 47) & \$13911\(64 to 95) & "11110111" & eclat_resize(
                    work.Int.add(\$13911\(96 to 103), "00000011"),16);
                    state_var7460 := \$13923_MAKE_BLOCK579\;
                  end if;
                when "00110000" =>
                  \$13925_offsetclosure_n639_id\ := "000010011000";
                  \$13925_offsetclosure_n639_arg\ := work.Int.add(\$13911\(0 to 15), X"000" & X"2") & \$13911\(48 to 63) & eclat_resize(\$15851_argument1\,16) & \$13911\(64 to 119) & \$13911\(120 to 121) & \$13911\(64 to 95);
                  state_var7460 := \$13925_OFFSETCLOSURE_N639\;
                when "00110100" =>
                  \$v7236\ := \$ram_lock\;
                  if \$v7236\(0) = '1' then
                    state_var7460 := Q_WAIT7235;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET7234;
                  end if;
                when "00110101" =>
                  \$v7239\ := \$ram_lock\;
                  if \$v7239\(0) = '1' then
                    state_var7460 := Q_WAIT7238;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(X"3e80", eclat_resize(\$15851_argument1\,16))));
                    state_var7460 := PAUSE_GET7237;
                  end if;
                when "00110110" =>
                  \$v7245\ := \$ram_lock\;
                  if \$v7245\(0) = '1' then
                    state_var7460 := Q_WAIT7244;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET7243;
                  end if;
                when "00111001" =>
                  \$v7248\ := \$ram_lock\;
                  if \$v7248\(0) = '1' then
                    state_var7460 := Q_WAIT7247;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            X"3e80", eclat_resize(\$15851_argument1\,16))));
                    \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET7246;
                  end if;
                when "00111011" =>
                  \$13926_make_block_n646_id\ := "000010011010";
                  \$13926_make_block_n646_arg\ := work.Int.add(\$13911\(0 to 15), X"000" & X"2") & \$13911\(48 to 63) & eclat_false & eclat_false & eclat_false & \$15851_argument1\ & X"000" & X"0" & \$13911\(16 to 47) & \$13911\(120 to 121) & \$13911\(64 to 95) & \$13911\(96 to 103) & \$13911\(104 to 119);
                  state_var7460 := \$13926_MAKE_BLOCK_N646\;
                when "00111101" =>
                  \$v7251\ := \$ram_lock\;
                  if \$v7251\(0) = '1' then
                    state_var7460 := Q_WAIT7250;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET7249;
                  end if;
                when "00111111" =>
                  \$13926_make_block_n646_id\ := "000010011100";
                  \$13926_make_block_n646_arg\ := work.Int.add(\$13911\(0 to 15), X"000" & X"2") & \$13911\(48 to 63) & eclat_true & eclat_false & eclat_false & \$15851_argument1\ & X"000" & X"1" & \$13911\(16 to 47) & \$13911\(120 to 121) & \$13911\(64 to 95) & \$13911\(96 to 103) & \$13911\(104 to 119);
                  state_var7460 := \$13926_MAKE_BLOCK_N646\;
                when "01000000" =>
                  \$13926_make_block_n646_id\ := "000010011101";
                  \$13926_make_block_n646_arg\ := work.Int.add(\$13911\(0 to 15), X"000" & X"2") & \$13911\(48 to 63) & eclat_true & eclat_true & eclat_false & \$15851_argument1\ & X"000" & X"2" & \$13911\(16 to 47) & \$13911\(120 to 121) & \$13911\(64 to 95) & \$13911\(96 to 103) & \$13911\(104 to 119);
                  state_var7460 := \$13926_MAKE_BLOCK_N646\;
                when "01000001" =>
                  \$13926_make_block_n646_id\ := "000010011110";
                  \$13926_make_block_n646_arg\ := work.Int.add(\$13911\(0 to 15), X"000" & X"2") & \$13911\(48 to 63) & eclat_true & eclat_true & eclat_true & \$15851_argument1\ & X"000" & X"3" & \$13911\(16 to 47) & \$13911\(120 to 121) & \$13911\(64 to 95) & \$13911\(96 to 103) & \$13911\(104 to 119);
                  state_var7460 := \$13926_MAKE_BLOCK_N646\;
                when "01000010" =>
                  \$16155\ := work.Print.print_string(clk,of_string("fatal error: "));
                  \$16156\ := work.Print.print_string(clk,of_string("unsupported instruction SETFLOATFIELD"));
                  \$16157\ := work.Print.print_newline(clk,eclat_unit);
                  \$16158_forever6705923_id\ := "000010011111";
                  \$16158_forever6705923_arg\ := eclat_unit;
                  state_var7460 := \$16158_FOREVER6705923\;
                when "01000111" =>
                  \$16165\ := work.Assertion.ok(work.Bool.lnot(""&\$13911\(47)));
                  \$v7254\ := \$ram_lock\;
                  if \$v7254\(0) = '1' then
                    state_var7460 := Q_WAIT7253;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$13911\(16 to 46),16), eclat_resize(\$15851_argument1\,16)), X"000" & X"1")));
                    state_var7460 := PAUSE_GET7252;
                  end if;
                when "01001101" =>
                  \$v7260\ := \$ram_lock\;
                  if \$v7260\(0) = '1' then
                    state_var7460 := Q_WAIT7259;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13911\(48 to 63), X"000" & X"1")));
                    state_var7460 := PAUSE_GET7258;
                  end if;
                when "01001110" =>
                  \$16192\ := work.Print.print_string(clk,of_string("fatal error: "));
                  \$16193\ := work.Print.print_string(clk,of_string("unsupported instruction SETFLOATFIELD"));
                  \$16194\ := work.Print.print_newline(clk,eclat_unit);
                  \$16195_forever6705924_id\ := "000010100000";
                  \$16195_forever6705924_arg\ := eclat_unit;
                  state_var7460 := \$16195_FOREVER6705924\;
                when "01010111" =>
                  \$v7267\ := ""&\$13911\(47);
                  if \$v7267\(0) = '1' then
                    \$16202_ofs\ := eclat_resize(\$13911\(16 to 46),16);
                    \$v7263\ := \$code_lock\;
                    if \$v7263\(0) = '1' then
                      state_var7460 := Q_WAIT7262;
                    else
                      acquire(\$code_lock\);
                      \$code_ptr\ <= to_integer(unsigned(work.Int.add(
                                                         work.Int.add(
                                                         \$13911\(0 to 15), X"000" & X"2"), \$16202_ofs\)));
                      state_var7460 := PAUSE_GET7261;
                    end if;
                  else
                    \$v7266\ := \$ram_lock\;
                    if \$v7266\(0) = '1' then
                      state_var7460 := Q_WAIT7265;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$13911\(16 to 46),16)));
                      state_var7460 := PAUSE_GET7264;
                    end if;
                  end if;
                when "01010100" =>
                  result6468 := work.Int.add(work.Int.add(\$13911\(0 to 15), X"000" & X"1"), eclat_resize(\$15851_argument1\,16)) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when "01011001" =>
                  \$v7279\ := \$ram_lock\;
                  if \$v7279\(0) = '1' then
                    state_var7460 := Q_WAIT7278;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= eclat_resize(\$13911\(96 to 103),31) & eclat_true; \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET7277;
                  end if;
                when "01011100" =>
                  result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 95) & \$13911\(96 to 103) & \$13911\(104 to 119) & \$13911\(120 to 121);
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when "01011101" =>
                  \$v7286\ := \$ram_lock\;
                  if \$v7286\(0) = '1' then
                    state_var7460 := Q_WAIT7285;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= \$13911\(64 to 95); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET7284;
                  end if;
                when "01011110" =>
                  \$v7296\ := \$ram_lock\;
                  if \$v7296\(0) = '1' then
                    state_var7460 := Q_WAIT7295;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13911\(48 to 63), X"000" & X"1")));
                    state_var7460 := PAUSE_GET7294;
                  end if;
                when "01011111" =>
                  \$v7309\ := \$ram_lock\;
                  if \$v7309\(0) = '1' then
                    state_var7460 := Q_WAIT7308;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13911\(48 to 63), X"000" & X"1")));
                    state_var7460 := PAUSE_GET7307;
                  end if;
                when "01100000" =>
                  \$v7325\ := \$ram_lock\;
                  if \$v7325\(0) = '1' then
                    state_var7460 := Q_WAIT7324;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13911\(48 to 63), X"000" & X"1")));
                    state_var7460 := PAUSE_GET7323;
                  end if;
                when "01100001" =>
                  \$v7344\ := \$ram_lock\;
                  if \$v7344\(0) = '1' then
                    state_var7460 := Q_WAIT7343;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13911\(48 to 63), X"000" & X"1")));
                    state_var7460 := PAUSE_GET7342;
                  end if;
                when "01100010" =>
                  \$16507\ := work.Print.print_string(clk,of_string("fatal error: "));
                  \$16508\ := work.Print.print_string(clk,of_string("unsupported instruction CALLN"));
                  \$16509\ := work.Print.print_newline(clk,eclat_unit);
                  \$16510_forever6705925_id\ := "000010100001";
                  \$16510_forever6705925_arg\ := eclat_unit;
                  state_var7460 := \$16510_FOREVER6705925\;
                when "01100111" =>
                  result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"2") & \$15851_argument1\ & eclat_true & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when "01101100" =>
                  \$v7347\ := \$ram_lock\;
                  if \$v7347\(0) = '1' then
                    state_var7460 := Q_WAIT7346;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET7345;
                  end if;
                when "01111111" =>
                  result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"2") & 
                  work.Int.add(\$13911\(16 to 46), \$15851_argument1\) & eclat_true & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when "10000000" =>
                  \$v7353\ := \$ram_lock\;
                  if \$v7353\(0) = '1' then
                    state_var7460 := Q_WAIT7352;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$13911\(16 to 46),16), X"000" & X"0"), X"000" & X"1")));
                    state_var7460 := PAUSE_GET7351;
                  end if;
                when "10001011" =>
                  \$16551_compbranch6505926_id\ := "000010100011";
                  \$16551_compbranch6505926_arg\ := X"0000000" & X"2" & \$15851_argument1\ & \$13911\(16 to 46) & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  state_var7460 := \$16551_COMPBRANCH6505926\;
                when "10001100" =>
                  \$16589_compbranch6505927_id\ := "000010100101";
                  \$16589_compbranch6505927_arg\ := X"0000000" & X"5" & \$15851_argument1\ & \$13911\(16 to 46) & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  state_var7460 := \$16589_COMPBRANCH6505927\;
                when others =>
                  \$v7445\ := \$code_lock\;
                  if \$v7445\(0) = '1' then
                    state_var7460 := Q_WAIT7444;
                  else
                    acquire(\$code_lock\);
                    \$code_ptr\ <= to_integer(unsigned(work.Int.add(\$13911\(0 to 15), X"000" & X"2")));
                    state_var7460 := PAUSE_GET7443;
                  end if;
                end case;
              when PAUSE_GET7451 =>
                \$13965\ := \$code_value\;
                release(\$code_lock\);
                \$v7450\ := eclat_resize(\$13965\,8);
                case \$v7450\ is
                when "00000000" =>
                  \$v6784\ := \$ram_lock\;
                  if \$v6784\(0) = '1' then
                    state_var7460 := Q_WAIT6783;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                   \$13911\(48 to 63), X"000" & X"0"), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6782;
                  end if;
                when "00000001" =>
                  \$v6787\ := \$ram_lock\;
                  if \$v6787\(0) = '1' then
                    state_var7460 := Q_WAIT6786;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                   \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6785;
                  end if;
                when "00000010" =>
                  \$v6790\ := \$ram_lock\;
                  if \$v6790\(0) = '1' then
                    state_var7460 := Q_WAIT6789;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                   \$13911\(48 to 63), X"000" & X"2"), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6788;
                  end if;
                when "00000011" =>
                  \$v6793\ := \$ram_lock\;
                  if \$v6793\(0) = '1' then
                    state_var7460 := Q_WAIT6792;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                   \$13911\(48 to 63), X"000" & X"3"), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6791;
                  end if;
                when "00000100" =>
                  \$v6796\ := \$ram_lock\;
                  if \$v6796\(0) = '1' then
                    state_var7460 := Q_WAIT6795;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                   \$13911\(48 to 63), X"000" & X"4"), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6794;
                  end if;
                when "00000101" =>
                  \$v6799\ := \$ram_lock\;
                  if \$v6799\(0) = '1' then
                    state_var7460 := Q_WAIT6798;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                   \$13911\(48 to 63), X"000" & X"5"), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6797;
                  end if;
                when "00000110" =>
                  \$v6802\ := \$ram_lock\;
                  if \$v6802\(0) = '1' then
                    state_var7460 := Q_WAIT6801;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                   \$13911\(48 to 63), X"000" & X"6"), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6800;
                  end if;
                when "00000111" =>
                  \$v6805\ := \$ram_lock\;
                  if \$v6805\(0) = '1' then
                    state_var7460 := Q_WAIT6804;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                   \$13911\(48 to 63), X"000" & X"7"), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6803;
                  end if;
                when "00001001" =>
                  \$v6808\ := \$ram_lock\;
                  if \$v6808\(0) = '1' then
                    state_var7460 := Q_WAIT6807;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET6806;
                  end if;
                when "00001010" =>
                  \$v6811\ := \$ram_lock\;
                  if \$v6811\(0) = '1' then
                    state_var7460 := Q_WAIT6810;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET6809;
                  end if;
                when "00001011" =>
                  \$v6817\ := \$ram_lock\;
                  if \$v6817\(0) = '1' then
                    state_var7460 := Q_WAIT6816;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET6815;
                  end if;
                when "00001100" =>
                  \$v6823\ := \$ram_lock\;
                  if \$v6823\(0) = '1' then
                    state_var7460 := Q_WAIT6822;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET6821;
                  end if;
                when "00001101" =>
                  \$v6829\ := \$ram_lock\;
                  if \$v6829\(0) = '1' then
                    state_var7460 := Q_WAIT6828;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET6827;
                  end if;
                when "00001110" =>
                  \$v6835\ := \$ram_lock\;
                  if \$v6835\(0) = '1' then
                    state_var7460 := Q_WAIT6834;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET6833;
                  end if;
                when "00001111" =>
                  \$v6841\ := \$ram_lock\;
                  if \$v6841\(0) = '1' then
                    state_var7460 := Q_WAIT6840;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET6839;
                  end if;
                when "00010000" =>
                  \$v6847\ := \$ram_lock\;
                  if \$v6847\(0) = '1' then
                    state_var7460 := Q_WAIT6846;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET6845;
                  end if;
                when "00010001" =>
                  \$v6853\ := \$ram_lock\;
                  if \$v6853\(0) = '1' then
                    state_var7460 := Q_WAIT6852;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET6851;
                  end if;
                when "00010101" =>
                  \$v6856\ := \$ram_lock\;
                  if \$v6856\(0) = '1' then
                    state_var7460 := Q_WAIT6855;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$13911\(64 to 94),16), 
                                                                   work.Int.sub(
                                                                   X"000" & X"1", X"000" & X"1")), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6854;
                  end if;
                when "00010110" =>
                  \$v6859\ := \$ram_lock\;
                  if \$v6859\(0) = '1' then
                    state_var7460 := Q_WAIT6858;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$13911\(64 to 94),16), 
                                                                   work.Int.sub(
                                                                   X"000" & X"2", X"000" & X"1")), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6857;
                  end if;
                when "00010111" =>
                  \$v6862\ := \$ram_lock\;
                  if \$v6862\(0) = '1' then
                    state_var7460 := Q_WAIT6861;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$13911\(64 to 94),16), 
                                                                   work.Int.sub(
                                                                   X"000" & X"3", X"000" & X"1")), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6860;
                  end if;
                when "00011000" =>
                  \$v6865\ := \$ram_lock\;
                  if \$v6865\(0) = '1' then
                    state_var7460 := Q_WAIT6864;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$13911\(64 to 94),16), 
                                                                   work.Int.sub(
                                                                   X"000" & X"4", X"000" & X"1")), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6863;
                  end if;
                when "00011010" =>
                  \$v6871\ := \$ram_lock\;
                  if \$v6871\(0) = '1' then
                    state_var7460 := Q_WAIT6870;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET6869;
                  end if;
                when "00011011" =>
                  \$v6877\ := \$ram_lock\;
                  if \$v6877\(0) = '1' then
                    state_var7460 := Q_WAIT6876;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET6875;
                  end if;
                when "00011100" =>
                  \$v6883\ := \$ram_lock\;
                  if \$v6883\(0) = '1' then
                    state_var7460 := Q_WAIT6882;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET6881;
                  end if;
                when "00011101" =>
                  \$v6889\ := \$ram_lock\;
                  if \$v6889\(0) = '1' then
                    state_var7460 := Q_WAIT6888;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET6887;
                  end if;
                when "00100001" =>
                  \$13924_apply638_id\ := "000000110101";
                  \$13924_apply638_arg\ := eclat_true & eclat_false & eclat_false & "00000000" & eclat_false & X"000" & X"0" & X"000" & X"0" & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(120 to 121) & \$13911\(64 to 95) & \$13911\(96 to 103) & \$13911\(104 to 119);
                  state_var7460 := \$13924_APPLY638\;
                when "00100010" =>
                  \$13924_apply638_id\ := "000000110110";
                  \$13924_apply638_arg\ := eclat_true & eclat_true & eclat_false & "00000001" & eclat_false & X"000" & X"0" & X"000" & X"0" & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(120 to 121) & \$13911\(64 to 95) & \$13911\(96 to 103) & \$13911\(104 to 119);
                  state_var7460 := \$13924_APPLY638\;
                when "00100011" =>
                  \$13924_apply638_id\ := "000000110111";
                  \$13924_apply638_arg\ := eclat_true & eclat_true & eclat_true & "00000010" & eclat_false & X"000" & X"0" & X"000" & X"0" & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(120 to 121) & \$13911\(64 to 95) & \$13911\(96 to 103) & \$13911\(104 to 119);
                  state_var7460 := \$13924_APPLY638\;
                when "00101001" =>
                  \$v6902\ := \$ram_lock\;
                  if \$v6902\(0) = '1' then
                    state_var7460 := Q_WAIT6901;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$13911\(64 to 94),16)));
                    state_var7460 := PAUSE_GET6900;
                  end if;
                when "00101101" =>
                  \$13925_offsetclosure_n639_id\ := "000000111001";
                  \$13925_offsetclosure_n639_arg\ := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$13911\(48 to 63) & 
                  work.Int.neg(X"000" & X"2") & \$13911\(64 to 119) & \$13911\(120 to 121) & \$13911\(64 to 95);
                  state_var7460 := \$13925_OFFSETCLOSURE_N639\;
                when "00101110" =>
                  \$13925_offsetclosure_n639_id\ := "000000111010";
                  \$13925_offsetclosure_n639_arg\ := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$13911\(48 to 63) & X"000" & X"0" & \$13911\(64 to 119) & \$13911\(120 to 121) & \$13911\(64 to 95);
                  state_var7460 := \$13925_OFFSETCLOSURE_N639\;
                when "00101111" =>
                  \$13925_offsetclosure_n639_id\ := "000000111011";
                  \$13925_offsetclosure_n639_arg\ := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$13911\(48 to 63) & X"000" & X"2" & \$13911\(64 to 119) & \$13911\(120 to 121) & \$13911\(64 to 95);
                  state_var7460 := \$13925_OFFSETCLOSURE_N639\;
                when "00110001" =>
                  \$v6905\ := \$ram_lock\;
                  if \$v6905\(0) = '1' then
                    state_var7460 := Q_WAIT6904;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET6903;
                  end if;
                when "00110010" =>
                  \$v6908\ := \$ram_lock\;
                  if \$v6908\(0) = '1' then
                    state_var7460 := Q_WAIT6907;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET6906;
                  end if;
                when "00110011" =>
                  \$v6911\ := \$ram_lock\;
                  if \$v6911\(0) = '1' then
                    state_var7460 := Q_WAIT6910;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET6909;
                  end if;
                when "00111010" =>
                  \$13926_make_block_n646_id\ := "000000111111";
                  \$13926_make_block_n646_arg\ := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$13911\(48 to 63) & eclat_false & eclat_false & eclat_false & "000"& X"000000" & X"0" & X"000" & X"0" & \$13911\(16 to 47) & \$13911\(120 to 121) & \$13911\(64 to 95) & \$13911\(96 to 103) & \$13911\(104 to 119);
                  state_var7460 := \$13926_MAKE_BLOCK_N646\;
                when "00111100" =>
                  \$v6914\ := \$ram_lock\;
                  if \$v6914\(0) = '1' then
                    state_var7460 := Q_WAIT6913;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET6912;
                  end if;
                when "01000011" =>
                  \$14281\ := work.Assertion.ok(work.Bool.lnot(""&\$13911\(47)));
                  \$v6917\ := \$ram_lock\;
                  if \$v6917\(0) = '1' then
                    state_var7460 := Q_WAIT6916;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$13911\(16 to 46),16), X"000" & X"0"), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6915;
                  end if;
                when "01000100" =>
                  \$14296\ := work.Assertion.ok(work.Bool.lnot(""&\$13911\(47)));
                  \$v6920\ := \$ram_lock\;
                  if \$v6920\(0) = '1' then
                    state_var7460 := Q_WAIT6919;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$13911\(16 to 46),16), X"000" & X"1"), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6918;
                  end if;
                when "01000101" =>
                  \$14311\ := work.Assertion.ok(work.Bool.lnot(""&\$13911\(47)));
                  \$v6923\ := \$ram_lock\;
                  if \$v6923\(0) = '1' then
                    state_var7460 := Q_WAIT6922;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$13911\(16 to 46),16), X"000" & X"2"), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6921;
                  end if;
                when "01000110" =>
                  \$14326\ := work.Assertion.ok(work.Bool.lnot(""&\$13911\(47)));
                  \$v6926\ := \$ram_lock\;
                  if \$v6926\(0) = '1' then
                    state_var7460 := Q_WAIT6925;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$13911\(16 to 46),16), X"000" & X"3"), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6924;
                  end if;
                when "01001001" =>
                  \$v6932\ := \$ram_lock\;
                  if \$v6932\(0) = '1' then
                    state_var7460 := Q_WAIT6931;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13911\(48 to 63), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6930;
                  end if;
                when "01001010" =>
                  \$v6938\ := \$ram_lock\;
                  if \$v6938\(0) = '1' then
                    state_var7460 := Q_WAIT6937;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13911\(48 to 63), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6936;
                  end if;
                when "01001011" =>
                  \$v6944\ := \$ram_lock\;
                  if \$v6944\(0) = '1' then
                    state_var7460 := Q_WAIT6943;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13911\(48 to 63), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6942;
                  end if;
                when "01001100" =>
                  \$v6950\ := \$ram_lock\;
                  if \$v6950\(0) = '1' then
                    state_var7460 := Q_WAIT6949;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13911\(48 to 63), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6948;
                  end if;
                when "01001111" =>
                  \$v6953\ := \$ram_lock\;
                  if \$v6953\(0) = '1' then
                    state_var7460 := Q_WAIT6952;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$13911\(16 to 46),16)));
                    state_var7460 := PAUSE_GET6951;
                  end if;
                when "01010000" =>
                  \$v6959\ := \$ram_lock\;
                  if \$v6959\(0) = '1' then
                    state_var7460 := Q_WAIT6958;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13911\(48 to 63), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6957;
                  end if;
                when "01010001" =>
                  \$v6968\ := \$ram_lock\;
                  if \$v6968\(0) = '1' then
                    state_var7460 := Q_WAIT6967;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13911\(48 to 63), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6966;
                  end if;
                when "01010010" =>
                  \$v6974\ := \$ram_lock\;
                  if \$v6974\(0) = '1' then
                    state_var7460 := Q_WAIT6973;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13911\(48 to 63), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6972;
                  end if;
                when "01010011" =>
                  \$v6983\ := \$ram_lock\;
                  if \$v6983\(0) = '1' then
                    state_var7460 := Q_WAIT6982;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13911\(48 to 63), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6981;
                  end if;
                when "01010101" =>
                  \$13927_branch_if648_id\ := "000001000001";
                  \$13927_branch_if648_arg\ := eclat_false & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  state_var7460 := \$13927_BRANCH_IF648\;
                when "01010110" =>
                  \$13927_branch_if648_id\ := "000001000010";
                  \$13927_branch_if648_arg\ := eclat_true & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  state_var7460 := \$13927_BRANCH_IF648\;
                when "01011000" =>
                  result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & 
                  eclat_if(work.Int.eq(\$13911\(16 to 46), "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when "01011010" =>
                  \$v6986\ := \$ram_lock\;
                  if \$v6986\(0) = '1' then
                    state_var7460 := Q_WAIT6985;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                   \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6984;
                  end if;
                when "01011011" =>
                  \$v6998\ := \$ram_lock\;
                  if \$v6998\(0) = '1' then
                    state_var7460 := Q_WAIT6997;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13911\(104 to 119), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6996;
                  end if;
                when "01100011" =>
                  result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & "000"& X"000000" & X"0" & eclat_true & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when "01100100" =>
                  result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when "01100101" =>
                  result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & "000"& X"000000" & X"2" & eclat_true & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when "01100110" =>
                  result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & "000"& X"000000" & X"3" & eclat_true & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when "01101000" =>
                  \$v7001\ := \$ram_lock\;
                  if \$v7001\(0) = '1' then
                    state_var7460 := Q_WAIT7000;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET6999;
                  end if;
                when "01101001" =>
                  \$v7004\ := \$ram_lock\;
                  if \$v7004\(0) = '1' then
                    state_var7460 := Q_WAIT7003;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET7002;
                  end if;
                when "01101010" =>
                  \$v7007\ := \$ram_lock\;
                  if \$v7007\(0) = '1' then
                    state_var7460 := Q_WAIT7006;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET7005;
                  end if;
                when "01101011" =>
                  \$v7010\ := \$ram_lock\;
                  if \$v7010\(0) = '1' then
                    state_var7460 := Q_WAIT7009;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                    \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET7008;
                  end if;
                when "01101110" =>
                  \$14564_binop_int6435900_id\ := "000001000111";
                  \$14564_binop_int6435900_arg\ := X"0000000" & X"0" & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  state_var7460 := \$14564_BINOP_INT6435900\;
                when "01101111" =>
                  \$14644_binop_int6435901_id\ := "000001001100";
                  \$14644_binop_int6435901_arg\ := X"0000000" & X"1" & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  state_var7460 := \$14644_BINOP_INT6435901\;
                when "01110000" =>
                  \$14724_binop_int6435902_id\ := "000001010001";
                  \$14724_binop_int6435902_arg\ := X"0000000" & X"2" & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  state_var7460 := \$14724_BINOP_INT6435902\;
                when "01110001" =>
                  \$14804_binop_int6435903_id\ := "000001010110";
                  \$14804_binop_int6435903_arg\ := X"0000000" & X"3" & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  state_var7460 := \$14804_BINOP_INT6435903\;
                when "01110010" =>
                  \$14884_binop_int6435904_id\ := "000001011011";
                  \$14884_binop_int6435904_arg\ := X"0000000" & X"4" & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  state_var7460 := \$14884_BINOP_INT6435904\;
                when "01110011" =>
                  \$14964_binop_int6435905_id\ := "000001100000";
                  \$14964_binop_int6435905_arg\ := X"0000000" & X"5" & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  state_var7460 := \$14964_BINOP_INT6435905\;
                when "01110100" =>
                  \$15044_binop_int6435906_id\ := "000001100101";
                  \$15044_binop_int6435906_arg\ := X"0000000" & X"6" & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  state_var7460 := \$15044_BINOP_INT6435906\;
                when "01110101" =>
                  \$15124_binop_int6435907_id\ := "000001101010";
                  \$15124_binop_int6435907_arg\ := X"0000000" & X"7" & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  state_var7460 := \$15124_BINOP_INT6435907\;
                when "01110110" =>
                  \$15204_binop_int6435908_id\ := "000001101111";
                  \$15204_binop_int6435908_arg\ := X"0000000" & X"8" & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  state_var7460 := \$15204_BINOP_INT6435908\;
                when "01110111" =>
                  \$15284_binop_int6435909_id\ := "000001110100";
                  \$15284_binop_int6435909_arg\ := X"0000000" & X"9" & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  state_var7460 := \$15284_BINOP_INT6435909\;
                when "01111000" =>
                  \$15364_binop_int6435910_id\ := "000001111001";
                  \$15364_binop_int6435910_arg\ := X"0000000" & X"a" & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  state_var7460 := \$15364_BINOP_INT6435910\;
                when "10000010" =>
                  \$15444\ := work.Print.print_string(clk,of_string("fatal error: "));
                  \$15445\ := work.Print.print_string(clk,of_string("unsupported instruction GETMETHOD"));
                  \$15446\ := work.Print.print_newline(clk,eclat_unit);
                  \$15447_forever6705911_id\ := "000001111010";
                  \$15447_forever6705911_arg\ := eclat_unit;
                  state_var7460 := \$15447_FOREVER6705911\;
                when "10001001" =>
                  \$15451_binop_int6435912_id\ := "000001111111";
                  \$15451_binop_int6435912_arg\ := X"0000000" & X"b" & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  state_var7460 := \$15451_BINOP_INT6435912\;
                when "10001010" =>
                  \$15531_binop_int6435913_id\ := "000010000100";
                  \$15531_binop_int6435913_arg\ := X"0000000" & X"c" & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  state_var7460 := \$15531_BINOP_INT6435913\;
                when "10001101" =>
                  \$15611\ := work.Print.print_string(clk,of_string("fatal error: "));
                  \$15612\ := work.Print.print_string(clk,of_string("unsupported instruction GETPUBMET"));
                  \$15613\ := work.Print.print_newline(clk,eclat_unit);
                  \$15614_forever6705914_id\ := "000010000101";
                  \$15614_forever6705914_arg\ := eclat_unit;
                  state_var7460 := \$15614_FOREVER6705914\;
                when "10001110" =>
                  \$15618\ := work.Print.print_string(clk,of_string("fatal error: "));
                  \$15619\ := work.Print.print_string(clk,of_string("unsupported instruction GETDYNMET"));
                  \$15620\ := work.Print.print_newline(clk,eclat_unit);
                  \$15621_forever6705915_id\ := "000010000110";
                  \$15621_forever6705915_arg\ := eclat_unit;
                  state_var7460 := \$15621_FOREVER6705915\;
                when "01111001" =>
                  \$15625_binop_compare6455916_id\ := "000010001000";
                  \$15625_binop_compare6455916_arg\ := X"0000000" & X"0" & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  state_var7460 := \$15625_BINOP_COMPARE6455916\;
                when "01111010" =>
                  \$15661_binop_compare6455917_id\ := "000010001010";
                  \$15661_binop_compare6455917_arg\ := X"0000000" & X"1" & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  state_var7460 := \$15661_BINOP_COMPARE6455917\;
                when "01111011" =>
                  \$15697_binop_compare6455918_id\ := "000010001100";
                  \$15697_binop_compare6455918_arg\ := X"0000000" & X"2" & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  state_var7460 := \$15697_BINOP_COMPARE6455918\;
                when "01111100" =>
                  \$15733_binop_compare6455919_id\ := "000010001110";
                  \$15733_binop_compare6455919_arg\ := X"0000000" & X"3" & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  state_var7460 := \$15733_BINOP_COMPARE6455919\;
                when "01111101" =>
                  \$15769_binop_compare6455920_id\ := "000010010000";
                  \$15769_binop_compare6455920_arg\ := X"0000000" & X"4" & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  state_var7460 := \$15769_BINOP_COMPARE6455920\;
                when "01111110" =>
                  \$15805_binop_compare6455921_id\ := "000010010010";
                  \$15805_binop_compare6455921_arg\ := X"0000000" & X"5" & \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  state_var7460 := \$15805_BINOP_COMPARE6455921\;
                when "10000001" =>
                  result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & 
                  eclat_if(""&\$13911\(47) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when "10001111" =>
                  \$15847\ := work.Print.print_string(clk,of_string("STOP : "));
                  result6468 := \$13911\(0 to 15) & \$13911\(16 to 47) & \$13911\(48 to 63) & \$13911\(64 to 119) & eclat_true & ""&\$13911\(121);
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                when others =>
                  \$v7449\ := \$code_lock\;
                  if \$v7449\(0) = '1' then
                    state_var7460 := Q_WAIT7448;
                  else
                    acquire(\$code_lock\);
                    \$code_ptr\ <= to_integer(unsigned(work.Int.add(\$13911\(0 to 15), X"000" & X"1")));
                    state_var7460 := PAUSE_GET7447;
                  end if;
                end case;
              when PAUSE_SET6471 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18546\ := eclat_unit;
                \$13920_loop666_arg\ := work.Int.add(\$13920_loop666_arg\(0 to 15), X"000" & X"1") & \$13920_loop666_arg\(16 to 31) & \$13920_loop666_arg\(32 to 47) & \$13920_loop666_arg\(48 to 63);
                state_var7460 := \$13920_LOOP666\;
              when PAUSE_SET6478 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18450\ := eclat_unit;
                \$13921_loop665_arg\ := work.Int.add(\$13921_loop665_arg\(0 to 15), X"000" & X"1") & \$18447\(32 to 47) & \$13921_loop665_arg\(32 to 47) & \$13921_loop665_arg\(48 to 63) & \$13921_loop665_arg\(64 to 79) & \$13921_loop665_arg\(80 to 95);
                state_var7460 := \$13921_LOOP665\;
              when PAUSE_SET6481 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18480\ := eclat_unit;
                \$18447\ := eclat_resize(\$13921_loop665_arg\(16 to 31),31) & eclat_false & 
                work.Int.add(\$13921_loop665_arg\(16 to 31), work.Int.add(
                                                             eclat_resize(
                                                             work.Int.lsr(
                                                             \$18464_hd\(0 to 30), X"0000000" & X"2"),16), X"000" & X"1"));
                \$v6480\ := \$ram_lock\;
                if \$v6480\(0) = '1' then
                  state_var7460 := Q_WAIT6479;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$13921_loop665_arg\(64 to 79), \$13921_loop665_arg\(0 to 15))));
                  \$ram_write\ <= \$18447\(0 to 31); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6478;
                end if;
              when PAUSE_SET6484 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18479\ := eclat_unit;
                \$v6483\ := \$ram_lock\;
                if \$v6483\(0) = '1' then
                  state_var7460 := Q_WAIT6482;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$18443\(0 to 30),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$13921_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6481;
                end if;
              when PAUSE_SET6487 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$18477\ := eclat_unit;
                \$13920_loop666_id\ := "000000100000";
                \$13920_loop666_arg\ := X"000" & X"1" & \$13921_loop665_arg\(16 to 31) & eclat_resize(\$18443\(0 to 30),16) & eclat_resize(
                work.Int.lsr(\$18464_hd\(0 to 30), X"0000000" & X"2"),16);
                state_var7460 := \$13920_LOOP666\;
              when PAUSE_SET6712 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$17396\ := eclat_unit;
                \$13923_make_block579_result\ := \$17389\(0 to 31) & \$17389\(32 to 63) & eclat_resize(\$17389\(64 to 79),31) & eclat_false;
                case \$13923_make_block579_id\ is
                when "000000110100" =>
                  \$17232\ := \$13923_make_block579_result\;
                  \$v6770\ := ""&\$13926_make_block_n646_arg\(32);
                  if \$v6770\(0) = '1' then
                    \$v6769\ := \$ram_lock\;
                    if \$v6769\(0) = '1' then
                      state_var7460 := Q_WAIT6768;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                              work.Int.add(
                                                              eclat_resize(\$17232\(64 to 94),16), X"000" & X"0"), X"000" & X"1")));
                      \$ram_write\ <= \$17232\(0 to 31); \$ram_write_request\ <= '1';
                      state_var7460 := PAUSE_SET6767;
                    end if;
                  else
                    \$17236\ := eclat_unit;
                    \$v6766\ := ""&\$13926_make_block_n646_arg\(33);
                    if \$v6766\(0) = '1' then
                      \$v6765\ := \$ram_lock\;
                      if \$v6765\(0) = '1' then
                        state_var7460 := Q_WAIT6764;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(
                                                          \$13926_make_block_n646_arg\(16 to 31), X"000" & X"1")));
                        state_var7460 := PAUSE_GET6763;
                      end if;
                    else
                      \$17237_sp\ := \$13926_make_block_n646_arg\(16 to 31);
                      \$v6759\ := ""&\$13926_make_block_n646_arg\(34);
                      if \$v6759\(0) = '1' then
                        \$v6758\ := \$ram_lock\;
                        if \$v6758\(0) = '1' then
                          state_var7460 := Q_WAIT6757;
                        else
                          acquire(\$ram_lock\);
                          \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(
                                                            \$17237_sp\, X"000" & X"1")));
                          state_var7460 := PAUSE_GET6756;
                        end if;
                      else
                        \$17238_sp\ := \$17237_sp\;
                        \$13926_make_block_n646_result\ := \$13926_make_block_n646_arg\(0 to 15) & \$17232\(64 to 95) & \$17238_sp\ & \$17232\(32 to 63) & \$13926_make_block_n646_arg\(148 to 155) & \$13926_make_block_n646_arg\(156 to 171) & \$13926_make_block_n646_arg\(114 to 115);
                        result6468 := \$13926_make_block_n646_result\;
                        rdy6469 := eclat_true;
                        state_var7460 := IDLE6470;
                      end if;
                    end if;
                  end if;
                when "000010010111" =>
                  \$16024\ := \$13923_make_block579_result\;
                  \$v7232\ := \$ram_lock\;
                  if \$v7232\(0) = '1' then
                    state_var7460 := Q_WAIT7231;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            work.Int.add(
                                                            eclat_resize(\$16024\(64 to 94),16), X"000" & X"0"), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(work.Int.sub(work.Int.add(
                                                              \$13911\(0 to 15), X"000" & X"2"), X"000" & X"3"),31) & eclat_true; \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET7230;
                  end if;
                when "000010101000" =>
                  \$16651\ := \$13923_make_block579_result\;
                  \$v7368\ := \$ram_lock\;
                  if \$v7368\(0) = '1' then
                    state_var7460 := Q_WAIT7367;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            work.Int.add(
                                                            eclat_resize(\$16651\(64 to 94),16), X"000" & X"0"), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(work.Int.add(work.Int.add(
                                                              \$13911\(0 to 15), X"000" & X"2"), eclat_resize(\$16624_argument2\,16)),31) & eclat_true; \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET7366;
                  end if;
                when "000010101010" =>
                  \$16741\ := \$13923_make_block579_result\;
                  \$v7397\ := \$ram_lock\;
                  if \$v7397\(0) = '1' then
                    state_var7460 := Q_WAIT7396;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            work.Int.add(
                                                            eclat_resize(\$16741\(64 to 94),16), X"000" & X"0"), X"000" & X"1")));
                    \$ram_write\ <= \$16741\(0 to 31); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET7395;
                  end if;
                when "000010111010" =>
                  \$17001\ := \$13923_make_block579_result\;
                  \$v7430\ := \$ram_lock\;
                  if \$v7430\(0) = '1' then
                    state_var7460 := Q_WAIT7429;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                            work.Int.add(
                                                            eclat_resize(\$17001\(64 to 94),16), X"000" & X"0"), X"000" & X"1")));
                    \$ram_write\ <= eclat_resize(work.Int.add(work.Int.add(
                                                              \$13911\(0 to 15), X"000" & X"3"), eclat_resize(\$16998_argument3\,16)),31) & eclat_true; \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET7428;
                  end if;
                when others =>
                  
                end case;
              when PAUSE_SET6718 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$17347\ := eclat_unit;
                \$17333_sp\ := work.Int.add(\$17332_sp\, X"000" & X"1");
                \$v6717\ := \$ram_lock\;
                if \$v6717\(0) = '1' then
                  state_var7460 := Q_WAIT6716;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13924_apply638_arg\(60 to 90),16), X"000" & X"0"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6715;
                end if;
              when PAUSE_SET6722 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$17348\ := eclat_unit;
                \$17332_sp\ := work.Int.add(\$17331_sp\, X"000" & X"1");
                \$v6721\ := ""&\$13924_apply638_arg\(0);
                if \$v6721\(0) = '1' then
                  \$v6720\ := \$ram_lock\;
                  if \$v6720\(0) = '1' then
                    state_var7460 := Q_WAIT6719;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17332_sp\));
                    \$ram_write\ <= \$17321\(0 to 31); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET6718;
                  end if;
                else
                  \$17333_sp\ := \$17332_sp\;
                  \$v6717\ := \$ram_lock\;
                  if \$v6717\(0) = '1' then
                    state_var7460 := Q_WAIT6716;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                   eclat_resize(\$13924_apply638_arg\(60 to 90),16), X"000" & X"0"), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6715;
                  end if;
                end if;
              when PAUSE_SET6726 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$17349\ := eclat_unit;
                \$17331_sp\ := work.Int.add(\$17330_sp\, X"000" & X"1");
                \$v6725\ := ""&\$13924_apply638_arg\(1);
                if \$v6725\(0) = '1' then
                  \$v6724\ := \$ram_lock\;
                  if \$v6724\(0) = '1' then
                    state_var7460 := Q_WAIT6723;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17331_sp\));
                    \$ram_write\ <= \$17324\(0 to 31); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET6722;
                  end if;
                else
                  \$17332_sp\ := \$17331_sp\;
                  \$v6721\ := ""&\$13924_apply638_arg\(0);
                  if \$v6721\(0) = '1' then
                    \$v6720\ := \$ram_lock\;
                    if \$v6720\(0) = '1' then
                      state_var7460 := Q_WAIT6719;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(\$17332_sp\));
                      \$ram_write\ <= \$17321\(0 to 31); \$ram_write_request\ <= '1';
                      state_var7460 := PAUSE_SET6718;
                    end if;
                  else
                    \$17333_sp\ := \$17332_sp\;
                    \$v6717\ := \$ram_lock\;
                    if \$v6717\(0) = '1' then
                      state_var7460 := Q_WAIT6716;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                        work.Int.add(
                                                        eclat_resize(\$13924_apply638_arg\(60 to 90),16), X"000" & X"0"), X"000" & X"1")));
                      state_var7460 := PAUSE_GET6715;
                    end if;
                  end if;
                end if;
              when PAUSE_SET6730 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$17354\ := eclat_unit;
                \$17330_sp\ := work.Int.add(work.Int.add(work.Int.add(
                                                         \$17327\(32 to 47), X"000" & X"1"), X"000" & X"1"), X"000" & X"1");
                \$v6729\ := ""&\$13924_apply638_arg\(2);
                if \$v6729\(0) = '1' then
                  \$v6728\ := \$ram_lock\;
                  if \$v6728\(0) = '1' then
                    state_var7460 := Q_WAIT6727;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$17330_sp\));
                    \$ram_write\ <= \$17327\(0 to 31); \$ram_write_request\ <= '1';
                    state_var7460 := PAUSE_SET6726;
                  end if;
                else
                  \$17331_sp\ := \$17330_sp\;
                  \$v6725\ := ""&\$13924_apply638_arg\(1);
                  if \$v6725\(0) = '1' then
                    \$v6724\ := \$ram_lock\;
                    if \$v6724\(0) = '1' then
                      state_var7460 := Q_WAIT6723;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr_write\ <= to_integer(unsigned(\$17331_sp\));
                      \$ram_write\ <= \$17324\(0 to 31); \$ram_write_request\ <= '1';
                      state_var7460 := PAUSE_SET6722;
                    end if;
                  else
                    \$17332_sp\ := \$17331_sp\;
                    \$v6721\ := ""&\$13924_apply638_arg\(0);
                    if \$v6721\(0) = '1' then
                      \$v6720\ := \$ram_lock\;
                      if \$v6720\(0) = '1' then
                        state_var7460 := Q_WAIT6719;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr_write\ <= to_integer(unsigned(\$17332_sp\));
                        \$ram_write\ <= \$17321\(0 to 31); \$ram_write_request\ <= '1';
                        state_var7460 := PAUSE_SET6718;
                      end if;
                    else
                      \$17333_sp\ := \$17332_sp\;
                      \$v6717\ := \$ram_lock\;
                      if \$v6717\(0) = '1' then
                        state_var7460 := Q_WAIT6716;
                      else
                        acquire(\$ram_lock\);
                        \$ram_ptr\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$13924_apply638_arg\(60 to 90),16), X"000" & X"0"), X"000" & X"1")));
                        state_var7460 := PAUSE_GET6715;
                      end if;
                    end if;
                  end if;
                end if;
              when PAUSE_SET6733 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$17353\ := eclat_unit;
                \$v6732\ := \$ram_lock\;
                if \$v6732\(0) = '1' then
                  state_var7460 := Q_WAIT6731;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          \$17327\(32 to 47), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(work.Int.add(\$13924_apply638_arg\(44 to 59), X"000" & X"1"),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6730;
                end if;
              when PAUSE_SET6736 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$17352\ := eclat_unit;
                \$v6735\ := \$ram_lock\;
                if \$v6735\(0) = '1' then
                  state_var7460 := Q_WAIT6734;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$17327\(32 to 47), X"000" & X"1")));
                  \$ram_write\ <= \$13924_apply638_arg\(110 to 141); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6733;
                end if;
              when PAUSE_SET6753 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$17243\ := eclat_unit;
                \$17238_sp\ := work.Int.sub(\$17237_sp\, X"000" & X"1");
                \$13926_make_block_n646_result\ := \$13926_make_block_n646_arg\(0 to 15) & \$17232\(64 to 95) & \$17238_sp\ & \$17232\(32 to 63) & \$13926_make_block_n646_arg\(148 to 155) & \$13926_make_block_n646_arg\(156 to 171) & \$13926_make_block_n646_arg\(114 to 115);
                result6468 := \$13926_make_block_n646_result\;
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_SET6760 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$17254\ := eclat_unit;
                \$17237_sp\ := work.Int.sub(\$13926_make_block_n646_arg\(16 to 31), X"000" & X"1");
                \$v6759\ := ""&\$13926_make_block_n646_arg\(34);
                if \$v6759\(0) = '1' then
                  \$v6758\ := \$ram_lock\;
                  if \$v6758\(0) = '1' then
                    state_var7460 := Q_WAIT6757;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$17237_sp\, X"000" & X"1")));
                    state_var7460 := PAUSE_GET6756;
                  end if;
                else
                  \$17238_sp\ := \$17237_sp\;
                  \$13926_make_block_n646_result\ := \$13926_make_block_n646_arg\(0 to 15) & \$17232\(64 to 95) & \$17238_sp\ & \$17232\(32 to 63) & \$13926_make_block_n646_arg\(148 to 155) & \$13926_make_block_n646_arg\(156 to 171) & \$13926_make_block_n646_arg\(114 to 115);
                  result6468 := \$13926_make_block_n646_result\;
                  rdy6469 := eclat_true;
                  state_var7460 := IDLE6470;
                end if;
              when PAUSE_SET6767 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$17236\ := eclat_unit;
                \$v6766\ := ""&\$13926_make_block_n646_arg\(33);
                if \$v6766\(0) = '1' then
                  \$v6765\ := \$ram_lock\;
                  if \$v6765\(0) = '1' then
                    state_var7460 := Q_WAIT6764;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13926_make_block_n646_arg\(16 to 31), X"000" & X"1")));
                    state_var7460 := PAUSE_GET6763;
                  end if;
                else
                  \$17237_sp\ := \$13926_make_block_n646_arg\(16 to 31);
                  \$v6759\ := ""&\$13926_make_block_n646_arg\(34);
                  if \$v6759\(0) = '1' then
                    \$v6758\ := \$ram_lock\;
                    if \$v6758\(0) = '1' then
                      state_var7460 := Q_WAIT6757;
                    else
                      acquire(\$ram_lock\);
                      \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(
                                                        \$17237_sp\, X"000" & X"1")));
                      state_var7460 := PAUSE_GET6756;
                    end if;
                  else
                    \$17238_sp\ := \$17237_sp\;
                    \$13926_make_block_n646_result\ := \$13926_make_block_n646_arg\(0 to 15) & \$17232\(64 to 95) & \$17238_sp\ & \$17232\(32 to 63) & \$13926_make_block_n646_arg\(148 to 155) & \$13926_make_block_n646_arg\(156 to 171) & \$13926_make_block_n646_arg\(114 to 115);
                    result6468 := \$13926_make_block_n646_result\;
                    rdy6469 := eclat_true;
                    state_var7460 := IDLE6470;
                  end if;
                end if;
              when PAUSE_SET6775 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$17184\ := eclat_unit;
                \$13928_w652_arg\ := work.Int.add(\$13928_w652_arg\(0 to 15), X"000" & X"1") & \$13928_w652_arg\(16 to 31) & \$13928_w652_arg\(32 to 47) & \$13928_w652_arg\(48 to 63);
                state_var7460 := \$13928_W652\;
              when PAUSE_SET6806 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$14008\ := eclat_unit;
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$13911\(16 to 47) & 
                work.Int.add(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_SET6809 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$14012\ := eclat_unit;
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & \$13911\(16 to 47) & 
                work.Int.add(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_SET6815 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$14015\ := eclat_unit;
                \$v6814\ := \$ram_lock\;
                if \$v6814\(0) = '1' then
                  state_var7460 := Q_WAIT6813;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6812;
                end if;
              when PAUSE_SET6821 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$14024\ := eclat_unit;
                \$v6820\ := \$ram_lock\;
                if \$v6820\(0) = '1' then
                  state_var7460 := Q_WAIT6819;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"2"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6818;
                end if;
              when PAUSE_SET6827 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$14033\ := eclat_unit;
                \$v6826\ := \$ram_lock\;
                if \$v6826\(0) = '1' then
                  state_var7460 := Q_WAIT6825;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"3"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6824;
                end if;
              when PAUSE_SET6833 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$14042\ := eclat_unit;
                \$v6832\ := \$ram_lock\;
                if \$v6832\(0) = '1' then
                  state_var7460 := Q_WAIT6831;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"4"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6830;
                end if;
              when PAUSE_SET6839 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$14051\ := eclat_unit;
                \$v6838\ := \$ram_lock\;
                if \$v6838\(0) = '1' then
                  state_var7460 := Q_WAIT6837;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"5"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6836;
                end if;
              when PAUSE_SET6845 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$14060\ := eclat_unit;
                \$v6844\ := \$ram_lock\;
                if \$v6844\(0) = '1' then
                  state_var7460 := Q_WAIT6843;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"6"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6842;
                end if;
              when PAUSE_SET6851 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$14069\ := eclat_unit;
                \$v6850\ := \$ram_lock\;
                if \$v6850\(0) = '1' then
                  state_var7460 := Q_WAIT6849;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"7"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6848;
                end if;
              when PAUSE_SET6869 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$14122\ := eclat_unit;
                \$v6868\ := \$ram_lock\;
                if \$v6868\(0) = '1' then
                  state_var7460 := Q_WAIT6867;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13911\(64 to 94),16), 
                                                                 work.Int.sub(
                                                                 X"000" & X"1", X"000" & X"1")), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6866;
                end if;
              when PAUSE_SET6875 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$14135\ := eclat_unit;
                \$v6874\ := \$ram_lock\;
                if \$v6874\(0) = '1' then
                  state_var7460 := Q_WAIT6873;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13911\(64 to 94),16), 
                                                                 work.Int.sub(
                                                                 X"000" & X"2", X"000" & X"1")), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6872;
                end if;
              when PAUSE_SET6881 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$14148\ := eclat_unit;
                \$v6880\ := \$ram_lock\;
                if \$v6880\(0) = '1' then
                  state_var7460 := Q_WAIT6879;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13911\(64 to 94),16), 
                                                                 work.Int.sub(
                                                                 X"000" & X"3", X"000" & X"1")), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6878;
                end if;
              when PAUSE_SET6887 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$14161\ := eclat_unit;
                \$v6886\ := \$ram_lock\;
                if \$v6886\(0) = '1' then
                  state_var7460 := Q_WAIT6885;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13911\(64 to 94),16), 
                                                                 work.Int.sub(
                                                                 X"000" & X"4", X"000" & X"1")), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6884;
                end if;
              when PAUSE_SET6893 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$14222\ := eclat_unit;
                \$14207_loop_push6495899_arg\ := work.Int.add(\$14207_loop_push6495899_arg\(0 to 15), X"000" & X"1") & 
                work.Int.add(\$14207_loop_push6495899_arg\(16 to 23), "00000001") & \$14207_loop_push6495899_arg\(24 to 55) & \$14207_loop_push6495899_arg\(56 to 63);
                state_var7460 := \$14207_LOOP_PUSH6495899\;
              when PAUSE_SET6903 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$14254\ := eclat_unit;
                \$13925_offsetclosure_n639_id\ := "000000111100";
                \$13925_offsetclosure_n639_arg\ := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & 
                work.Int.add(\$13911\(48 to 63), X"000" & X"1") & work.Int.neg(
                                                                  X"000" & X"2") & \$13911\(64 to 119) & \$13911\(120 to 121) & \$13911\(64 to 95);
                state_var7460 := \$13925_OFFSETCLOSURE_N639\;
              when PAUSE_SET6906 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$14260\ := eclat_unit;
                \$13925_offsetclosure_n639_id\ := "000000111101";
                \$13925_offsetclosure_n639_arg\ := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & 
                work.Int.add(\$13911\(48 to 63), X"000" & X"1") & X"000" & X"0" & \$13911\(64 to 119) & \$13911\(120 to 121) & \$13911\(64 to 95);
                state_var7460 := \$13925_OFFSETCLOSURE_N639\;
              when PAUSE_SET6909 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$14265\ := eclat_unit;
                \$13925_offsetclosure_n639_id\ := "000000111110";
                \$13925_offsetclosure_n639_arg\ := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & 
                work.Int.add(\$13911\(48 to 63), X"000" & X"1") & X"000" & X"2" & \$13911\(64 to 119) & \$13911\(120 to 121) & \$13911\(64 to 95);
                state_var7460 := \$13925_OFFSETCLOSURE_N639\;
              when PAUSE_SET6912 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$14273\ := eclat_unit;
                \$13926_make_block_n646_id\ := "000001000000";
                \$13926_make_block_n646_arg\ := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & 
                work.Int.add(\$13911\(48 to 63), X"000" & X"1") & eclat_false & eclat_false & eclat_false & "000"& X"000000" & X"0" & X"000" & X"0" & \$13911\(16 to 47) & \$13911\(120 to 121) & \$13911\(64 to 95) & \$13911\(96 to 103) & \$13911\(104 to 119);
                state_var7460 := \$13926_MAKE_BLOCK_N646\;
              when PAUSE_SET6927 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$14342\ := eclat_unit;
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & 
                work.Int.sub(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_SET6933 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$14355\ := eclat_unit;
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & 
                work.Int.sub(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_SET6939 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$14368\ := eclat_unit;
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & 
                work.Int.sub(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_SET6945 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$14381\ := eclat_unit;
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & 
                work.Int.sub(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_SET6960 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$14431\ := eclat_unit;
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & 
                work.Int.sub(work.Int.sub(\$13911\(48 to 63), X"000" & X"1"), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_SET6975 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$14471\ := eclat_unit;
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & 
                work.Int.sub(work.Int.sub(\$13911\(48 to 63), X"000" & X"1"), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_SET6999 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$14552\ := eclat_unit;
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & "000"& X"000000" & X"0" & eclat_true & 
                work.Int.add(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_SET7002 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$14555\ := eclat_unit;
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & 
                work.Int.add(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_SET7005 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$14558\ := eclat_unit;
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & "000"& X"000000" & X"2" & eclat_true & 
                work.Int.add(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_SET7008 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$14561\ := eclat_unit;
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"1") & "000"& X"000000" & X"3" & eclat_true & 
                work.Int.add(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_SET7171 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$15860\ := eclat_unit;
                \$v7170\ := \$ram_lock\;
                if \$v7170\(0) = '1' then
                  state_var7460 := Q_WAIT7169;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$13911\(48 to 63), X"000" & X"1"), eclat_resize(\$15851_argument1\,16)), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7168;
                end if;
              when PAUSE_SET7174 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$15874\ := eclat_unit;
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"2") & "000"& X"000000" & X"1" & eclat_true & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_SET7183 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$15893\ := eclat_unit;
                \$v7182\ := \$ram_lock\;
                if \$v7182\(0) = '1' then
                  state_var7460 := Q_WAIT7181;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13911\(64 to 94),16), 
                                                                 work.Int.sub(
                                                                 eclat_resize(\$15851_argument1\,16), X"000" & X"1")), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7180;
                end if;
              when PAUSE_SET7186 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$15910\ := eclat_unit;
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"2") & \$13911\(16 to 47) & 
                work.Int.add(work.Int.add(work.Int.add(\$13911\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_SET7189 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$15909\ := eclat_unit;
                \$v7188\ := \$ram_lock\;
                if \$v7188\(0) = '1' then
                  state_var7460 := Q_WAIT7187;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(work.Int.add(work.Int.add(
                                                            \$13911\(0 to 15), X"000" & X"1"), eclat_resize(\$15851_argument1\,16)),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7186;
                end if;
              when PAUSE_SET7192 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$15908\ := eclat_unit;
                \$v7191\ := \$ram_lock\;
                if \$v7191\(0) = '1' then
                  state_var7460 := Q_WAIT7190;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$13911\(48 to 63), X"000" & X"1")));
                  \$ram_write\ <= \$13911\(64 to 95); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7189;
                end if;
              when PAUSE_SET7220 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$16078\ := eclat_unit;
                \$16063_w6515922_arg\ := work.Int.add(\$16063_w6515922_arg\(0 to 7), "00000001") & 
                work.Int.sub(\$16063_w6515922_arg\(8 to 23), X"000" & X"1") & \$16063_w6515922_arg\(24 to 31) & \$16063_w6515922_arg\(32 to 63);
                state_var7460 := \$16063_W6515922\;
              when PAUSE_SET7227 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$16035\ := eclat_unit;
                \$16063_w6515922_id\ := "000010010110";
                \$16063_w6515922_arg\ := "00000000" & \$13911\(48 to 63) & \$13911\(96 to 103) & \$16024\(64 to 95);
                state_var7460 := \$16063_W6515922\;
              when PAUSE_SET7230 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$16031\ := eclat_unit;
                \$v7229\ := \$ram_lock\;
                if \$v7229\(0) = '1' then
                  state_var7460 := Q_WAIT7228;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$16024\(64 to 94),16), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= \$16024\(32 to 63); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7227;
                end if;
              when PAUSE_SET7234 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$16115\ := eclat_unit;
                \$13925_offsetclosure_n639_id\ := "000010011001";
                \$13925_offsetclosure_n639_arg\ := work.Int.add(\$13911\(0 to 15), X"000" & X"2") & 
                work.Int.add(\$13911\(48 to 63), X"000" & X"1") & eclat_resize(\$15851_argument1\,16) & \$13911\(64 to 119) & \$13911\(120 to 121) & \$13911\(64 to 95);
                state_var7460 := \$13925_OFFSETCLOSURE_N639\;
              when PAUSE_SET7243 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$16126\ := eclat_unit;
                \$v7242\ := \$ram_lock\;
                if \$v7242\(0) = '1' then
                  state_var7460 := Q_WAIT7241;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(X"3e80", eclat_resize(\$15851_argument1\,16))));
                  state_var7460 := PAUSE_GET7240;
                end if;
              when PAUSE_SET7246 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$16133\ := eclat_unit;
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"2") & "000"& X"000000" & X"1" & eclat_true & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_SET7249 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$16141\ := eclat_unit;
                \$13926_make_block_n646_id\ := "000010011011";
                \$13926_make_block_n646_arg\ := work.Int.add(\$13911\(0 to 15), X"000" & X"2") & 
                work.Int.add(\$13911\(48 to 63), X"000" & X"1") & eclat_false & eclat_false & eclat_false & \$15851_argument1\ & X"000" & X"0" & \$13911\(16 to 47) & \$13911\(120 to 121) & \$13911\(64 to 95) & \$13911\(96 to 103) & \$13911\(104 to 119);
                state_var7460 := \$13926_MAKE_BLOCK_N646\;
              when PAUSE_SET7255 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$16182\ := eclat_unit;
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"2") & "000"& X"000000" & X"1" & eclat_true & 
                work.Int.sub(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_SET7268 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$16234\ := eclat_unit;
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"2") & \$13911\(16 to 47) & 
                work.Int.add(work.Int.add(work.Int.add(work.Int.add(\$13911\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1"), X"000" & X"1") & \$13911\(64 to 95) & \$13911\(96 to 103) & 
                work.Int.add(work.Int.add(work.Int.add(work.Int.add(\$13911\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1"), X"000" & X"1") & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_SET7271 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$16233\ := eclat_unit;
                \$v7270\ := \$ram_lock\;
                if \$v7270\(0) = '1' then
                  state_var7460 := Q_WAIT7269;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          work.Int.add(
                                                          \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(work.Int.add(work.Int.add(
                                                            \$13911\(0 to 15), X"000" & X"1"), eclat_resize(\$15851_argument1\,16)),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7268;
                end if;
              when PAUSE_SET7274 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$16232\ := eclat_unit;
                \$v7273\ := \$ram_lock\;
                if \$v7273\(0) = '1' then
                  state_var7460 := Q_WAIT7272;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$13911\(104 to 119),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7271;
                end if;
              when PAUSE_SET7277 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$16231\ := eclat_unit;
                \$v7276\ := \$ram_lock\;
                if \$v7276\(0) = '1' then
                  state_var7460 := Q_WAIT7275;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$13911\(48 to 63), X"000" & X"1")));
                  \$ram_write\ <= \$13911\(64 to 95); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7274;
                end if;
              when PAUSE_SET7284 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$16271\ := eclat_unit;
                \$v7283\ := \$15851_argument1\;
                case \$v7283\ is
                when "000"& X"000000" & X"0" =>
                  \$16288\ := work.Print.print_string(clk,of_string("======> "));
                  \$16292\ := work.Int.print(clk,\$13911\(16 to 46));
                  \$16293\ := work.Print.print_newline(clk,eclat_unit);
                  \$16272\ := "000"& X"000000" & X"1" & eclat_true & \$13911\(0 to 15) & \$13911\(16 to 47) & 
                  work.Int.add(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 95) & \$13911\(96 to 103) & \$13911\(104 to 119) & \$13911\(120 to 121);
                  \$v7282\ := \$ram_lock\;
                  if \$v7282\(0) = '1' then
                    state_var7460 := Q_WAIT7281;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$16272\(80 to 95), X"000" & X"1")));
                    state_var7460 := PAUSE_GET7280;
                  end if;
                when others =>
                  \$16296\ := work.Print.print_string(clk,of_string("unknown primitive"));
                  \$16272\ := "000"& X"000000" & X"1" & eclat_true & \$13911\(0 to 15) & \$13911\(16 to 47) & 
                  work.Int.add(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 95) & \$13911\(96 to 103) & \$13911\(104 to 119) & \$13911\(120 to 121);
                  \$v7282\ := \$ram_lock\;
                  if \$v7282\(0) = '1' then
                    state_var7460 := Q_WAIT7281;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$16272\(80 to 95), X"000" & X"1")));
                    state_var7460 := PAUSE_GET7280;
                  end if;
                end case;
              when PAUSE_SET7291 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$16300\ := eclat_unit;
                \$v7290\ := \$15851_argument1\;
                case \$v7290\ is
                when "000"& X"000000" & X"0" =>
                  \$16317\ := work.Print.print_string(clk,of_string("======> "));
                  \$16321\ := work.Int.print(clk,\$13911\(16 to 46));
                  \$16322\ := work.Print.print_newline(clk,eclat_unit);
                  \$16301\ := "000"& X"000000" & X"1" & eclat_true & \$13911\(0 to 15) & \$13911\(16 to 47) & 
                  work.Int.add(work.Int.sub(\$13911\(48 to 63), X"000" & X"1"), X"000" & X"1") & \$13911\(64 to 95) & \$13911\(96 to 103) & \$13911\(104 to 119) & \$13911\(120 to 121);
                  \$v7289\ := \$ram_lock\;
                  if \$v7289\(0) = '1' then
                    state_var7460 := Q_WAIT7288;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$16301\(80 to 95), X"000" & X"1")));
                    state_var7460 := PAUSE_GET7287;
                  end if;
                when others =>
                  \$16327\ := work.Print.print_string(clk,of_string("unknown primitive"));
                  \$16301\ := "000"& X"000000" & X"1" & eclat_true & \$13911\(0 to 15) & \$13911\(16 to 47) & 
                  work.Int.add(work.Int.sub(\$13911\(48 to 63), X"000" & X"1"), X"000" & X"1") & \$13911\(64 to 95) & \$13911\(96 to 103) & \$13911\(104 to 119) & \$13911\(120 to 121);
                  \$v7289\ := \$ram_lock\;
                  if \$v7289\(0) = '1' then
                    state_var7460 := Q_WAIT7288;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$16301\(80 to 95), X"000" & X"1")));
                    state_var7460 := PAUSE_GET7287;
                  end if;
                end case;
              when PAUSE_SET7301 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$16336\ := eclat_unit;
                \$v7300\ := \$15851_argument1\;
                case \$v7300\ is
                when "000"& X"000000" & X"0" =>
                  \$16353\ := work.Print.print_string(clk,of_string("======> "));
                  \$16357\ := work.Int.print(clk,\$13911\(16 to 46));
                  \$16358\ := work.Print.print_newline(clk,eclat_unit);
                  \$16337\ := "000"& X"000000" & X"1" & eclat_true & \$13911\(0 to 15) & \$13911\(16 to 47) & 
                  work.Int.add(work.Int.sub(work.Int.sub(\$13911\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1") & \$13911\(64 to 95) & \$13911\(96 to 103) & \$13911\(104 to 119) & \$13911\(120 to 121);
                  \$v7299\ := \$ram_lock\;
                  if \$v7299\(0) = '1' then
                    state_var7460 := Q_WAIT7298;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$16337\(80 to 95), X"000" & X"1")));
                    state_var7460 := PAUSE_GET7297;
                  end if;
                when others =>
                  \$16365\ := work.Print.print_string(clk,of_string("unknown primitive"));
                  \$16337\ := "000"& X"000000" & X"1" & eclat_true & \$13911\(0 to 15) & \$13911\(16 to 47) & 
                  work.Int.add(work.Int.sub(work.Int.sub(\$13911\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1") & \$13911\(64 to 95) & \$13911\(96 to 103) & \$13911\(104 to 119) & \$13911\(120 to 121);
                  \$v7299\ := \$ram_lock\;
                  if \$v7299\(0) = '1' then
                    state_var7460 := Q_WAIT7298;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$16337\(80 to 95), X"000" & X"1")));
                    state_var7460 := PAUSE_GET7297;
                  end if;
                end case;
              when PAUSE_SET7314 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$16382\ := eclat_unit;
                \$v7313\ := \$15851_argument1\;
                case \$v7313\ is
                when "000"& X"000000" & X"0" =>
                  \$16399\ := work.Print.print_string(clk,of_string("======> "));
                  \$16403\ := work.Int.print(clk,\$13911\(16 to 46));
                  \$16404\ := work.Print.print_newline(clk,eclat_unit);
                  \$16383\ := "000"& X"000000" & X"1" & eclat_true & \$13911\(0 to 15) & \$13911\(16 to 47) & 
                  work.Int.add(work.Int.sub(work.Int.sub(work.Int.sub(
                                                         \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1"), X"000" & X"1") & \$13911\(64 to 95) & \$13911\(96 to 103) & \$13911\(104 to 119) & \$13911\(120 to 121);
                  \$v7312\ := \$ram_lock\;
                  if \$v7312\(0) = '1' then
                    state_var7460 := Q_WAIT7311;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$16383\(80 to 95), X"000" & X"1")));
                    state_var7460 := PAUSE_GET7310;
                  end if;
                when others =>
                  \$16413\ := work.Print.print_string(clk,of_string("unknown primitive"));
                  \$16383\ := "000"& X"000000" & X"1" & eclat_true & \$13911\(0 to 15) & \$13911\(16 to 47) & 
                  work.Int.add(work.Int.sub(work.Int.sub(work.Int.sub(
                                                         \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1"), X"000" & X"1") & \$13911\(64 to 95) & \$13911\(96 to 103) & \$13911\(104 to 119) & \$13911\(120 to 121);
                  \$v7312\ := \$ram_lock\;
                  if \$v7312\(0) = '1' then
                    state_var7460 := Q_WAIT7311;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$16383\(80 to 95), X"000" & X"1")));
                    state_var7460 := PAUSE_GET7310;
                  end if;
                end case;
              when PAUSE_SET7330 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$16440\ := eclat_unit;
                \$v7329\ := \$15851_argument1\;
                case \$v7329\ is
                when "000"& X"000000" & X"0" =>
                  \$16457\ := work.Print.print_string(clk,of_string("======> "));
                  \$16461\ := work.Int.print(clk,\$13911\(16 to 46));
                  \$16462\ := work.Print.print_newline(clk,eclat_unit);
                  \$16441\ := "000"& X"000000" & X"1" & eclat_true & \$13911\(0 to 15) & \$13911\(16 to 47) & 
                  work.Int.add(work.Int.sub(work.Int.sub(work.Int.sub(
                                                         work.Int.sub(
                                                         \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1"), X"000" & X"1"), X"000" & X"1") & \$13911\(64 to 95) & \$13911\(96 to 103) & \$13911\(104 to 119) & \$13911\(120 to 121);
                  \$v7328\ := \$ram_lock\;
                  if \$v7328\(0) = '1' then
                    state_var7460 := Q_WAIT7327;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$16441\(80 to 95), X"000" & X"1")));
                    state_var7460 := PAUSE_GET7326;
                  end if;
                when others =>
                  \$16473\ := work.Print.print_string(clk,of_string("unknown primitive"));
                  \$16441\ := "000"& X"000000" & X"1" & eclat_true & \$13911\(0 to 15) & \$13911\(16 to 47) & 
                  work.Int.add(work.Int.sub(work.Int.sub(work.Int.sub(
                                                         work.Int.sub(
                                                         \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1"), X"000" & X"1"), X"000" & X"1") & \$13911\(64 to 95) & \$13911\(96 to 103) & \$13911\(104 to 119) & \$13911\(120 to 121);
                  \$v7328\ := \$ram_lock\;
                  if \$v7328\(0) = '1' then
                    state_var7460 := Q_WAIT7327;
                  else
                    acquire(\$ram_lock\);
                    \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$16441\(80 to 95), X"000" & X"1")));
                    state_var7460 := PAUSE_GET7326;
                  end if;
                end case;
              when PAUSE_SET7345 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$16515\ := eclat_unit;
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"2") & \$15851_argument1\ & eclat_true & 
                work.Int.add(\$13911\(48 to 63), X"000" & X"1") & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_SET7348 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$16534\ := eclat_unit;
                result6468 := work.Int.add(\$13911\(0 to 15), X"000" & X"2") & "000"& X"000000" & X"1" & eclat_true & \$13911\(48 to 63) & \$13911\(64 to 119) & \$13911\(120 to 121);
                rdy6469 := eclat_true;
                state_var7460 := IDLE6470;
              when PAUSE_SET7359 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$16677\ := eclat_unit;
                \$16662_fill6535928_arg\ := work.Int.add(\$16662_fill6535928_arg\(0 to 15), X"000" & X"1") & 
                work.Int.sub(\$16662_fill6535928_arg\(16 to 31), X"000" & X"1") & \$16662_fill6535928_arg\(32 to 47) & \$16662_fill6535928_arg\(48 to 79);
                state_var7460 := \$16662_FILL6535928\;
              when PAUSE_SET7366 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$16658\ := eclat_unit;
                \$16662_fill6535928_id\ := "000010100111";
                \$16662_fill6535928_arg\ := X"000" & X"1" & \$16650_sp\ & eclat_resize(\$15851_argument1\,16) & \$16651\(64 to 95);
                state_var7460 := \$16662_FILL6535928\;
              when PAUSE_SET7369 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$16706\ := eclat_unit;
                \$16650_sp\ := work.Int.add(\$13911\(48 to 63), X"000" & X"1");
                \$13923_make_block579_id\ := "000010101000";
                \$13923_make_block579_arg\ := \$16650_sp\ & \$13911\(16 to 47) & \$13911\(64 to 95) & "11110111" & 
                work.Int.add(eclat_resize(\$15851_argument1\,16), X"000" & X"1");
                state_var7460 := \$13923_MAKE_BLOCK579\;
              when PAUSE_SET7385 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$16724\ := eclat_unit;
                \$v7384\ := \$ram_lock\;
                if \$v7384\(0) = '1' then
                  state_var7460 := Q_WAIT7383;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(X"3e80", eclat_resize(\$15851_argument1\,16))));
                  state_var7460 := PAUSE_GET7382;
                end if;
              when PAUSE_SET7388 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$16767\ := eclat_unit;
                \$16752_fill6545929_arg\ := work.Int.add(\$16752_fill6545929_arg\(0 to 15), X"000" & X"1") & 
                work.Int.sub(\$16752_fill6545929_arg\(16 to 31), X"000" & X"1") & \$16752_fill6545929_arg\(32 to 47) & \$16752_fill6545929_arg\(48 to 79);
                state_var7460 := \$16752_FILL6545929\;
              when PAUSE_SET7395 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$16748\ := eclat_unit;
                \$16752_fill6545929_id\ := "000010101001";
                \$16752_fill6545929_arg\ := X"000" & X"1" & \$13911\(48 to 63) & eclat_resize(\$15851_argument1\,16) & \$16741\(64 to 95);
                state_var7460 := \$16752_FILL6545929\;
              when PAUSE_SET7404 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$17032\ := eclat_unit;
                \$17018_w36575938_arg\ := work.Int.add(\$17018_w36575938_arg\(0 to 15), X"000" & X"1") & 
                work.Int.add(\$17018_w36575938_arg\(16 to 31), X"000" & X"1") & \$17018_w36575938_arg\(32 to 47) & \$17018_w36575938_arg\(48 to 79);
                state_var7460 := \$17018_W36575938\;
              when PAUSE_SET7408 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$17011\ := eclat_unit;
                \$17018_w36575938_id\ := "000010110111";
                \$17018_w36575938_arg\ := X"000" & X"1" & work.Int.add(
                                                          \$17009_sp\, X"000" & X"1") & eclat_resize(\$15851_argument1\,16) & \$17001\(64 to 95);
                state_var7460 := \$17018_W36575938\;
              when PAUSE_SET7411 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$17066\ := eclat_unit;
                \$17048_w16565937_arg\ := work.Int.add(\$17048_w16565937_arg\(0 to 15), X"000" & X"1") & \$17048_w16565937_arg\(16 to 31) & \$17048_w16565937_arg\(32 to 47) & \$17048_w16565937_arg\(48 to 79);
                state_var7460 := \$17048_W16565937\;
              when PAUSE_SET7417 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$17061\ := eclat_unit;
                \$v7416\ := \$code_lock\;
                if \$v7416\(0) = '1' then
                  state_var7460 := Q_WAIT7415;
                else
                  acquire(\$code_lock\);
                  \$code_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                  \$17048_w16565937_arg\(16 to 31), X"000" & X"3"), \$17048_w16565937_arg\(0 to 15))));
                  state_var7460 := PAUSE_GET7414;
                end if;
              when PAUSE_SET7421 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$17121\ := eclat_unit;
                \$17105_w06555936_arg\ := work.Int.add(\$17105_w06555936_arg\(0 to 15), X"000" & X"1") & 
                work.Int.sub(\$17105_w06555936_arg\(16 to 31), X"000" & X"1") & \$17105_w06555936_arg\(32 to 47) & \$17105_w06555936_arg\(48 to 63) & \$17105_w06555936_arg\(64 to 95);
                state_var7460 := \$17105_W06555936\;
              when PAUSE_SET7428 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$17008\ := eclat_unit;
                \$17105_w06555936_id\ := "000010111001";
                \$17105_w06555936_arg\ := X"000" & X"0" & \$17000_sp\ & eclat_resize(\$15851_argument1\,16) & eclat_resize(\$16624_argument2\,16) & \$17001\(64 to 95);
                state_var7460 := \$17105_W06555936\;
              when PAUSE_SET7431 =>
                \$ram_write_request\ <= '0';
                release(\$ram_lock\);
                \$17161\ := eclat_unit;
                \$17000_sp\ := work.Int.add(\$13911\(48 to 63), X"000" & X"1");
                \$13923_make_block579_id\ := "000010111010";
                \$13923_make_block579_arg\ := \$17000_sp\ & \$13911\(16 to 47) & \$13911\(64 to 95) & "11110111" & 
                work.Int.add(work.Int.sub(work.Int.mul(X"000" & X"2", eclat_resize(\$15851_argument1\,16)), X"000" & X"1"), eclat_resize(\$16624_argument2\,16));
                state_var7460 := \$13923_MAKE_BLOCK579\;
              when Q_WAIT6472 =>
                \$v6473\ := \$ram_lock\;
                if \$v6473\(0) = '1' then
                  state_var7460 := Q_WAIT6472;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$13920_loop666_arg\(16 to 31), \$13920_loop666_arg\(0 to 15))));
                  \$ram_write\ <= \$18545\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6471;
                end if;
              when Q_WAIT6475 =>
                \$v6476\ := \$ram_lock\;
                if \$v6476\(0) = '1' then
                  state_var7460 := Q_WAIT6475;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$13920_loop666_arg\(32 to 47), \$13920_loop666_arg\(0 to 15))));
                  state_var7460 := PAUSE_GET6474;
                end if;
              when Q_WAIT6479 =>
                \$v6480\ := \$ram_lock\;
                if \$v6480\(0) = '1' then
                  state_var7460 := Q_WAIT6479;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$13921_loop665_arg\(64 to 79), \$13921_loop665_arg\(0 to 15))));
                  \$ram_write\ <= \$18447\(0 to 31); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6478;
                end if;
              when Q_WAIT6482 =>
                \$v6483\ := \$ram_lock\;
                if \$v6483\(0) = '1' then
                  state_var7460 := Q_WAIT6482;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          eclat_resize(\$18443\(0 to 30),16), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$13921_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6481;
                end if;
              when Q_WAIT6485 =>
                \$v6486\ := \$ram_lock\;
                if \$v6486\(0) = '1' then
                  state_var7460 := Q_WAIT6485;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$18443\(0 to 30),16)));
                  \$ram_write\ <= eclat_resize(\$13921_loop665_arg\(16 to 31),31) & eclat_false; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6484;
                end if;
              when Q_WAIT6488 =>
                \$v6489\ := \$ram_lock\;
                if \$v6489\(0) = '1' then
                  state_var7460 := Q_WAIT6488;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13921_loop665_arg\(16 to 31)));
                  \$ram_write\ <= \$18464_hd\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6487;
                end if;
              when Q_WAIT6491 =>
                \$v6492\ := \$ram_lock\;
                if \$v6492\(0) = '1' then
                  state_var7460 := Q_WAIT6491;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$18443\(0 to 30),16)));
                  state_var7460 := PAUSE_GET6490;
                end if;
              when Q_WAIT6495 =>
                \$v6496\ := \$ram_lock\;
                if \$v6496\(0) = '1' then
                  state_var7460 := Q_WAIT6495;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(eclat_resize(\$18443\(0 to 30),16), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6494;
                end if;
              when Q_WAIT6499 =>
                \$v6500\ := \$ram_lock\;
                if \$v6500\(0) = '1' then
                  state_var7460 := Q_WAIT6499;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(\$13921_loop665_arg\(64 to 79), \$13921_loop665_arg\(0 to 15))));
                  state_var7460 := PAUSE_GET6498;
                end if;
              when Q_WAIT6713 =>
                \$v6714\ := \$ram_lock\;
                if \$v6714\(0) = '1' then
                  state_var7460 := Q_WAIT6713;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$17389\(64 to 79)));
                  \$ram_write\ <= work.Int.lor(work.Int.lsl(eclat_resize(\$13923_make_block579_arg\(80 to 87),31), X"000000" & X"18"), 
                                               work.Int.lsl(eclat_resize(
                                                            eclat_if(
                                                            work.Int.eq(
                                                            \$13923_make_block579_arg\(88 to 103), X"000" & X"0") & X"000" & X"1" & \$13923_make_block579_arg\(88 to 103)),31), X"0000000" & X"2")) & eclat_true; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6712;
                end if;
              when Q_WAIT6716 =>
                \$v6717\ := \$ram_lock\;
                if \$v6717\(0) = '1' then
                  state_var7460 := Q_WAIT6716;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13924_apply638_arg\(60 to 90),16), X"000" & X"0"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6715;
                end if;
              when Q_WAIT6719 =>
                \$v6720\ := \$ram_lock\;
                if \$v6720\(0) = '1' then
                  state_var7460 := Q_WAIT6719;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$17332_sp\));
                  \$ram_write\ <= \$17321\(0 to 31); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6718;
                end if;
              when Q_WAIT6723 =>
                \$v6724\ := \$ram_lock\;
                if \$v6724\(0) = '1' then
                  state_var7460 := Q_WAIT6723;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$17331_sp\));
                  \$ram_write\ <= \$17324\(0 to 31); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6722;
                end if;
              when Q_WAIT6727 =>
                \$v6728\ := \$ram_lock\;
                if \$v6728\(0) = '1' then
                  state_var7460 := Q_WAIT6727;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$17330_sp\));
                  \$ram_write\ <= \$17327\(0 to 31); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6726;
                end if;
              when Q_WAIT6731 =>
                \$v6732\ := \$ram_lock\;
                if \$v6732\(0) = '1' then
                  state_var7460 := Q_WAIT6731;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          \$17327\(32 to 47), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(work.Int.add(\$13924_apply638_arg\(44 to 59), X"000" & X"1"),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6730;
                end if;
              when Q_WAIT6734 =>
                \$v6735\ := \$ram_lock\;
                if \$v6735\(0) = '1' then
                  state_var7460 := Q_WAIT6734;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$17327\(32 to 47), X"000" & X"1")));
                  \$ram_write\ <= \$13924_apply638_arg\(110 to 141); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6733;
                end if;
              when Q_WAIT6737 =>
                \$v6738\ := \$ram_lock\;
                if \$v6738\(0) = '1' then
                  state_var7460 := Q_WAIT6737;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$17327\(32 to 47)));
                  \$ram_write\ <= eclat_resize(\$13924_apply638_arg\(142 to 149),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6736;
                end if;
              when Q_WAIT6741 =>
                \$v6742\ := \$ram_lock\;
                if \$v6742\(0) = '1' then
                  state_var7460 := Q_WAIT6741;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$17324\(32 to 47), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6740;
                end if;
              when Q_WAIT6745 =>
                \$v6746\ := \$ram_lock\;
                if \$v6746\(0) = '1' then
                  state_var7460 := Q_WAIT6745;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$17321\(32 to 47), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6744;
                end if;
              when Q_WAIT6749 =>
                \$v6750\ := \$ram_lock\;
                if \$v6750\(0) = '1' then
                  state_var7460 := Q_WAIT6749;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13924_apply638_arg\(92 to 107), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6748;
                end if;
              when Q_WAIT6754 =>
                \$v6755\ := \$ram_lock\;
                if \$v6755\(0) = '1' then
                  state_var7460 := Q_WAIT6754;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$17232\(64 to 94),16), X"000" & X"2"), X"000" & X"1")));
                  \$ram_write\ <= \$17239_v\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6753;
                end if;
              when Q_WAIT6757 =>
                \$v6758\ := \$ram_lock\;
                if \$v6758\(0) = '1' then
                  state_var7460 := Q_WAIT6757;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$17237_sp\, X"000" & X"1")));
                  state_var7460 := PAUSE_GET6756;
                end if;
              when Q_WAIT6761 =>
                \$v6762\ := \$ram_lock\;
                if \$v6762\(0) = '1' then
                  state_var7460 := Q_WAIT6761;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$17232\(64 to 94),16), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= \$17250_v\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6760;
                end if;
              when Q_WAIT6764 =>
                \$v6765\ := \$ram_lock\;
                if \$v6765\(0) = '1' then
                  state_var7460 := Q_WAIT6764;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13926_make_block_n646_arg\(16 to 31), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6763;
                end if;
              when Q_WAIT6768 =>
                \$v6769\ := \$ram_lock\;
                if \$v6769\(0) = '1' then
                  state_var7460 := Q_WAIT6768;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$17232\(64 to 94),16), X"000" & X"0"), X"000" & X"1")));
                  \$ram_write\ <= \$17232\(0 to 31); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6767;
                end if;
              when Q_WAIT6772 =>
                \$v6773\ := \$code_lock\;
                if \$v6773\(0) = '1' then
                  state_var7460 := Q_WAIT6772;
                else
                  acquire(\$code_lock\);
                  \$code_ptr\ <= to_integer(unsigned(work.Int.add(\$13927_branch_if648_arg\(1 to 16), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6771;
                end if;
              when Q_WAIT6776 =>
                \$v6777\ := \$ram_lock\;
                if \$v6777\(0) = '1' then
                  state_var7460 := Q_WAIT6776;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.sub(
                                                          work.Int.sub(
                                                          work.Int.sub(
                                                          \$13928_w652_arg\(16 to 31), \$13928_w652_arg\(32 to 47)), \$13928_w652_arg\(48 to 63)), \$13928_w652_arg\(0 to 15))));
                  \$ram_write\ <= \$17183\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6775;
                end if;
              when Q_WAIT6779 =>
                \$v6780\ := \$ram_lock\;
                if \$v6780\(0) = '1' then
                  state_var7460 := Q_WAIT6779;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13928_w652_arg\(16 to 31), \$13928_w652_arg\(0 to 15))));
                  state_var7460 := PAUSE_GET6778;
                end if;
              when Q_WAIT6783 =>
                \$v6784\ := \$ram_lock\;
                if \$v6784\(0) = '1' then
                  state_var7460 := Q_WAIT6783;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$13911\(48 to 63), X"000" & X"0"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6782;
                end if;
              when Q_WAIT6786 =>
                \$v6787\ := \$ram_lock\;
                if \$v6787\(0) = '1' then
                  state_var7460 := Q_WAIT6786;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6785;
                end if;
              when Q_WAIT6789 =>
                \$v6790\ := \$ram_lock\;
                if \$v6790\(0) = '1' then
                  state_var7460 := Q_WAIT6789;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$13911\(48 to 63), X"000" & X"2"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6788;
                end if;
              when Q_WAIT6792 =>
                \$v6793\ := \$ram_lock\;
                if \$v6793\(0) = '1' then
                  state_var7460 := Q_WAIT6792;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$13911\(48 to 63), X"000" & X"3"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6791;
                end if;
              when Q_WAIT6795 =>
                \$v6796\ := \$ram_lock\;
                if \$v6796\(0) = '1' then
                  state_var7460 := Q_WAIT6795;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$13911\(48 to 63), X"000" & X"4"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6794;
                end if;
              when Q_WAIT6798 =>
                \$v6799\ := \$ram_lock\;
                if \$v6799\(0) = '1' then
                  state_var7460 := Q_WAIT6798;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$13911\(48 to 63), X"000" & X"5"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6797;
                end if;
              when Q_WAIT6801 =>
                \$v6802\ := \$ram_lock\;
                if \$v6802\(0) = '1' then
                  state_var7460 := Q_WAIT6801;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$13911\(48 to 63), X"000" & X"6"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6800;
                end if;
              when Q_WAIT6804 =>
                \$v6805\ := \$ram_lock\;
                if \$v6805\(0) = '1' then
                  state_var7460 := Q_WAIT6804;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$13911\(48 to 63), X"000" & X"7"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6803;
                end if;
              when Q_WAIT6807 =>
                \$v6808\ := \$ram_lock\;
                if \$v6808\(0) = '1' then
                  state_var7460 := Q_WAIT6807;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6806;
                end if;
              when Q_WAIT6810 =>
                \$v6811\ := \$ram_lock\;
                if \$v6811\(0) = '1' then
                  state_var7460 := Q_WAIT6810;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6809;
                end if;
              when Q_WAIT6813 =>
                \$v6814\ := \$ram_lock\;
                if \$v6814\(0) = '1' then
                  state_var7460 := Q_WAIT6813;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6812;
                end if;
              when Q_WAIT6816 =>
                \$v6817\ := \$ram_lock\;
                if \$v6817\(0) = '1' then
                  state_var7460 := Q_WAIT6816;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6815;
                end if;
              when Q_WAIT6819 =>
                \$v6820\ := \$ram_lock\;
                if \$v6820\(0) = '1' then
                  state_var7460 := Q_WAIT6819;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"2"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6818;
                end if;
              when Q_WAIT6822 =>
                \$v6823\ := \$ram_lock\;
                if \$v6823\(0) = '1' then
                  state_var7460 := Q_WAIT6822;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6821;
                end if;
              when Q_WAIT6825 =>
                \$v6826\ := \$ram_lock\;
                if \$v6826\(0) = '1' then
                  state_var7460 := Q_WAIT6825;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"3"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6824;
                end if;
              when Q_WAIT6828 =>
                \$v6829\ := \$ram_lock\;
                if \$v6829\(0) = '1' then
                  state_var7460 := Q_WAIT6828;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6827;
                end if;
              when Q_WAIT6831 =>
                \$v6832\ := \$ram_lock\;
                if \$v6832\(0) = '1' then
                  state_var7460 := Q_WAIT6831;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"4"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6830;
                end if;
              when Q_WAIT6834 =>
                \$v6835\ := \$ram_lock\;
                if \$v6835\(0) = '1' then
                  state_var7460 := Q_WAIT6834;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6833;
                end if;
              when Q_WAIT6837 =>
                \$v6838\ := \$ram_lock\;
                if \$v6838\(0) = '1' then
                  state_var7460 := Q_WAIT6837;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"5"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6836;
                end if;
              when Q_WAIT6840 =>
                \$v6841\ := \$ram_lock\;
                if \$v6841\(0) = '1' then
                  state_var7460 := Q_WAIT6840;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6839;
                end if;
              when Q_WAIT6843 =>
                \$v6844\ := \$ram_lock\;
                if \$v6844\(0) = '1' then
                  state_var7460 := Q_WAIT6843;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"6"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6842;
                end if;
              when Q_WAIT6846 =>
                \$v6847\ := \$ram_lock\;
                if \$v6847\(0) = '1' then
                  state_var7460 := Q_WAIT6846;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6845;
                end if;
              when Q_WAIT6849 =>
                \$v6850\ := \$ram_lock\;
                if \$v6850\(0) = '1' then
                  state_var7460 := Q_WAIT6849;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"7"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6848;
                end if;
              when Q_WAIT6852 =>
                \$v6853\ := \$ram_lock\;
                if \$v6853\(0) = '1' then
                  state_var7460 := Q_WAIT6852;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6851;
                end if;
              when Q_WAIT6855 =>
                \$v6856\ := \$ram_lock\;
                if \$v6856\(0) = '1' then
                  state_var7460 := Q_WAIT6855;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13911\(64 to 94),16), 
                                                                 work.Int.sub(
                                                                 X"000" & X"1", X"000" & X"1")), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6854;
                end if;
              when Q_WAIT6858 =>
                \$v6859\ := \$ram_lock\;
                if \$v6859\(0) = '1' then
                  state_var7460 := Q_WAIT6858;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13911\(64 to 94),16), 
                                                                 work.Int.sub(
                                                                 X"000" & X"2", X"000" & X"1")), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6857;
                end if;
              when Q_WAIT6861 =>
                \$v6862\ := \$ram_lock\;
                if \$v6862\(0) = '1' then
                  state_var7460 := Q_WAIT6861;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13911\(64 to 94),16), 
                                                                 work.Int.sub(
                                                                 X"000" & X"3", X"000" & X"1")), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6860;
                end if;
              when Q_WAIT6864 =>
                \$v6865\ := \$ram_lock\;
                if \$v6865\(0) = '1' then
                  state_var7460 := Q_WAIT6864;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13911\(64 to 94),16), 
                                                                 work.Int.sub(
                                                                 X"000" & X"4", X"000" & X"1")), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6863;
                end if;
              when Q_WAIT6867 =>
                \$v6868\ := \$ram_lock\;
                if \$v6868\(0) = '1' then
                  state_var7460 := Q_WAIT6867;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13911\(64 to 94),16), 
                                                                 work.Int.sub(
                                                                 X"000" & X"1", X"000" & X"1")), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6866;
                end if;
              when Q_WAIT6870 =>
                \$v6871\ := \$ram_lock\;
                if \$v6871\(0) = '1' then
                  state_var7460 := Q_WAIT6870;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6869;
                end if;
              when Q_WAIT6873 =>
                \$v6874\ := \$ram_lock\;
                if \$v6874\(0) = '1' then
                  state_var7460 := Q_WAIT6873;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13911\(64 to 94),16), 
                                                                 work.Int.sub(
                                                                 X"000" & X"2", X"000" & X"1")), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6872;
                end if;
              when Q_WAIT6876 =>
                \$v6877\ := \$ram_lock\;
                if \$v6877\(0) = '1' then
                  state_var7460 := Q_WAIT6876;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6875;
                end if;
              when Q_WAIT6879 =>
                \$v6880\ := \$ram_lock\;
                if \$v6880\(0) = '1' then
                  state_var7460 := Q_WAIT6879;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13911\(64 to 94),16), 
                                                                 work.Int.sub(
                                                                 X"000" & X"3", X"000" & X"1")), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6878;
                end if;
              when Q_WAIT6882 =>
                \$v6883\ := \$ram_lock\;
                if \$v6883\(0) = '1' then
                  state_var7460 := Q_WAIT6882;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6881;
                end if;
              when Q_WAIT6885 =>
                \$v6886\ := \$ram_lock\;
                if \$v6886\(0) = '1' then
                  state_var7460 := Q_WAIT6885;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13911\(64 to 94),16), 
                                                                 work.Int.sub(
                                                                 X"000" & X"4", X"000" & X"1")), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6884;
                end if;
              when Q_WAIT6888 =>
                \$v6889\ := \$ram_lock\;
                if \$v6889\(0) = '1' then
                  state_var7460 := Q_WAIT6888;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6887;
                end if;
              when Q_WAIT6891 =>
                \$v6892\ := \$ram_lock\;
                if \$v6892\(0) = '1' then
                  state_var7460 := Q_WAIT6891;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13911\(64 to 94),16), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6890;
                end if;
              when Q_WAIT6894 =>
                \$v6895\ := \$ram_lock\;
                if \$v6895\(0) = '1' then
                  state_var7460 := Q_WAIT6894;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$14207_loop_push6495899_arg\(0 to 15)));
                  \$ram_write\ <= \$14221\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6893;
                end if;
              when Q_WAIT6897 =>
                \$v6898\ := \$ram_lock\;
                if \$v6898\(0) = '1' then
                  state_var7460 := Q_WAIT6897;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$14207_loop_push6495899_arg\(24 to 54),16), eclat_resize(
                                                                 work.Int.add(
                                                                 \$14207_loop_push6495899_arg\(16 to 23), "00000010"),16)), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6896;
                end if;
              when Q_WAIT6901 =>
                \$v6902\ := \$ram_lock\;
                if \$v6902\(0) = '1' then
                  state_var7460 := Q_WAIT6901;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$13911\(64 to 94),16)));
                  state_var7460 := PAUSE_GET6900;
                end if;
              when Q_WAIT6904 =>
                \$v6905\ := \$ram_lock\;
                if \$v6905\(0) = '1' then
                  state_var7460 := Q_WAIT6904;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6903;
                end if;
              when Q_WAIT6907 =>
                \$v6908\ := \$ram_lock\;
                if \$v6908\(0) = '1' then
                  state_var7460 := Q_WAIT6907;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6906;
                end if;
              when Q_WAIT6910 =>
                \$v6911\ := \$ram_lock\;
                if \$v6911\(0) = '1' then
                  state_var7460 := Q_WAIT6910;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6909;
                end if;
              when Q_WAIT6913 =>
                \$v6914\ := \$ram_lock\;
                if \$v6914\(0) = '1' then
                  state_var7460 := Q_WAIT6913;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6912;
                end if;
              when Q_WAIT6916 =>
                \$v6917\ := \$ram_lock\;
                if \$v6917\(0) = '1' then
                  state_var7460 := Q_WAIT6916;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13911\(16 to 46),16), X"000" & X"0"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6915;
                end if;
              when Q_WAIT6919 =>
                \$v6920\ := \$ram_lock\;
                if \$v6920\(0) = '1' then
                  state_var7460 := Q_WAIT6919;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13911\(16 to 46),16), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6918;
                end if;
              when Q_WAIT6922 =>
                \$v6923\ := \$ram_lock\;
                if \$v6923\(0) = '1' then
                  state_var7460 := Q_WAIT6922;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13911\(16 to 46),16), X"000" & X"2"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6921;
                end if;
              when Q_WAIT6925 =>
                \$v6926\ := \$ram_lock\;
                if \$v6926\(0) = '1' then
                  state_var7460 := Q_WAIT6925;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13911\(16 to 46),16), X"000" & X"3"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6924;
                end if;
              when Q_WAIT6928 =>
                \$v6929\ := \$ram_lock\;
                if \$v6929\(0) = '1' then
                  state_var7460 := Q_WAIT6928;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$13911\(16 to 46),16), X"000" & X"0"), X"000" & X"1")));
                  \$ram_write\ <= \$14338_v\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6927;
                end if;
              when Q_WAIT6931 =>
                \$v6932\ := \$ram_lock\;
                if \$v6932\(0) = '1' then
                  state_var7460 := Q_WAIT6931;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13911\(48 to 63), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6930;
                end if;
              when Q_WAIT6934 =>
                \$v6935\ := \$ram_lock\;
                if \$v6935\(0) = '1' then
                  state_var7460 := Q_WAIT6934;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$13911\(16 to 46),16), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= \$14351_v\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6933;
                end if;
              when Q_WAIT6937 =>
                \$v6938\ := \$ram_lock\;
                if \$v6938\(0) = '1' then
                  state_var7460 := Q_WAIT6937;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13911\(48 to 63), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6936;
                end if;
              when Q_WAIT6940 =>
                \$v6941\ := \$ram_lock\;
                if \$v6941\(0) = '1' then
                  state_var7460 := Q_WAIT6940;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$13911\(16 to 46),16), X"000" & X"2"), X"000" & X"1")));
                  \$ram_write\ <= \$14364_v\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6939;
                end if;
              when Q_WAIT6943 =>
                \$v6944\ := \$ram_lock\;
                if \$v6944\(0) = '1' then
                  state_var7460 := Q_WAIT6943;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13911\(48 to 63), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6942;
                end if;
              when Q_WAIT6946 =>
                \$v6947\ := \$ram_lock\;
                if \$v6947\(0) = '1' then
                  state_var7460 := Q_WAIT6946;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$13911\(16 to 46),16), X"000" & X"3"), X"000" & X"1")));
                  \$ram_write\ <= \$14377_v\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6945;
                end if;
              when Q_WAIT6949 =>
                \$v6950\ := \$ram_lock\;
                if \$v6950\(0) = '1' then
                  state_var7460 := Q_WAIT6949;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13911\(48 to 63), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6948;
                end if;
              when Q_WAIT6952 =>
                \$v6953\ := \$ram_lock\;
                if \$v6953\(0) = '1' then
                  state_var7460 := Q_WAIT6952;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$13911\(16 to 46),16)));
                  state_var7460 := PAUSE_GET6951;
                end if;
              when Q_WAIT6955 =>
                \$v6956\ := \$ram_lock\;
                if \$v6956\(0) = '1' then
                  state_var7460 := Q_WAIT6955;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13911\(16 to 46),16), eclat_resize(\$14406_v\(0 to 30),16)), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6954;
                end if;
              when Q_WAIT6958 =>
                \$v6959\ := \$ram_lock\;
                if \$v6959\(0) = '1' then
                  state_var7460 := Q_WAIT6958;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13911\(48 to 63), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6957;
                end if;
              when Q_WAIT6961 =>
                \$v6962\ := \$ram_lock\;
                if \$v6962\(0) = '1' then
                  state_var7460 := Q_WAIT6961;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$13911\(16 to 46),16), eclat_resize(\$14423_v\(0 to 30),16)), X"000" & X"1")));
                  \$ram_write\ <= \$14424_v\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6960;
                end if;
              when Q_WAIT6964 =>
                \$v6965\ := \$ram_lock\;
                if \$v6965\(0) = '1' then
                  state_var7460 := Q_WAIT6964;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6963;
                end if;
              when Q_WAIT6967 =>
                \$v6968\ := \$ram_lock\;
                if \$v6968\(0) = '1' then
                  state_var7460 := Q_WAIT6967;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13911\(48 to 63), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6966;
                end if;
              when Q_WAIT6970 =>
                \$v6971\ := \$ram_lock\;
                if \$v6971\(0) = '1' then
                  state_var7460 := Q_WAIT6970;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13911\(16 to 46),16), eclat_resize(\$14446_v\(0 to 30),16)), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6969;
                end if;
              when Q_WAIT6973 =>
                \$v6974\ := \$ram_lock\;
                if \$v6974\(0) = '1' then
                  state_var7460 := Q_WAIT6973;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13911\(48 to 63), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6972;
                end if;
              when Q_WAIT6976 =>
                \$v6977\ := \$ram_lock\;
                if \$v6977\(0) = '1' then
                  state_var7460 := Q_WAIT6976;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$13911\(16 to 46),16), eclat_resize(\$14463_v\(0 to 30),16)), X"000" & X"1")));
                  \$ram_write\ <= \$14464_v\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6975;
                end if;
              when Q_WAIT6979 =>
                \$v6980\ := \$ram_lock\;
                if \$v6980\(0) = '1' then
                  state_var7460 := Q_WAIT6979;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6978;
                end if;
              when Q_WAIT6982 =>
                \$v6983\ := \$ram_lock\;
                if \$v6983\(0) = '1' then
                  state_var7460 := Q_WAIT6982;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13911\(48 to 63), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6981;
                end if;
              when Q_WAIT6985 =>
                \$v6986\ := \$ram_lock\;
                if \$v6986\(0) = '1' then
                  state_var7460 := Q_WAIT6985;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6984;
                end if;
              when Q_WAIT6988 =>
                \$v6989\ := \$ram_lock\;
                if \$v6989\(0) = '1' then
                  state_var7460 := Q_WAIT6988;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$13911\(104 to 119), X"000" & X"1"), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6987;
                end if;
              when Q_WAIT6991 =>
                \$v6992\ := \$ram_lock\;
                if \$v6992\(0) = '1' then
                  state_var7460 := Q_WAIT6991;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$13911\(104 to 119), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6990;
                end if;
              when Q_WAIT6994 =>
                \$v6995\ := \$ram_lock\;
                if \$v6995\(0) = '1' then
                  state_var7460 := Q_WAIT6994;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$13911\(104 to 119), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6993;
                end if;
              when Q_WAIT6997 =>
                \$v6998\ := \$ram_lock\;
                if \$v6998\(0) = '1' then
                  state_var7460 := Q_WAIT6997;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13911\(104 to 119), X"000" & X"1")));
                  state_var7460 := PAUSE_GET6996;
                end if;
              when Q_WAIT7000 =>
                \$v7001\ := \$ram_lock\;
                if \$v7001\(0) = '1' then
                  state_var7460 := Q_WAIT7000;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET6999;
                end if;
              when Q_WAIT7003 =>
                \$v7004\ := \$ram_lock\;
                if \$v7004\(0) = '1' then
                  state_var7460 := Q_WAIT7003;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7002;
                end if;
              when Q_WAIT7006 =>
                \$v7007\ := \$ram_lock\;
                if \$v7007\(0) = '1' then
                  state_var7460 := Q_WAIT7006;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7005;
                end if;
              when Q_WAIT7009 =>
                \$v7010\ := \$ram_lock\;
                if \$v7010\(0) = '1' then
                  state_var7460 := Q_WAIT7009;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7008;
                end if;
              when Q_WAIT7019 =>
                \$v7020\ := \$ram_lock\;
                if \$v7020\(0) = '1' then
                  state_var7460 := Q_WAIT7019;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$14564_binop_int6435900_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7018;
                end if;
              when Q_WAIT7029 =>
                \$v7030\ := \$ram_lock\;
                if \$v7030\(0) = '1' then
                  state_var7460 := Q_WAIT7029;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$14644_binop_int6435901_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7028;
                end if;
              when Q_WAIT7039 =>
                \$v7040\ := \$ram_lock\;
                if \$v7040\(0) = '1' then
                  state_var7460 := Q_WAIT7039;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$14724_binop_int6435902_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7038;
                end if;
              when Q_WAIT7049 =>
                \$v7050\ := \$ram_lock\;
                if \$v7050\(0) = '1' then
                  state_var7460 := Q_WAIT7049;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$14804_binop_int6435903_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7048;
                end if;
              when Q_WAIT7059 =>
                \$v7060\ := \$ram_lock\;
                if \$v7060\(0) = '1' then
                  state_var7460 := Q_WAIT7059;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$14884_binop_int6435904_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7058;
                end if;
              when Q_WAIT7069 =>
                \$v7070\ := \$ram_lock\;
                if \$v7070\(0) = '1' then
                  state_var7460 := Q_WAIT7069;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$14964_binop_int6435905_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7068;
                end if;
              when Q_WAIT7079 =>
                \$v7080\ := \$ram_lock\;
                if \$v7080\(0) = '1' then
                  state_var7460 := Q_WAIT7079;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$15044_binop_int6435906_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7078;
                end if;
              when Q_WAIT7089 =>
                \$v7090\ := \$ram_lock\;
                if \$v7090\(0) = '1' then
                  state_var7460 := Q_WAIT7089;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$15124_binop_int6435907_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7088;
                end if;
              when Q_WAIT7099 =>
                \$v7100\ := \$ram_lock\;
                if \$v7100\(0) = '1' then
                  state_var7460 := Q_WAIT7099;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$15204_binop_int6435908_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7098;
                end if;
              when Q_WAIT7109 =>
                \$v7110\ := \$ram_lock\;
                if \$v7110\(0) = '1' then
                  state_var7460 := Q_WAIT7109;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$15284_binop_int6435909_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7108;
                end if;
              when Q_WAIT7119 =>
                \$v7120\ := \$ram_lock\;
                if \$v7120\(0) = '1' then
                  state_var7460 := Q_WAIT7119;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$15364_binop_int6435910_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7118;
                end if;
              when Q_WAIT7129 =>
                \$v7130\ := \$ram_lock\;
                if \$v7130\(0) = '1' then
                  state_var7460 := Q_WAIT7129;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$15451_binop_int6435912_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7128;
                end if;
              when Q_WAIT7139 =>
                \$v7140\ := \$ram_lock\;
                if \$v7140\(0) = '1' then
                  state_var7460 := Q_WAIT7139;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$15531_binop_int6435913_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7138;
                end if;
              when Q_WAIT7143 =>
                \$v7144\ := \$ram_lock\;
                if \$v7144\(0) = '1' then
                  state_var7460 := Q_WAIT7143;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$15625_binop_compare6455916_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7142;
                end if;
              when Q_WAIT7147 =>
                \$v7148\ := \$ram_lock\;
                if \$v7148\(0) = '1' then
                  state_var7460 := Q_WAIT7147;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$15661_binop_compare6455917_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7146;
                end if;
              when Q_WAIT7151 =>
                \$v7152\ := \$ram_lock\;
                if \$v7152\(0) = '1' then
                  state_var7460 := Q_WAIT7151;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$15697_binop_compare6455918_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7150;
                end if;
              when Q_WAIT7155 =>
                \$v7156\ := \$ram_lock\;
                if \$v7156\(0) = '1' then
                  state_var7460 := Q_WAIT7155;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$15733_binop_compare6455919_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7154;
                end if;
              when Q_WAIT7159 =>
                \$v7160\ := \$ram_lock\;
                if \$v7160\(0) = '1' then
                  state_var7460 := Q_WAIT7159;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$15769_binop_compare6455920_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7158;
                end if;
              when Q_WAIT7163 =>
                \$v7164\ := \$ram_lock\;
                if \$v7164\(0) = '1' then
                  state_var7460 := Q_WAIT7163;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$15805_binop_compare6455921_arg\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7162;
                end if;
              when Q_WAIT7166 =>
                \$v7167\ := \$ram_lock\;
                if \$v7167\(0) = '1' then
                  state_var7460 := Q_WAIT7166;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$13911\(48 to 63), eclat_resize(\$15851_argument1\,16)), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7165;
                end if;
              when Q_WAIT7169 =>
                \$v7170\ := \$ram_lock\;
                if \$v7170\(0) = '1' then
                  state_var7460 := Q_WAIT7169;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.add(
                                                                 \$13911\(48 to 63), X"000" & X"1"), eclat_resize(\$15851_argument1\,16)), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7168;
                end if;
              when Q_WAIT7172 =>
                \$v7173\ := \$ram_lock\;
                if \$v7173\(0) = '1' then
                  state_var7460 := Q_WAIT7172;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7171;
                end if;
              when Q_WAIT7175 =>
                \$v7176\ := \$ram_lock\;
                if \$v7176\(0) = '1' then
                  state_var7460 := Q_WAIT7175;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.sub(
                                                          work.Int.sub(
                                                          \$13911\(48 to 63), X"000" & X"1"), eclat_resize(\$15851_argument1\,16))));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7174;
                end if;
              when Q_WAIT7178 =>
                \$v7179\ := \$ram_lock\;
                if \$v7179\(0) = '1' then
                  state_var7460 := Q_WAIT7178;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13911\(64 to 94),16), 
                                                                 work.Int.sub(
                                                                 eclat_resize(\$15851_argument1\,16), X"000" & X"1")), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7177;
                end if;
              when Q_WAIT7181 =>
                \$v7182\ := \$ram_lock\;
                if \$v7182\(0) = '1' then
                  state_var7460 := Q_WAIT7181;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13911\(64 to 94),16), 
                                                                 work.Int.sub(
                                                                 eclat_resize(\$15851_argument1\,16), X"000" & X"1")), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7180;
                end if;
              when Q_WAIT7184 =>
                \$v7185\ := \$ram_lock\;
                if \$v7185\(0) = '1' then
                  state_var7460 := Q_WAIT7184;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7183;
                end if;
              when Q_WAIT7187 =>
                \$v7188\ := \$ram_lock\;
                if \$v7188\(0) = '1' then
                  state_var7460 := Q_WAIT7187;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(work.Int.add(work.Int.add(
                                                            \$13911\(0 to 15), X"000" & X"1"), eclat_resize(\$15851_argument1\,16)),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7186;
                end if;
              when Q_WAIT7190 =>
                \$v7191\ := \$ram_lock\;
                if \$v7191\(0) = '1' then
                  state_var7460 := Q_WAIT7190;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$13911\(48 to 63), X"000" & X"1")));
                  \$ram_write\ <= \$13911\(64 to 95); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7189;
                end if;
              when Q_WAIT7193 =>
                \$v7194\ := \$ram_lock\;
                if \$v7194\(0) = '1' then
                  state_var7460 := Q_WAIT7193;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= eclat_resize(\$13911\(96 to 103),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7192;
                end if;
              when Q_WAIT7196 =>
                \$v7197\ := \$ram_lock\;
                if \$v7197\(0) = '1' then
                  state_var7460 := Q_WAIT7196;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13911\(16 to 46),16), X"000" & X"0"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7195;
                end if;
              when Q_WAIT7199 =>
                \$v7200\ := \$ram_lock\;
                if \$v7200\(0) = '1' then
                  state_var7460 := Q_WAIT7199;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13911\(16 to 46),16), X"000" & X"0"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7198;
                end if;
              when Q_WAIT7202 =>
                \$v7203\ := \$ram_lock\;
                if \$v7203\(0) = '1' then
                  state_var7460 := Q_WAIT7202;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$13911\(48 to 63), eclat_resize(\$15851_argument1\,16)), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7201;
                end if;
              when Q_WAIT7205 =>
                \$v7206\ := \$ram_lock\;
                if \$v7206\(0) = '1' then
                  state_var7460 := Q_WAIT7205;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$13911\(48 to 63), eclat_resize(\$15851_argument1\,16)), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7204;
                end if;
              when Q_WAIT7208 =>
                \$v7209\ := \$ram_lock\;
                if \$v7209\(0) = '1' then
                  state_var7460 := Q_WAIT7208;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$13911\(48 to 63), eclat_resize(\$15851_argument1\,16)), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7207;
                end if;
              when Q_WAIT7212 =>
                \$v7213\ := \$ram_lock\;
                if \$v7213\(0) = '1' then
                  state_var7460 := Q_WAIT7212;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$16036_sp\, X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7211;
                end if;
              when Q_WAIT7215 =>
                \$v7216\ := \$ram_lock\;
                if \$v7216\(0) = '1' then
                  state_var7460 := Q_WAIT7215;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$16036_sp\, X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7214;
                end if;
              when Q_WAIT7218 =>
                \$v7219\ := \$ram_lock\;
                if \$v7219\(0) = '1' then
                  state_var7460 := Q_WAIT7218;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$16036_sp\, X"000" & X"1")));
                  state_var7460 := PAUSE_GET7217;
                end if;
              when Q_WAIT7221 =>
                \$v7222\ := \$ram_lock\;
                if \$v7222\(0) = '1' then
                  state_var7460 := Q_WAIT7221;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$16063_w6515922_arg\(32 to 62),16), eclat_resize(
                                                          work.Int.add(
                                                          \$16063_w6515922_arg\(0 to 7), "00000010"),16)), X"000" & X"1")));
                  \$ram_write\ <= \$16074_v\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7220;
                end if;
              when Q_WAIT7224 =>
                \$v7225\ := \$ram_lock\;
                if \$v7225\(0) = '1' then
                  state_var7460 := Q_WAIT7224;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$16063_w6515922_arg\(8 to 23), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7223;
                end if;
              when Q_WAIT7228 =>
                \$v7229\ := \$ram_lock\;
                if \$v7229\(0) = '1' then
                  state_var7460 := Q_WAIT7228;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$16024\(64 to 94),16), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= \$16024\(32 to 63); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7227;
                end if;
              when Q_WAIT7231 =>
                \$v7232\ := \$ram_lock\;
                if \$v7232\(0) = '1' then
                  state_var7460 := Q_WAIT7231;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$16024\(64 to 94),16), X"000" & X"0"), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(work.Int.sub(work.Int.add(
                                                            \$13911\(0 to 15), X"000" & X"2"), X"000" & X"3"),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7230;
                end if;
              when Q_WAIT7235 =>
                \$v7236\ := \$ram_lock\;
                if \$v7236\(0) = '1' then
                  state_var7460 := Q_WAIT7235;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7234;
                end if;
              when Q_WAIT7238 =>
                \$v7239\ := \$ram_lock\;
                if \$v7239\(0) = '1' then
                  state_var7460 := Q_WAIT7238;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(X"3e80", eclat_resize(\$15851_argument1\,16))));
                  state_var7460 := PAUSE_GET7237;
                end if;
              when Q_WAIT7241 =>
                \$v7242\ := \$ram_lock\;
                if \$v7242\(0) = '1' then
                  state_var7460 := Q_WAIT7241;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(X"3e80", eclat_resize(\$15851_argument1\,16))));
                  state_var7460 := PAUSE_GET7240;
                end if;
              when Q_WAIT7244 =>
                \$v7245\ := \$ram_lock\;
                if \$v7245\(0) = '1' then
                  state_var7460 := Q_WAIT7244;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7243;
                end if;
              when Q_WAIT7247 =>
                \$v7248\ := \$ram_lock\;
                if \$v7248\(0) = '1' then
                  state_var7460 := Q_WAIT7247;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          X"3e80", eclat_resize(\$15851_argument1\,16))));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7246;
                end if;
              when Q_WAIT7250 =>
                \$v7251\ := \$ram_lock\;
                if \$v7251\(0) = '1' then
                  state_var7460 := Q_WAIT7250;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7249;
                end if;
              when Q_WAIT7253 =>
                \$v7254\ := \$ram_lock\;
                if \$v7254\(0) = '1' then
                  state_var7460 := Q_WAIT7253;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13911\(16 to 46),16), eclat_resize(\$15851_argument1\,16)), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7252;
                end if;
              when Q_WAIT7256 =>
                \$v7257\ := \$ram_lock\;
                if \$v7257\(0) = '1' then
                  state_var7460 := Q_WAIT7256;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$13911\(16 to 46),16), eclat_resize(\$15851_argument1\,16)), X"000" & X"1")));
                  \$ram_write\ <= \$16178_v\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7255;
                end if;
              when Q_WAIT7259 =>
                \$v7260\ := \$ram_lock\;
                if \$v7260\(0) = '1' then
                  state_var7460 := Q_WAIT7259;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13911\(48 to 63), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7258;
                end if;
              when Q_WAIT7262 =>
                \$v7263\ := \$code_lock\;
                if \$v7263\(0) = '1' then
                  state_var7460 := Q_WAIT7262;
                else
                  acquire(\$code_lock\);
                  \$code_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                  \$13911\(0 to 15), X"000" & X"2"), \$16202_ofs\)));
                  state_var7460 := PAUSE_GET7261;
                end if;
              when Q_WAIT7265 =>
                \$v7266\ := \$ram_lock\;
                if \$v7266\(0) = '1' then
                  state_var7460 := Q_WAIT7265;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$13911\(16 to 46),16)));
                  state_var7460 := PAUSE_GET7264;
                end if;
              when Q_WAIT7269 =>
                \$v7270\ := \$ram_lock\;
                if \$v7270\(0) = '1' then
                  state_var7460 := Q_WAIT7269;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          work.Int.add(
                                                          \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(work.Int.add(work.Int.add(
                                                            \$13911\(0 to 15), X"000" & X"1"), eclat_resize(\$15851_argument1\,16)),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7268;
                end if;
              when Q_WAIT7272 =>
                \$v7273\ := \$ram_lock\;
                if \$v7273\(0) = '1' then
                  state_var7460 := Q_WAIT7272;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(\$13911\(104 to 119),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7271;
                end if;
              when Q_WAIT7275 =>
                \$v7276\ := \$ram_lock\;
                if \$v7276\(0) = '1' then
                  state_var7460 := Q_WAIT7275;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          \$13911\(48 to 63), X"000" & X"1")));
                  \$ram_write\ <= \$13911\(64 to 95); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7274;
                end if;
              when Q_WAIT7278 =>
                \$v7279\ := \$ram_lock\;
                if \$v7279\(0) = '1' then
                  state_var7460 := Q_WAIT7278;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= eclat_resize(\$13911\(96 to 103),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7277;
                end if;
              when Q_WAIT7281 =>
                \$v7282\ := \$ram_lock\;
                if \$v7282\(0) = '1' then
                  state_var7460 := Q_WAIT7281;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$16272\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7280;
                end if;
              when Q_WAIT7285 =>
                \$v7286\ := \$ram_lock\;
                if \$v7286\(0) = '1' then
                  state_var7460 := Q_WAIT7285;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(64 to 95); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7284;
                end if;
              when Q_WAIT7288 =>
                \$v7289\ := \$ram_lock\;
                if \$v7289\(0) = '1' then
                  state_var7460 := Q_WAIT7288;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$16301\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7287;
                end if;
              when Q_WAIT7292 =>
                \$v7293\ := \$ram_lock\;
                if \$v7293\(0) = '1' then
                  state_var7460 := Q_WAIT7292;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.sub(
                                                          \$13911\(48 to 63), X"000" & X"1")));
                  \$ram_write\ <= \$13911\(64 to 95); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7291;
                end if;
              when Q_WAIT7295 =>
                \$v7296\ := \$ram_lock\;
                if \$v7296\(0) = '1' then
                  state_var7460 := Q_WAIT7295;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13911\(48 to 63), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7294;
                end if;
              when Q_WAIT7298 =>
                \$v7299\ := \$ram_lock\;
                if \$v7299\(0) = '1' then
                  state_var7460 := Q_WAIT7298;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$16337\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7297;
                end if;
              when Q_WAIT7302 =>
                \$v7303\ := \$ram_lock\;
                if \$v7303\(0) = '1' then
                  state_var7460 := Q_WAIT7302;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.sub(
                                                          work.Int.sub(
                                                          \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= \$13911\(64 to 95); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7301;
                end if;
              when Q_WAIT7305 =>
                \$v7306\ := \$ram_lock\;
                if \$v7306\(0) = '1' then
                  state_var7460 := Q_WAIT7305;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7304;
                end if;
              when Q_WAIT7308 =>
                \$v7309\ := \$ram_lock\;
                if \$v7309\(0) = '1' then
                  state_var7460 := Q_WAIT7308;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13911\(48 to 63), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7307;
                end if;
              when Q_WAIT7311 =>
                \$v7312\ := \$ram_lock\;
                if \$v7312\(0) = '1' then
                  state_var7460 := Q_WAIT7311;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$16383\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7310;
                end if;
              when Q_WAIT7315 =>
                \$v7316\ := \$ram_lock\;
                if \$v7316\(0) = '1' then
                  state_var7460 := Q_WAIT7315;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.sub(
                                                          work.Int.sub(
                                                          work.Int.sub(
                                                          \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= \$13911\(64 to 95); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7314;
                end if;
              when Q_WAIT7318 =>
                \$v7319\ := \$ram_lock\;
                if \$v7319\(0) = '1' then
                  state_var7460 := Q_WAIT7318;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7317;
                end if;
              when Q_WAIT7321 =>
                \$v7322\ := \$ram_lock\;
                if \$v7322\(0) = '1' then
                  state_var7460 := Q_WAIT7321;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7320;
                end if;
              when Q_WAIT7324 =>
                \$v7325\ := \$ram_lock\;
                if \$v7325\(0) = '1' then
                  state_var7460 := Q_WAIT7324;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13911\(48 to 63), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7323;
                end if;
              when Q_WAIT7327 =>
                \$v7328\ := \$ram_lock\;
                if \$v7328\(0) = '1' then
                  state_var7460 := Q_WAIT7327;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$16441\(80 to 95), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7326;
                end if;
              when Q_WAIT7331 =>
                \$v7332\ := \$ram_lock\;
                if \$v7332\(0) = '1' then
                  state_var7460 := Q_WAIT7331;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.sub(
                                                          work.Int.sub(
                                                          work.Int.sub(
                                                          work.Int.sub(
                                                          \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  \$ram_write\ <= \$13911\(64 to 95); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7330;
                end if;
              when Q_WAIT7334 =>
                \$v7335\ := \$ram_lock\;
                if \$v7335\(0) = '1' then
                  state_var7460 := Q_WAIT7334;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7333;
                end if;
              when Q_WAIT7337 =>
                \$v7338\ := \$ram_lock\;
                if \$v7338\(0) = '1' then
                  state_var7460 := Q_WAIT7337;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 work.Int.sub(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7336;
                end if;
              when Q_WAIT7340 =>
                \$v7341\ := \$ram_lock\;
                if \$v7341\(0) = '1' then
                  state_var7460 := Q_WAIT7340;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(work.Int.sub(
                                                                 \$13911\(48 to 63), X"000" & X"1"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7339;
                end if;
              when Q_WAIT7343 =>
                \$v7344\ := \$ram_lock\;
                if \$v7344\(0) = '1' then
                  state_var7460 := Q_WAIT7343;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$13911\(48 to 63), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7342;
                end if;
              when Q_WAIT7346 =>
                \$v7347\ := \$ram_lock\;
                if \$v7347\(0) = '1' then
                  state_var7460 := Q_WAIT7346;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7345;
                end if;
              when Q_WAIT7349 =>
                \$v7350\ := \$ram_lock\;
                if \$v7350\(0) = '1' then
                  state_var7460 := Q_WAIT7349;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$13911\(16 to 46),16), X"000" & X"0"), X"000" & X"1")));
                  \$ram_write\ <= work.Int.add(\$16527_f0\(0 to 30), \$15851_argument1\) & eclat_true; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7348;
                end if;
              when Q_WAIT7352 =>
                \$v7353\ := \$ram_lock\;
                if \$v7353\(0) = '1' then
                  state_var7460 := Q_WAIT7352;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13911\(16 to 46),16), X"000" & X"0"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7351;
                end if;
              when Q_WAIT7357 =>
                \$v7358\ := \$ram_lock\;
                if \$v7358\(0) = '1' then
                  state_var7460 := Q_WAIT7357;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$13911\(16 to 46),16), X"000" & X"0"), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7356;
                end if;
              when Q_WAIT7360 =>
                \$v7361\ := \$ram_lock\;
                if \$v7361\(0) = '1' then
                  state_var7460 := Q_WAIT7360;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$16662_fill6535928_arg\(48 to 78),16), \$16662_fill6535928_arg\(0 to 15)), X"000" & X"1")));
                  \$ram_write\ <= \$16673_v\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7359;
                end if;
              when Q_WAIT7363 =>
                \$v7364\ := \$ram_lock\;
                if \$v7364\(0) = '1' then
                  state_var7460 := Q_WAIT7363;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$16662_fill6535928_arg\(16 to 31), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7362;
                end if;
              when Q_WAIT7367 =>
                \$v7368\ := \$ram_lock\;
                if \$v7368\(0) = '1' then
                  state_var7460 := Q_WAIT7367;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$16651\(64 to 94),16), X"000" & X"0"), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(work.Int.add(work.Int.add(
                                                            \$13911\(0 to 15), X"000" & X"2"), eclat_resize(\$16624_argument2\,16)),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7366;
                end if;
              when Q_WAIT7370 =>
                \$v7371\ := \$ram_lock\;
                if \$v7371\(0) = '1' then
                  state_var7460 := Q_WAIT7370;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7369;
                end if;
              when Q_WAIT7374 =>
                \$v7375\ := \$ram_lock\;
                if \$v7375\(0) = '1' then
                  state_var7460 := Q_WAIT7374;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$16709\(0 to 30),16), eclat_resize(\$16624_argument2\,16)), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7373;
                end if;
              when Q_WAIT7377 =>
                \$v7378\ := \$ram_lock\;
                if \$v7378\(0) = '1' then
                  state_var7460 := Q_WAIT7377;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(X"3e80", eclat_resize(\$15851_argument1\,16))));
                  state_var7460 := PAUSE_GET7376;
                end if;
              when Q_WAIT7380 =>
                \$v7381\ := \$ram_lock\;
                if \$v7381\(0) = '1' then
                  state_var7460 := Q_WAIT7380;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                 eclat_resize(\$16725\(0 to 30),16), eclat_resize(\$16624_argument2\,16)), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7379;
                end if;
              when Q_WAIT7383 =>
                \$v7384\ := \$ram_lock\;
                if \$v7384\(0) = '1' then
                  state_var7460 := Q_WAIT7383;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.add(X"3e80", eclat_resize(\$15851_argument1\,16))));
                  state_var7460 := PAUSE_GET7382;
                end if;
              when Q_WAIT7386 =>
                \$v7387\ := \$ram_lock\;
                if \$v7387\(0) = '1' then
                  state_var7460 := Q_WAIT7386;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7385;
                end if;
              when Q_WAIT7389 =>
                \$v7390\ := \$ram_lock\;
                if \$v7390\(0) = '1' then
                  state_var7460 := Q_WAIT7389;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$16752_fill6545929_arg\(48 to 78),16), \$16752_fill6545929_arg\(0 to 15)), X"000" & X"1")));
                  \$ram_write\ <= \$16763_v\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7388;
                end if;
              when Q_WAIT7392 =>
                \$v7393\ := \$ram_lock\;
                if \$v7393\(0) = '1' then
                  state_var7460 := Q_WAIT7392;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$16752_fill6545929_arg\(16 to 31), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7391;
                end if;
              when Q_WAIT7396 =>
                \$v7397\ := \$ram_lock\;
                if \$v7397\(0) = '1' then
                  state_var7460 := Q_WAIT7396;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$16741\(64 to 94),16), X"000" & X"0"), X"000" & X"1")));
                  \$ram_write\ <= \$16741\(0 to 31); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7395;
                end if;
              when Q_WAIT7405 =>
                \$v7406\ := \$ram_lock\;
                if \$v7406\(0) = '1' then
                  state_var7460 := Q_WAIT7405;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$17018_w36575938_arg\(16 to 31)));
                  \$ram_write\ <= eclat_resize(work.Int.add(eclat_resize(\$17018_w36575938_arg\(48 to 78),16), 
                                                            work.Int.mul(
                                                            X"000" & X"2", \$17018_w36575938_arg\(0 to 15))),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7404;
                end if;
              when Q_WAIT7409 =>
                \$v7410\ := \$ram_lock\;
                if \$v7410\(0) = '1' then
                  state_var7460 := Q_WAIT7409;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$17009_sp\));
                  \$ram_write\ <= \$17001\(64 to 95); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7408;
                end if;
              when Q_WAIT7412 =>
                \$v7413\ := \$ram_lock\;
                if \$v7413\(0) = '1' then
                  state_var7460 := Q_WAIT7412;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$17048_w16565937_arg\(48 to 78),16), 
                                                          work.Int.mul(
                                                          X"000" & X"2", \$17048_w16565937_arg\(0 to 15))), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(work.Int.add(work.Int.add(
                                                            \$17048_w16565937_arg\(16 to 31), X"000" & X"2"), eclat_resize(\$17062\,16)),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7411;
                end if;
              when Q_WAIT7415 =>
                \$v7416\ := \$code_lock\;
                if \$v7416\(0) = '1' then
                  state_var7460 := Q_WAIT7415;
                else
                  acquire(\$code_lock\);
                  \$code_ptr\ <= to_integer(unsigned(work.Int.add(work.Int.add(
                                                                  \$17048_w16565937_arg\(16 to 31), X"000" & X"3"), \$17048_w16565937_arg\(0 to 15))));
                  state_var7460 := PAUSE_GET7414;
                end if;
              when Q_WAIT7418 =>
                \$v7419\ := \$ram_lock\;
                if \$v7419\(0) = '1' then
                  state_var7460 := Q_WAIT7418;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$17048_w16565937_arg\(48 to 78),16), 
                                                          work.Int.sub(
                                                          work.Int.mul(
                                                          X"000" & X"2", \$17048_w16565937_arg\(0 to 15)), X"000" & X"1")), X"000" & X"1")));
                  \$ram_write\ <= work.Int.lor(work.Int.lsl(eclat_resize("11111001",31), X"000000" & X"18"), 
                                               work.Int.lsl(eclat_resize(
                                                            work.Int.mul(
                                                            X"000" & X"2", \$17048_w16565937_arg\(0 to 15)),31), X"0000000" & X"2")) & eclat_true; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7417;
                end if;
              when Q_WAIT7422 =>
                \$v7423\ := \$ram_lock\;
                if \$v7423\(0) = '1' then
                  state_var7460 := Q_WAIT7422;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$17105_w06555936_arg\(64 to 94),16), 
                                                          work.Int.sub(
                                                          work.Int.add(
                                                          \$17105_w06555936_arg\(0 to 15), 
                                                          work.Int.mul(
                                                          X"000" & X"2", \$17105_w06555936_arg\(32 to 47))), X"000" & X"1")), X"000" & X"1")));
                  \$ram_write\ <= \$17117_v\; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7421;
                end if;
              when Q_WAIT7425 =>
                \$v7426\ := \$ram_lock\;
                if \$v7426\(0) = '1' then
                  state_var7460 := Q_WAIT7425;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr\ <= to_integer(unsigned(work.Int.sub(\$17105_w06555936_arg\(16 to 31), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7424;
                end if;
              when Q_WAIT7429 =>
                \$v7430\ := \$ram_lock\;
                if \$v7430\(0) = '1' then
                  state_var7460 := Q_WAIT7429;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(work.Int.add(
                                                          work.Int.add(
                                                          eclat_resize(\$17001\(64 to 94),16), X"000" & X"0"), X"000" & X"1")));
                  \$ram_write\ <= eclat_resize(work.Int.add(work.Int.add(
                                                            \$13911\(0 to 15), X"000" & X"3"), eclat_resize(\$16998_argument3\,16)),31) & eclat_true; \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7428;
                end if;
              when Q_WAIT7432 =>
                \$v7433\ := \$ram_lock\;
                if \$v7433\(0) = '1' then
                  state_var7460 := Q_WAIT7432;
                else
                  acquire(\$ram_lock\);
                  \$ram_ptr_write\ <= to_integer(unsigned(\$13911\(48 to 63)));
                  \$ram_write\ <= \$13911\(16 to 47); \$ram_write_request\ <= '1';
                  state_var7460 := PAUSE_SET7431;
                end if;
              when Q_WAIT7436 =>
                \$v7437\ := \$code_lock\;
                if \$v7437\(0) = '1' then
                  state_var7460 := Q_WAIT7436;
                else
                  acquire(\$code_lock\);
                  \$code_ptr\ <= to_integer(unsigned(\$13911\(0 to 15)));
                  state_var7460 := PAUSE_GET7435;
                end if;
              when Q_WAIT7440 =>
                \$v7441\ := \$code_lock\;
                if \$v7441\(0) = '1' then
                  state_var7460 := Q_WAIT7440;
                else
                  acquire(\$code_lock\);
                  \$code_ptr\ <= to_integer(unsigned(work.Int.add(\$13911\(0 to 15), X"000" & X"3")));
                  state_var7460 := PAUSE_GET7439;
                end if;
              when Q_WAIT7444 =>
                \$v7445\ := \$code_lock\;
                if \$v7445\(0) = '1' then
                  state_var7460 := Q_WAIT7444;
                else
                  acquire(\$code_lock\);
                  \$code_ptr\ <= to_integer(unsigned(work.Int.add(\$13911\(0 to 15), X"000" & X"2")));
                  state_var7460 := PAUSE_GET7443;
                end if;
              when Q_WAIT7448 =>
                \$v7449\ := \$code_lock\;
                if \$v7449\(0) = '1' then
                  state_var7460 := Q_WAIT7448;
                else
                  acquire(\$code_lock\);
                  \$code_ptr\ <= to_integer(unsigned(work.Int.add(\$13911\(0 to 15), X"000" & X"1")));
                  state_var7460 := PAUSE_GET7447;
                end if;
              when Q_WAIT7452 =>
                \$v7453\ := \$code_lock\;
                if \$v7453\(0) = '1' then
                  state_var7460 := Q_WAIT7452;
                else
                  acquire(\$code_lock\);
                  \$code_ptr\ <= to_integer(unsigned(\$13911\(0 to 15)));
                  state_var7460 := PAUSE_GET7451;
                end if;
              when IDLE6470 =>
                rdy6469 := eclat_false;
                \$13939\ := work.Print.print_string(clk,of_string("pc:"));
                \$13940\ := work.Int.print(clk,\$13911\(0 to 15));
                \$13941\ := work.Print.print_string(clk,of_string("|acc:"));
                \$13945\ := work.Int.print(clk,\$13911\(16 to 46));
                \$13946\ := work.Print.print_string(clk,of_string("<"));
                \$v7455\ := ""&\$13911\(47);
                if \$v7455\(0) = '1' then
                  \$17173\ := work.Print.print_string(clk,of_string("int"));
                  \$13950\ := work.Print.print_string(clk,of_string(">"));
                  \$13951\ := work.Print.print_string(clk,of_string("|sp:"));
                  \$13952\ := work.Int.print(clk,\$13911\(48 to 63));
                  \$13953\ := work.Print.print_string(clk,of_string("|env:"));
                  \$13957\ := work.Int.print(clk,\$13911\(64 to 94));
                  \$13958\ := work.Print.print_string(clk,of_string("<"));
                  \$v7454\ := ""&\$13911\(95);
                  if \$v7454\(0) = '1' then
                    \$17172\ := work.Print.print_string(clk,of_string("int"));
                    \$13962\ := work.Print.print_string(clk,of_string(">"));
                    \$13963\ := work.Print.print_newline(clk,eclat_unit);
                    \$13964\ := work.Assertion.ok(work.Int.lt(\$13911\(0 to 15), std_logic_vector(to_unsigned(code'length,16))));
                    \$v7453\ := \$code_lock\;
                    if \$v7453\(0) = '1' then
                      state_var7460 := Q_WAIT7452;
                    else
                      acquire(\$code_lock\);
                      \$code_ptr\ <= to_integer(unsigned(\$13911\(0 to 15)));
                      state_var7460 := PAUSE_GET7451;
                    end if;
                  else
                    \$17172\ := work.Print.print_string(clk,of_string("ptr"));
                    \$13962\ := work.Print.print_string(clk,of_string(">"));
                    \$13963\ := work.Print.print_newline(clk,eclat_unit);
                    \$13964\ := work.Assertion.ok(work.Int.lt(\$13911\(0 to 15), std_logic_vector(to_unsigned(code'length,16))));
                    \$v7453\ := \$code_lock\;
                    if \$v7453\(0) = '1' then
                      state_var7460 := Q_WAIT7452;
                    else
                      acquire(\$code_lock\);
                      \$code_ptr\ <= to_integer(unsigned(\$13911\(0 to 15)));
                      state_var7460 := PAUSE_GET7451;
                    end if;
                  end if;
                else
                  \$17173\ := work.Print.print_string(clk,of_string("ptr"));
                  \$13950\ := work.Print.print_string(clk,of_string(">"));
                  \$13951\ := work.Print.print_string(clk,of_string("|sp:"));
                  \$13952\ := work.Int.print(clk,\$13911\(48 to 63));
                  \$13953\ := work.Print.print_string(clk,of_string("|env:"));
                  \$13957\ := work.Int.print(clk,\$13911\(64 to 94));
                  \$13958\ := work.Print.print_string(clk,of_string("<"));
                  \$v7454\ := ""&\$13911\(95);
                  if \$v7454\(0) = '1' then
                    \$17172\ := work.Print.print_string(clk,of_string("int"));
                    \$13962\ := work.Print.print_string(clk,of_string(">"));
                    \$13963\ := work.Print.print_newline(clk,eclat_unit);
                    \$13964\ := work.Assertion.ok(work.Int.lt(\$13911\(0 to 15), std_logic_vector(to_unsigned(code'length,16))));
                    \$v7453\ := \$code_lock\;
                    if \$v7453\(0) = '1' then
                      state_var7460 := Q_WAIT7452;
                    else
                      acquire(\$code_lock\);
                      \$code_ptr\ <= to_integer(unsigned(\$13911\(0 to 15)));
                      state_var7460 := PAUSE_GET7451;
                    end if;
                  else
                    \$17172\ := work.Print.print_string(clk,of_string("ptr"));
                    \$13962\ := work.Print.print_string(clk,of_string(">"));
                    \$13963\ := work.Print.print_newline(clk,eclat_unit);
                    \$13964\ := work.Assertion.ok(work.Int.lt(\$13911\(0 to 15), std_logic_vector(to_unsigned(code'length,16))));
                    \$v7453\ := \$code_lock\;
                    if \$v7453\(0) = '1' then
                      state_var7460 := Q_WAIT7452;
                    else
                      acquire(\$code_lock\);
                      \$code_ptr\ <= to_integer(unsigned(\$13911\(0 to 15)));
                      state_var7460 := PAUSE_GET7451;
                    end if;
                  end if;
                end if;
              end case;
              
              if rdy6469(0) = '1' then
                
              else
                result6468 := \$13911\(0 to 121);
              end if;
              \$13917\ := result6468 & rdy6469;
              \$13911\ := \$13917\(0 to 121) & ""&\$13917\(122);
            end if;
            \$13897\ := \$13911\;
            \$12662\ := ""&\$13897\(120) & ""&\$13897\(122) & ""&\$12662\(2) & ""&\$13897\(121);
          end if;
          \$12539\ := \$12662\;
          \$v6111\ := ""&\$12539\(0);
          if \$v6111\(0) = '1' then
            \$12659\ := work.Print.print_string(clk,of_string("(cy="));
            \$12660\ := work.Int.print(clk,\$12538_cy\);
            \$12661\ := work.Print.print_string(clk,of_string(")"));
            \$12544\ := work.Print.print_newline(clk,eclat_unit);
            if \$v5876\(0) = '1' then
              
            else
              \$v5876\ := eclat_true;
              \$12657\ := eclat_false;
            end if;
            \$12657\ := eclat_if(""&\$12539\(0) & eclat_true & \$12657\);
            \$12545_x\ := \$12657\;
            if \$v5877\(0) = '1' then
              
            else
              \$v5877\ := eclat_true;
              \$12654\ := X"0000000" & X"0";
            end if;
            \$12654\ := eclat_if(work.Bool.lnot(\$12545_x\) & work.Int.add(
                                                              \$12654\, X"0000000" & X"1") & \$12654\);
            \$12546_dur\ := \$12654\;
            \$v6110\ := \$12545_x\;
            if \$v6110\(0) = '1' then
              \$12547\ := work.Int.print(clk,\$12546_dur\);
              \$v6109\ := \$12545_x\;
              if \$v6109\(0) = '1' then
                \$v6108\ := eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"3") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"2") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"1") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"0");
                case \$v6108\ is
                when "0000" =>
                  \$12558\ := "00000011";
                when "0001" =>
                  \$12558\ := "10011111";
                when "0010" =>
                  \$12558\ := "00100101";
                when "0011" =>
                  \$12558\ := "00001101";
                when "0100" =>
                  \$12558\ := "10011001";
                when "0101" =>
                  \$12558\ := "01001001";
                when "0110" =>
                  \$12558\ := "01000001";
                when "0111" =>
                  \$12558\ := "00011111";
                when "1000" =>
                  \$12558\ := "00000001";
                when "1001" =>
                  \$12558\ := "00001001";
                when "1010" =>
                  \$12558\ := "00010001";
                when "1011" =>
                  \$12558\ := "11000001";
                when "1100" =>
                  \$12558\ := "01100011";
                when "1101" =>
                  \$12558\ := "10000101";
                when "1110" =>
                  \$12558\ := "01100001";
                when "1111" =>
                  \$12558\ := "01110001";
                when others =>
                  \$12558\ := "11100011";
                end case;
                \$v6107\ := eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"7") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"6") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"5") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"4");
                case \$v6107\ is
                when "0000" =>
                  \$12559\ := "00000011";
                when "0001" =>
                  \$12559\ := "10011111";
                when "0010" =>
                  \$12559\ := "00100101";
                when "0011" =>
                  \$12559\ := "00001101";
                when "0100" =>
                  \$12559\ := "10011001";
                when "0101" =>
                  \$12559\ := "01001001";
                when "0110" =>
                  \$12559\ := "01000001";
                when "0111" =>
                  \$12559\ := "00011111";
                when "1000" =>
                  \$12559\ := "00000001";
                when "1001" =>
                  \$12559\ := "00001001";
                when "1010" =>
                  \$12559\ := "00010001";
                when "1011" =>
                  \$12559\ := "11000001";
                when "1100" =>
                  \$12559\ := "01100011";
                when "1101" =>
                  \$12559\ := "10000101";
                when "1110" =>
                  \$12559\ := "01100001";
                when "1111" =>
                  \$12559\ := "01110001";
                when others =>
                  \$12559\ := "11100011";
                end case;
                \$v6106\ := eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"b") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"a") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"9") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"8");
                case \$v6106\ is
                when "0000" =>
                  \$12560\ := "00000011";
                when "0001" =>
                  \$12560\ := "10011111";
                when "0010" =>
                  \$12560\ := "00100101";
                when "0011" =>
                  \$12560\ := "00001101";
                when "0100" =>
                  \$12560\ := "10011001";
                when "0101" =>
                  \$12560\ := "01001001";
                when "0110" =>
                  \$12560\ := "01000001";
                when "0111" =>
                  \$12560\ := "00011111";
                when "1000" =>
                  \$12560\ := "00000001";
                when "1001" =>
                  \$12560\ := "00001001";
                when "1010" =>
                  \$12560\ := "00010001";
                when "1011" =>
                  \$12560\ := "11000001";
                when "1100" =>
                  \$12560\ := "01100011";
                when "1101" =>
                  \$12560\ := "10000101";
                when "1110" =>
                  \$12560\ := "01100001";
                when "1111" =>
                  \$12560\ := "01110001";
                when others =>
                  \$12560\ := "11100011";
                end case;
                \$v6105\ := eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"f") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"e") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"d") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"c");
                case \$v6105\ is
                when "0000" =>
                  \$12561\ := "00000011";
                when "0001" =>
                  \$12561\ := "10011111";
                when "0010" =>
                  \$12561\ := "00100101";
                when "0011" =>
                  \$12561\ := "00001101";
                when "0100" =>
                  \$12561\ := "10011001";
                when "0101" =>
                  \$12561\ := "01001001";
                when "0110" =>
                  \$12561\ := "01000001";
                when "0111" =>
                  \$12561\ := "00011111";
                when "1000" =>
                  \$12561\ := "00000001";
                when "1001" =>
                  \$12561\ := "00001001";
                when "1010" =>
                  \$12561\ := "00010001";
                when "1011" =>
                  \$12561\ := "11000001";
                when "1100" =>
                  \$12561\ := "01100011";
                when "1101" =>
                  \$12561\ := "10000101";
                when "1110" =>
                  \$12561\ := "01100001";
                when "1111" =>
                  \$12561\ := "01110001";
                when others =>
                  \$12561\ := "11100011";
                end case;
                \$v6104\ := eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"13") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"12") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"11") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"10");
                case \$v6104\ is
                when "0000" =>
                  \$12562\ := "00000011";
                when "0001" =>
                  \$12562\ := "10011111";
                when "0010" =>
                  \$12562\ := "00100101";
                when "0011" =>
                  \$12562\ := "00001101";
                when "0100" =>
                  \$12562\ := "10011001";
                when "0101" =>
                  \$12562\ := "01001001";
                when "0110" =>
                  \$12562\ := "01000001";
                when "0111" =>
                  \$12562\ := "00011111";
                when "1000" =>
                  \$12562\ := "00000001";
                when "1001" =>
                  \$12562\ := "00001001";
                when "1010" =>
                  \$12562\ := "00010001";
                when "1011" =>
                  \$12562\ := "11000001";
                when "1100" =>
                  \$12562\ := "01100011";
                when "1101" =>
                  \$12562\ := "10000101";
                when "1110" =>
                  \$12562\ := "01100001";
                when "1111" =>
                  \$12562\ := "01110001";
                when others =>
                  \$12562\ := "11100011";
                end case;
                \$v6103\ := eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"17") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"16") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"15") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"14");
                case \$v6103\ is
                when "0000" =>
                  \$12563\ := "00000011";
                when "0001" =>
                  \$12563\ := "10011111";
                when "0010" =>
                  \$12563\ := "00100101";
                when "0011" =>
                  \$12563\ := "00001101";
                when "0100" =>
                  \$12563\ := "10011001";
                when "0101" =>
                  \$12563\ := "01001001";
                when "0110" =>
                  \$12563\ := "01000001";
                when "0111" =>
                  \$12563\ := "00011111";
                when "1000" =>
                  \$12563\ := "00000001";
                when "1001" =>
                  \$12563\ := "00001001";
                when "1010" =>
                  \$12563\ := "00010001";
                when "1011" =>
                  \$12563\ := "11000001";
                when "1100" =>
                  \$12563\ := "01100011";
                when "1101" =>
                  \$12563\ := "10000101";
                when "1110" =>
                  \$12563\ := "01100001";
                when "1111" =>
                  \$12563\ := "01110001";
                when others =>
                  \$12563\ := "11100011";
                end case;
                \$12548_dis\ := \$12558\ & \$12559\ & \$12560\ & \$12561\ & \$12562\ & \$12563\;
              else
                \$12548_dis\ := "00000011" & "00000011" & "00000011" & "00000011" & "00000011" & "00000011";
              end if;
              if \$v5878\(0) = '1' then
                
              else
                \$v5878\ := eclat_true;
                \$12553\ := X"0000000" & X"0";
              end if;
              \$12553\ := eclat_if(work.Int.eq(\$12553\, work.Int.add(
                                                         X"00" & X"989680", X"00" & X"989680")) & X"0000000" & X"0" & 
                          work.Int.add(\$12553\, X"0000000" & X"1"));
              \$12549\ := \$12553\;
              result5939 := ""&\$12539\(0) & work.Bool.lnot(""&\$12539\(1)) & 
              work.Int.gt(\$12549\, X"00" & X"989680") & ""&\$12539\(3) & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & \$12548_dis\;
              rdy5940 := eclat_true;
              state := IDLE5941;
            else
              \$12547\ := eclat_unit;
              \$v6109\ := \$12545_x\;
              if \$v6109\(0) = '1' then
                \$v6108\ := eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"3") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"2") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"1") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"0");
                case \$v6108\ is
                when "0000" =>
                  \$12558\ := "00000011";
                when "0001" =>
                  \$12558\ := "10011111";
                when "0010" =>
                  \$12558\ := "00100101";
                when "0011" =>
                  \$12558\ := "00001101";
                when "0100" =>
                  \$12558\ := "10011001";
                when "0101" =>
                  \$12558\ := "01001001";
                when "0110" =>
                  \$12558\ := "01000001";
                when "0111" =>
                  \$12558\ := "00011111";
                when "1000" =>
                  \$12558\ := "00000001";
                when "1001" =>
                  \$12558\ := "00001001";
                when "1010" =>
                  \$12558\ := "00010001";
                when "1011" =>
                  \$12558\ := "11000001";
                when "1100" =>
                  \$12558\ := "01100011";
                when "1101" =>
                  \$12558\ := "10000101";
                when "1110" =>
                  \$12558\ := "01100001";
                when "1111" =>
                  \$12558\ := "01110001";
                when others =>
                  \$12558\ := "11100011";
                end case;
                \$v6107\ := eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"7") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"6") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"5") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"4");
                case \$v6107\ is
                when "0000" =>
                  \$12559\ := "00000011";
                when "0001" =>
                  \$12559\ := "10011111";
                when "0010" =>
                  \$12559\ := "00100101";
                when "0011" =>
                  \$12559\ := "00001101";
                when "0100" =>
                  \$12559\ := "10011001";
                when "0101" =>
                  \$12559\ := "01001001";
                when "0110" =>
                  \$12559\ := "01000001";
                when "0111" =>
                  \$12559\ := "00011111";
                when "1000" =>
                  \$12559\ := "00000001";
                when "1001" =>
                  \$12559\ := "00001001";
                when "1010" =>
                  \$12559\ := "00010001";
                when "1011" =>
                  \$12559\ := "11000001";
                when "1100" =>
                  \$12559\ := "01100011";
                when "1101" =>
                  \$12559\ := "10000101";
                when "1110" =>
                  \$12559\ := "01100001";
                when "1111" =>
                  \$12559\ := "01110001";
                when others =>
                  \$12559\ := "11100011";
                end case;
                \$v6106\ := eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"b") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"a") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"9") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"8");
                case \$v6106\ is
                when "0000" =>
                  \$12560\ := "00000011";
                when "0001" =>
                  \$12560\ := "10011111";
                when "0010" =>
                  \$12560\ := "00100101";
                when "0011" =>
                  \$12560\ := "00001101";
                when "0100" =>
                  \$12560\ := "10011001";
                when "0101" =>
                  \$12560\ := "01001001";
                when "0110" =>
                  \$12560\ := "01000001";
                when "0111" =>
                  \$12560\ := "00011111";
                when "1000" =>
                  \$12560\ := "00000001";
                when "1001" =>
                  \$12560\ := "00001001";
                when "1010" =>
                  \$12560\ := "00010001";
                when "1011" =>
                  \$12560\ := "11000001";
                when "1100" =>
                  \$12560\ := "01100011";
                when "1101" =>
                  \$12560\ := "10000101";
                when "1110" =>
                  \$12560\ := "01100001";
                when "1111" =>
                  \$12560\ := "01110001";
                when others =>
                  \$12560\ := "11100011";
                end case;
                \$v6105\ := eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"f") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"e") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"d") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"c");
                case \$v6105\ is
                when "0000" =>
                  \$12561\ := "00000011";
                when "0001" =>
                  \$12561\ := "10011111";
                when "0010" =>
                  \$12561\ := "00100101";
                when "0011" =>
                  \$12561\ := "00001101";
                when "0100" =>
                  \$12561\ := "10011001";
                when "0101" =>
                  \$12561\ := "01001001";
                when "0110" =>
                  \$12561\ := "01000001";
                when "0111" =>
                  \$12561\ := "00011111";
                when "1000" =>
                  \$12561\ := "00000001";
                when "1001" =>
                  \$12561\ := "00001001";
                when "1010" =>
                  \$12561\ := "00010001";
                when "1011" =>
                  \$12561\ := "11000001";
                when "1100" =>
                  \$12561\ := "01100011";
                when "1101" =>
                  \$12561\ := "10000101";
                when "1110" =>
                  \$12561\ := "01100001";
                when "1111" =>
                  \$12561\ := "01110001";
                when others =>
                  \$12561\ := "11100011";
                end case;
                \$v6104\ := eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"13") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"12") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"11") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"10");
                case \$v6104\ is
                when "0000" =>
                  \$12562\ := "00000011";
                when "0001" =>
                  \$12562\ := "10011111";
                when "0010" =>
                  \$12562\ := "00100101";
                when "0011" =>
                  \$12562\ := "00001101";
                when "0100" =>
                  \$12562\ := "10011001";
                when "0101" =>
                  \$12562\ := "01001001";
                when "0110" =>
                  \$12562\ := "01000001";
                when "0111" =>
                  \$12562\ := "00011111";
                when "1000" =>
                  \$12562\ := "00000001";
                when "1001" =>
                  \$12562\ := "00001001";
                when "1010" =>
                  \$12562\ := "00010001";
                when "1011" =>
                  \$12562\ := "11000001";
                when "1100" =>
                  \$12562\ := "01100011";
                when "1101" =>
                  \$12562\ := "10000101";
                when "1110" =>
                  \$12562\ := "01100001";
                when "1111" =>
                  \$12562\ := "01110001";
                when others =>
                  \$12562\ := "11100011";
                end case;
                \$v6103\ := eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"17") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"16") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"15") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"14");
                case \$v6103\ is
                when "0000" =>
                  \$12563\ := "00000011";
                when "0001" =>
                  \$12563\ := "10011111";
                when "0010" =>
                  \$12563\ := "00100101";
                when "0011" =>
                  \$12563\ := "00001101";
                when "0100" =>
                  \$12563\ := "10011001";
                when "0101" =>
                  \$12563\ := "01001001";
                when "0110" =>
                  \$12563\ := "01000001";
                when "0111" =>
                  \$12563\ := "00011111";
                when "1000" =>
                  \$12563\ := "00000001";
                when "1001" =>
                  \$12563\ := "00001001";
                when "1010" =>
                  \$12563\ := "00010001";
                when "1011" =>
                  \$12563\ := "11000001";
                when "1100" =>
                  \$12563\ := "01100011";
                when "1101" =>
                  \$12563\ := "10000101";
                when "1110" =>
                  \$12563\ := "01100001";
                when "1111" =>
                  \$12563\ := "01110001";
                when others =>
                  \$12563\ := "11100011";
                end case;
                \$12548_dis\ := \$12558\ & \$12559\ & \$12560\ & \$12561\ & \$12562\ & \$12563\;
              else
                \$12548_dis\ := "00000011" & "00000011" & "00000011" & "00000011" & "00000011" & "00000011";
              end if;
              if \$v5878\(0) = '1' then
                
              else
                \$v5878\ := eclat_true;
                \$12553\ := X"0000000" & X"0";
              end if;
              \$12553\ := eclat_if(work.Int.eq(\$12553\, work.Int.add(
                                                         X"00" & X"989680", X"00" & X"989680")) & X"0000000" & X"0" & 
                          work.Int.add(\$12553\, X"0000000" & X"1"));
              \$12549\ := \$12553\;
              result5939 := ""&\$12539\(0) & work.Bool.lnot(""&\$12539\(1)) & 
              work.Int.gt(\$12549\, X"00" & X"989680") & ""&\$12539\(3) & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & \$12548_dis\;
              rdy5940 := eclat_true;
              state := IDLE5941;
            end if;
          else
            \$12544\ := eclat_unit;
            if \$v5876\(0) = '1' then
              
            else
              \$v5876\ := eclat_true;
              \$12657\ := eclat_false;
            end if;
            \$12657\ := eclat_if(""&\$12539\(0) & eclat_true & \$12657\);
            \$12545_x\ := \$12657\;
            if \$v5877\(0) = '1' then
              
            else
              \$v5877\ := eclat_true;
              \$12654\ := X"0000000" & X"0";
            end if;
            \$12654\ := eclat_if(work.Bool.lnot(\$12545_x\) & work.Int.add(
                                                              \$12654\, X"0000000" & X"1") & \$12654\);
            \$12546_dur\ := \$12654\;
            \$v6110\ := \$12545_x\;
            if \$v6110\(0) = '1' then
              \$12547\ := work.Int.print(clk,\$12546_dur\);
              \$v6109\ := \$12545_x\;
              if \$v6109\(0) = '1' then
                \$v6108\ := eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"3") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"2") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"1") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"0");
                case \$v6108\ is
                when "0000" =>
                  \$12558\ := "00000011";
                when "0001" =>
                  \$12558\ := "10011111";
                when "0010" =>
                  \$12558\ := "00100101";
                when "0011" =>
                  \$12558\ := "00001101";
                when "0100" =>
                  \$12558\ := "10011001";
                when "0101" =>
                  \$12558\ := "01001001";
                when "0110" =>
                  \$12558\ := "01000001";
                when "0111" =>
                  \$12558\ := "00011111";
                when "1000" =>
                  \$12558\ := "00000001";
                when "1001" =>
                  \$12558\ := "00001001";
                when "1010" =>
                  \$12558\ := "00010001";
                when "1011" =>
                  \$12558\ := "11000001";
                when "1100" =>
                  \$12558\ := "01100011";
                when "1101" =>
                  \$12558\ := "10000101";
                when "1110" =>
                  \$12558\ := "01100001";
                when "1111" =>
                  \$12558\ := "01110001";
                when others =>
                  \$12558\ := "11100011";
                end case;
                \$v6107\ := eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"7") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"6") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"5") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"4");
                case \$v6107\ is
                when "0000" =>
                  \$12559\ := "00000011";
                when "0001" =>
                  \$12559\ := "10011111";
                when "0010" =>
                  \$12559\ := "00100101";
                when "0011" =>
                  \$12559\ := "00001101";
                when "0100" =>
                  \$12559\ := "10011001";
                when "0101" =>
                  \$12559\ := "01001001";
                when "0110" =>
                  \$12559\ := "01000001";
                when "0111" =>
                  \$12559\ := "00011111";
                when "1000" =>
                  \$12559\ := "00000001";
                when "1001" =>
                  \$12559\ := "00001001";
                when "1010" =>
                  \$12559\ := "00010001";
                when "1011" =>
                  \$12559\ := "11000001";
                when "1100" =>
                  \$12559\ := "01100011";
                when "1101" =>
                  \$12559\ := "10000101";
                when "1110" =>
                  \$12559\ := "01100001";
                when "1111" =>
                  \$12559\ := "01110001";
                when others =>
                  \$12559\ := "11100011";
                end case;
                \$v6106\ := eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"b") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"a") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"9") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"8");
                case \$v6106\ is
                when "0000" =>
                  \$12560\ := "00000011";
                when "0001" =>
                  \$12560\ := "10011111";
                when "0010" =>
                  \$12560\ := "00100101";
                when "0011" =>
                  \$12560\ := "00001101";
                when "0100" =>
                  \$12560\ := "10011001";
                when "0101" =>
                  \$12560\ := "01001001";
                when "0110" =>
                  \$12560\ := "01000001";
                when "0111" =>
                  \$12560\ := "00011111";
                when "1000" =>
                  \$12560\ := "00000001";
                when "1001" =>
                  \$12560\ := "00001001";
                when "1010" =>
                  \$12560\ := "00010001";
                when "1011" =>
                  \$12560\ := "11000001";
                when "1100" =>
                  \$12560\ := "01100011";
                when "1101" =>
                  \$12560\ := "10000101";
                when "1110" =>
                  \$12560\ := "01100001";
                when "1111" =>
                  \$12560\ := "01110001";
                when others =>
                  \$12560\ := "11100011";
                end case;
                \$v6105\ := eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"f") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"e") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"d") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"c");
                case \$v6105\ is
                when "0000" =>
                  \$12561\ := "00000011";
                when "0001" =>
                  \$12561\ := "10011111";
                when "0010" =>
                  \$12561\ := "00100101";
                when "0011" =>
                  \$12561\ := "00001101";
                when "0100" =>
                  \$12561\ := "10011001";
                when "0101" =>
                  \$12561\ := "01001001";
                when "0110" =>
                  \$12561\ := "01000001";
                when "0111" =>
                  \$12561\ := "00011111";
                when "1000" =>
                  \$12561\ := "00000001";
                when "1001" =>
                  \$12561\ := "00001001";
                when "1010" =>
                  \$12561\ := "00010001";
                when "1011" =>
                  \$12561\ := "11000001";
                when "1100" =>
                  \$12561\ := "01100011";
                when "1101" =>
                  \$12561\ := "10000101";
                when "1110" =>
                  \$12561\ := "01100001";
                when "1111" =>
                  \$12561\ := "01110001";
                when others =>
                  \$12561\ := "11100011";
                end case;
                \$v6104\ := eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"13") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"12") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"11") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"10");
                case \$v6104\ is
                when "0000" =>
                  \$12562\ := "00000011";
                when "0001" =>
                  \$12562\ := "10011111";
                when "0010" =>
                  \$12562\ := "00100101";
                when "0011" =>
                  \$12562\ := "00001101";
                when "0100" =>
                  \$12562\ := "10011001";
                when "0101" =>
                  \$12562\ := "01001001";
                when "0110" =>
                  \$12562\ := "01000001";
                when "0111" =>
                  \$12562\ := "00011111";
                when "1000" =>
                  \$12562\ := "00000001";
                when "1001" =>
                  \$12562\ := "00001001";
                when "1010" =>
                  \$12562\ := "00010001";
                when "1011" =>
                  \$12562\ := "11000001";
                when "1100" =>
                  \$12562\ := "01100011";
                when "1101" =>
                  \$12562\ := "10000101";
                when "1110" =>
                  \$12562\ := "01100001";
                when "1111" =>
                  \$12562\ := "01110001";
                when others =>
                  \$12562\ := "11100011";
                end case;
                \$v6103\ := eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"17") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"16") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"15") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"14");
                case \$v6103\ is
                when "0000" =>
                  \$12563\ := "00000011";
                when "0001" =>
                  \$12563\ := "10011111";
                when "0010" =>
                  \$12563\ := "00100101";
                when "0011" =>
                  \$12563\ := "00001101";
                when "0100" =>
                  \$12563\ := "10011001";
                when "0101" =>
                  \$12563\ := "01001001";
                when "0110" =>
                  \$12563\ := "01000001";
                when "0111" =>
                  \$12563\ := "00011111";
                when "1000" =>
                  \$12563\ := "00000001";
                when "1001" =>
                  \$12563\ := "00001001";
                when "1010" =>
                  \$12563\ := "00010001";
                when "1011" =>
                  \$12563\ := "11000001";
                when "1100" =>
                  \$12563\ := "01100011";
                when "1101" =>
                  \$12563\ := "10000101";
                when "1110" =>
                  \$12563\ := "01100001";
                when "1111" =>
                  \$12563\ := "01110001";
                when others =>
                  \$12563\ := "11100011";
                end case;
                \$12548_dis\ := \$12558\ & \$12559\ & \$12560\ & \$12561\ & \$12562\ & \$12563\;
              else
                \$12548_dis\ := "00000011" & "00000011" & "00000011" & "00000011" & "00000011" & "00000011";
              end if;
              if \$v5878\(0) = '1' then
                
              else
                \$v5878\ := eclat_true;
                \$12553\ := X"0000000" & X"0";
              end if;
              \$12553\ := eclat_if(work.Int.eq(\$12553\, work.Int.add(
                                                         X"00" & X"989680", X"00" & X"989680")) & X"0000000" & X"0" & 
                          work.Int.add(\$12553\, X"0000000" & X"1"));
              \$12549\ := \$12553\;
              result5939 := ""&\$12539\(0) & work.Bool.lnot(""&\$12539\(1)) & 
              work.Int.gt(\$12549\, X"00" & X"989680") & ""&\$12539\(3) & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & \$12548_dis\;
              rdy5940 := eclat_true;
              state := IDLE5941;
            else
              \$12547\ := eclat_unit;
              \$v6109\ := \$12545_x\;
              if \$v6109\(0) = '1' then
                \$v6108\ := eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"3") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"2") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"1") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"0");
                case \$v6108\ is
                when "0000" =>
                  \$12558\ := "00000011";
                when "0001" =>
                  \$12558\ := "10011111";
                when "0010" =>
                  \$12558\ := "00100101";
                when "0011" =>
                  \$12558\ := "00001101";
                when "0100" =>
                  \$12558\ := "10011001";
                when "0101" =>
                  \$12558\ := "01001001";
                when "0110" =>
                  \$12558\ := "01000001";
                when "0111" =>
                  \$12558\ := "00011111";
                when "1000" =>
                  \$12558\ := "00000001";
                when "1001" =>
                  \$12558\ := "00001001";
                when "1010" =>
                  \$12558\ := "00010001";
                when "1011" =>
                  \$12558\ := "11000001";
                when "1100" =>
                  \$12558\ := "01100011";
                when "1101" =>
                  \$12558\ := "10000101";
                when "1110" =>
                  \$12558\ := "01100001";
                when "1111" =>
                  \$12558\ := "01110001";
                when others =>
                  \$12558\ := "11100011";
                end case;
                \$v6107\ := eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"7") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"6") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"5") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"4");
                case \$v6107\ is
                when "0000" =>
                  \$12559\ := "00000011";
                when "0001" =>
                  \$12559\ := "10011111";
                when "0010" =>
                  \$12559\ := "00100101";
                when "0011" =>
                  \$12559\ := "00001101";
                when "0100" =>
                  \$12559\ := "10011001";
                when "0101" =>
                  \$12559\ := "01001001";
                when "0110" =>
                  \$12559\ := "01000001";
                when "0111" =>
                  \$12559\ := "00011111";
                when "1000" =>
                  \$12559\ := "00000001";
                when "1001" =>
                  \$12559\ := "00001001";
                when "1010" =>
                  \$12559\ := "00010001";
                when "1011" =>
                  \$12559\ := "11000001";
                when "1100" =>
                  \$12559\ := "01100011";
                when "1101" =>
                  \$12559\ := "10000101";
                when "1110" =>
                  \$12559\ := "01100001";
                when "1111" =>
                  \$12559\ := "01110001";
                when others =>
                  \$12559\ := "11100011";
                end case;
                \$v6106\ := eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"b") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"a") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"9") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"8");
                case \$v6106\ is
                when "0000" =>
                  \$12560\ := "00000011";
                when "0001" =>
                  \$12560\ := "10011111";
                when "0010" =>
                  \$12560\ := "00100101";
                when "0011" =>
                  \$12560\ := "00001101";
                when "0100" =>
                  \$12560\ := "10011001";
                when "0101" =>
                  \$12560\ := "01001001";
                when "0110" =>
                  \$12560\ := "01000001";
                when "0111" =>
                  \$12560\ := "00011111";
                when "1000" =>
                  \$12560\ := "00000001";
                when "1001" =>
                  \$12560\ := "00001001";
                when "1010" =>
                  \$12560\ := "00010001";
                when "1011" =>
                  \$12560\ := "11000001";
                when "1100" =>
                  \$12560\ := "01100011";
                when "1101" =>
                  \$12560\ := "10000101";
                when "1110" =>
                  \$12560\ := "01100001";
                when "1111" =>
                  \$12560\ := "01110001";
                when others =>
                  \$12560\ := "11100011";
                end case;
                \$v6105\ := eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"f") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"e") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"d") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"0000000" & X"c");
                case \$v6105\ is
                when "0000" =>
                  \$12561\ := "00000011";
                when "0001" =>
                  \$12561\ := "10011111";
                when "0010" =>
                  \$12561\ := "00100101";
                when "0011" =>
                  \$12561\ := "00001101";
                when "0100" =>
                  \$12561\ := "10011001";
                when "0101" =>
                  \$12561\ := "01001001";
                when "0110" =>
                  \$12561\ := "01000001";
                when "0111" =>
                  \$12561\ := "00011111";
                when "1000" =>
                  \$12561\ := "00000001";
                when "1001" =>
                  \$12561\ := "00001001";
                when "1010" =>
                  \$12561\ := "00010001";
                when "1011" =>
                  \$12561\ := "11000001";
                when "1100" =>
                  \$12561\ := "01100011";
                when "1101" =>
                  \$12561\ := "10000101";
                when "1110" =>
                  \$12561\ := "01100001";
                when "1111" =>
                  \$12561\ := "01110001";
                when others =>
                  \$12561\ := "11100011";
                end case;
                \$v6104\ := eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"13") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"12") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"11") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"10");
                case \$v6104\ is
                when "0000" =>
                  \$12562\ := "00000011";
                when "0001" =>
                  \$12562\ := "10011111";
                when "0010" =>
                  \$12562\ := "00100101";
                when "0011" =>
                  \$12562\ := "00001101";
                when "0100" =>
                  \$12562\ := "10011001";
                when "0101" =>
                  \$12562\ := "01001001";
                when "0110" =>
                  \$12562\ := "01000001";
                when "0111" =>
                  \$12562\ := "00011111";
                when "1000" =>
                  \$12562\ := "00000001";
                when "1001" =>
                  \$12562\ := "00001001";
                when "1010" =>
                  \$12562\ := "00010001";
                when "1011" =>
                  \$12562\ := "11000001";
                when "1100" =>
                  \$12562\ := "01100011";
                when "1101" =>
                  \$12562\ := "10000101";
                when "1110" =>
                  \$12562\ := "01100001";
                when "1111" =>
                  \$12562\ := "01110001";
                when others =>
                  \$12562\ := "11100011";
                end case;
                \$v6103\ := eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"17") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"16") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"15") & eclat_getBit(eclat_resize(\$12546_dur\,25) & X"000000" & X"14");
                case \$v6103\ is
                when "0000" =>
                  \$12563\ := "00000011";
                when "0001" =>
                  \$12563\ := "10011111";
                when "0010" =>
                  \$12563\ := "00100101";
                when "0011" =>
                  \$12563\ := "00001101";
                when "0100" =>
                  \$12563\ := "10011001";
                when "0101" =>
                  \$12563\ := "01001001";
                when "0110" =>
                  \$12563\ := "01000001";
                when "0111" =>
                  \$12563\ := "00011111";
                when "1000" =>
                  \$12563\ := "00000001";
                when "1001" =>
                  \$12563\ := "00001001";
                when "1010" =>
                  \$12563\ := "00010001";
                when "1011" =>
                  \$12563\ := "11000001";
                when "1100" =>
                  \$12563\ := "01100011";
                when "1101" =>
                  \$12563\ := "10000101";
                when "1110" =>
                  \$12563\ := "01100001";
                when "1111" =>
                  \$12563\ := "01110001";
                when others =>
                  \$12563\ := "11100011";
                end case;
                \$12548_dis\ := \$12558\ & \$12559\ & \$12560\ & \$12561\ & \$12562\ & \$12563\;
              else
                \$12548_dis\ := "00000011" & "00000011" & "00000011" & "00000011" & "00000011" & "00000011";
              end if;
              if \$v5878\(0) = '1' then
                
              else
                \$v5878\ := eclat_true;
                \$12553\ := X"0000000" & X"0";
              end if;
              \$12553\ := eclat_if(work.Int.eq(\$12553\, work.Int.add(
                                                         X"00" & X"989680", X"00" & X"989680")) & X"0000000" & X"0" & 
                          work.Int.add(\$12553\, X"0000000" & X"1"));
              \$12549\ := \$12553\;
              result5939 := ""&\$12539\(0) & work.Bool.lnot(""&\$12539\(1)) & 
              work.Int.gt(\$12549\, X"00" & X"989680") & ""&\$12539\(3) & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & \$12548_dis\;
              rdy5940 := eclat_true;
              state := IDLE5941;
            end if;
          end if;
        end if;
      end case;
      \state%next\ <= state;
      \state_var7464%next\ <= state_var7464;
      \state_var7463%next\ <= state_var7463;
      \state_var7462%next\ <= state_var7462;
      \state_var7461%next\ <= state_var7461;
      \state_var7460%next\ <= state_var7460;
      \$12559%next\ <= \$12559\;
      \$14060%next\ <= \$14060\;
      \$v6454%next\ <= \$v6454\;
      \$14516_v%next\ <= \$14516_v\;
      \$15069_modulo6685895_arg%next\ <= \$15069_modulo6685895_arg\;
      \$18421%next\ <= \$18421\;
      \$v6570%next\ <= \$v6570\;
      \$14564_binop_int6435900_arg%next\ <= \$14564_binop_int6435900_arg\;
      \$17813%next\ <= \$17813\;
      \$v6841%next\ <= \$v6841\;
      \$14666_r%next\ <= \$14666_r\;
      \$v7022%next\ <= \$v7022\;
      \$14589_modulo6685895_result%next\ <= \$14589_modulo6685895_result\;
      \$13392%next\ <= \$13392\;
      \$18996%next\ <= \$18996\;
      \$12673_rdy%next\ <= \$12673_rdy\;
      \$v6130%next\ <= \$v6130\;
      \$v7263%next\ <= \$v7263\;
      \$14917_modulo6685888_arg%next\ <= \$14917_modulo6685888_arg\;
      \$v6197%next\ <= \$v6197\;
      \$19272%next\ <= \$19272\;
      \$v7123%next\ <= \$v7123\;
      \$v6642%next\ <= \$v6642\;
      \$18729%next\ <= \$18729\;
      \$18192%next\ <= \$18192\;
      \$13670%next\ <= \$13670\;
      \$v6127%next\ <= \$v6127\;
      \$15675_v%next\ <= \$15675_v\;
      \$15077_modulo6685888_result%next\ <= \$15077_modulo6685888_result\;
      \$v6725%next\ <= \$v6725\;
      \$16182%next\ <= \$16182\;
      \$14052_v%next\ <= \$14052_v\;
      \$18354%next\ <= \$18354\;
      \$14749_modulo6685895_result%next\ <= \$14749_modulo6685895_result\;
      \$v6451%next\ <= \$v6451\;
      \$12545_x%next\ <= \$12545_x\;
      \$v7062%next\ <= \$v7062\;
      \$17496_next%next\ <= \$17496_next\;
      \$12852%next\ <= \$12852\;
      \$13503%next\ <= \$13503\;
      \$v6473%next\ <= \$v6473\;
      \$15531_binop_int6435913_arg%next\ <= \$15531_binop_int6435913_arg\;
      \$17887%next\ <= \$17887\;
      \$18997%next\ <= \$18997\;
      \$18835%next\ <= \$18835\;
      \$v6567%next\ <= \$v6567\;
      \$v7313%next\ <= \$v7313\;
      \$14724_binop_int6435902_result%next\ <= \$14724_binop_int6435902_result\;
      \$12699%next\ <= \$12699\;
      \$v7125%next\ <= \$v7125\;
      \$14989_modulo6685895_arg%next\ <= \$14989_modulo6685895_arg\;
      \$13090%next\ <= \$13090\;
      \$19003%next\ <= \$19003\;
      \$12522_wait662_arg%next\ <= \$12522_wait662_arg\;
      \$16811_compare6445898_arg%next\ <= \$16811_compare6445898_arg\;
      \$17893%next\ <= \$17893\;
      \$15661_binop_compare6455917_arg%next\ <= \$15661_binop_compare6455917_arg\;
      \$14126%next\ <= \$14126\;
      \$v7437%next\ <= \$v7437\;
      \$17570%next\ <= \$17570\;
      \$16453_v%next\ <= \$16453_v\;
      \$17676%next\ <= \$17676\;
      \$18121%next\ <= \$18121\;
      \$v7222%next\ <= \$v7222\;
      \$v6512%next\ <= \$v6512\;
      \$13308%next\ <= \$13308\;
      \$17018_w36575938_arg%next\ <= \$17018_w36575938_arg\;
      \$v6206%next\ <= \$v6206\;
      \$15484_modulo6685888_result%next\ <= \$15484_modulo6685888_result\;
      \$v7170%next\ <= \$v7170\;
      \$15614_forever6705914_arg%next\ <= \$15614_forever6705914_arg\;
      \$16858_compbranch6505932_arg%next\ <= \$16858_compbranch6505932_arg\;
      \$v7236%next\ <= \$v7236\;
      \$v7153%next\ <= \$v7153\;
      \$16893_compbranch6505933_id%next\ <= \$16893_compbranch6505933_id\;
      \$14597_modulo6685888_arg%next\ <= \$14597_modulo6685888_arg\;
      \$16141%next\ <= \$16141\;
      \$v6105%next\ <= \$v6105\;
      \$v7446%next\ <= \$v7446\;
      \$13156%next\ <= \$13156\;
      \$v6575%next\ <= \$v6575\;
      \$19138%next\ <= \$19138\;
      \$16178_v%next\ <= \$16178_v\;
      \$13945%next\ <= \$13945\;
      \$v7094%next\ <= \$v7094\;
      \$v6391%next\ <= \$v6391\;
      \$18838%next\ <= \$18838\;
      \$13824%next\ <= \$13824\;
      \$v6959%next\ <= \$v6959\;
      \$13531%next\ <= \$13531\;
      \$16788_compbranch6505930_arg%next\ <= \$16788_compbranch6505930_arg\;
      \$17971%next\ <= \$17971\;
      \$v6348%next\ <= \$v6348\;
      \$17121%next\ <= \$17121\;
      \$16752_fill6545929_arg%next\ <= \$16752_fill6545929_arg\;
      \$v6382%next\ <= \$v6382\;
      \$12853_forever6705887_arg%next\ <= \$12853_forever6705887_arg\;
      \$v7251%next\ <= \$v7251\;
      \$15769_binop_compare6455920_arg%next\ <= \$15769_binop_compare6455920_arg\;
      \$17494%next\ <= \$17494\;
      \$v6385%next\ <= \$v6385\;
      \$14326%next\ <= \$14326\;
      \$v6240%next\ <= \$v6240\;
      \$19080_next%next\ <= \$19080_next\;
      \$17386%next\ <= \$17386\;
      \$13982_v%next\ <= \$13982_v\;
      \$17459_loop665_arg%next\ <= \$17459_loop665_arg\;
      \$18719_w%next\ <= \$18719_w\;
      \$15445%next\ <= \$15445\;
      \$v7353%next\ <= \$v7353\;
      \$16752_fill6545929_result%next\ <= \$16752_fill6545929_result\;
      \$14997_modulo6685888_id%next\ <= \$14997_modulo6685888_id\;
      \$18050%next\ <= \$18050\;
      \$12883%next\ <= \$12883\;
      \$16823_compbranch6505931_arg%next\ <= \$16823_compbranch6505931_arg\;
      \$16233%next\ <= \$16233\;
      \$16271%next\ <= \$16271\;
      \$12682_make_block579_arg%next\ <= \$12682_make_block579_arg\;
      \$18655%next\ <= \$18655\;
      \$v7371%next\ <= \$v7371\;
      \$18987_hd%next\ <= \$18987_hd\;
      \$v6619%next\ <= \$v6619\;
      \$v6427%next\ <= \$v6427\;
      \$16748%next\ <= \$16748\;
      \$v6974%next\ <= \$v6974\;
      \$18474%next\ <= \$18474\;
      \$17886%next\ <= \$17886\;
      \$15756_compare6445897_arg%next\ <= \$15756_compare6445897_arg\;
      \$13151%next\ <= \$13151\;
      \$v6805%next\ <= \$v6805\;
      \$17569%next\ <= \$17569\;
      \$12698%next\ <= \$12698\;
      \$15389_modulo6685895_arg%next\ <= \$15389_modulo6685895_arg\;
      \$v6035%next\ <= \$v6035\;
      \$15553_r%next\ <= \$15553_r\;
      \$15237_modulo6685888_result%next\ <= \$15237_modulo6685888_result\;
      \$12944%next\ <= \$12944\;
      \$14613_modulo6685896_result%next\ <= \$14613_modulo6685896_result\;
      \$v7381%next\ <= \$v7381\;
      \$18846%next\ <= \$18846\;
      \$18917%next\ <= \$18917\;
      \$v6092%next\ <= \$v6092\;
      \$18916%next\ <= \$18916\;
      \$15261_modulo6685888_id%next\ <= \$15261_modulo6685888_id\;
      \$17679%next\ <= \$17679\;
      \$13154%next\ <= \$13154\;
      \$v6336%next\ <= \$v6336\;
      \$16527_f0%next\ <= \$16527_f0\;
      \$18352%next\ <= \$18352\;
      \$13964%next\ <= \$13964\;
      \$v7420%next\ <= \$v7420\;
      \$13632_next%next\ <= \$13632_next\;
      \$v6502%next\ <= \$v6502\;
      \$v6370%next\ <= \$v6370\;
      \$18739%next\ <= \$18739\;
      \$12714%next\ <= \$12714\;
      \$17484%next\ <= \$17484\;
      \$17597%next\ <= \$17597\;
      \$15756_compare6445897_result%next\ <= \$15756_compare6445897_result\;
      \$v7137%next\ <= \$v7137\;
      \$13532%next\ <= \$13532\;
      \$v6823%next\ <= \$v6823\;
      \$14781_modulo6685888_result%next\ <= \$14781_modulo6685888_result\;
      \$v6721%next\ <= \$v6721\;
      \$17734_copy_root_in_ram6635892_id%next\ <= \$17734_copy_root_in_ram6635892_id\;
      \$v7338%next\ <= \$v7338\;
      \$14749_modulo6685895_arg%next\ <= \$14749_modulo6685895_arg\;
      \$v7050%next\ <= \$v7050\;
      \$16299_v%next\ <= \$16299_v\;
      \$12689%next\ <= \$12689\;
      \$18807%next\ <= \$18807\;
      \$13920_loop666_arg%next\ <= \$13920_loop666_arg\;
      \$17455_loop666_id%next\ <= \$17455_loop666_id\;
      \$v6027%next\ <= \$v6027\;
      \$18650%next\ <= \$18650\;
      \$18837%next\ <= \$18837\;
      \$16951_compare6445898_arg%next\ <= \$16951_compare6445898_arg\;
      \$14861_modulo6685888_result%next\ <= \$14861_modulo6685888_result\;
      \$18805%next\ <= \$18805\;
      \$17543%next\ <= \$17543\;
      \$13997_v%next\ <= \$13997_v\;
      \$16574_compare6445898_id%next\ <= \$16574_compare6445898_id\;
      \$v6728%next\ <= \$v6728\;
      \$v6500%next\ <= \$v6500\;
      \$v5869%next\ <= \$v5869\;
      \$v6496%next\ <= \$v6496\;
      \$14978_v%next\ <= \$14978_v\;
      \$v7454%next\ <= \$v7454\;
      \$13237%next\ <= \$13237\;
      \$v6146%next\ <= \$v6146\;
      \$15330_r%next\ <= \$15330_r\;
      \$12839%next\ <= \$12839\;
      \$14061_v%next\ <= \$14061_v\;
      \$14701_modulo6685888_arg%next\ <= \$14701_modulo6685888_arg\;
      \$12697%next\ <= \$12697\;
      \$17773%next\ <= \$17773\;
      \$v7344%next\ <= \$v7344\;
      \$12888%next\ <= \$12888\;
      \$13155%next\ <= \$13155\;
      \$12937%next\ <= \$12937\;
      \$16115%next\ <= \$16115\;
      \$12805_aux664_result%next\ <= \$12805_aux664_result\;
      \$v6021%next\ <= \$v6021\;
      \$13697%next\ <= \$13697\;
      \$v6466%next\ <= \$v6466\;
      \$18355%next\ <= \$18355\;
      \rdy5940%next\ <= rdy5940;
      \$13102%next\ <= \$13102\;
      \$13235%next\ <= \$13235\;
      \$15044_binop_int6435906_id%next\ <= \$15044_binop_int6435906_id\;
      \$16729_v%next\ <= \$16729_v\;
      \$v6376%next\ <= \$v6376\;
      \$13233%next\ <= \$13233\;
      \$17670%next\ <= \$17670\;
      \$14555%next\ <= \$14555\;
      \$14564_binop_int6435900_result%next\ <= \$14564_binop_int6435900_result\;
      \$v6802%next\ <= \$v6802\;
      \$15058_v%next\ <= \$15058_v\;
      \$17464%next\ <= \$17464\;
      \$v6599%next\ <= \$v6599\;
      \$v6430%next\ <= \$v6430\;
      \$v6318%next\ <= \$v6318\;
      \$v7161%next\ <= \$v7161\;
      \$17669%next\ <= \$17669\;
      \$16963_compbranch6505935_id%next\ <= \$16963_compbranch6505935_id\;
      \$13967_v%next\ <= \$13967_v\;
      \$13696%next\ <= \$13696\;
      \$v6015%next\ <= \$v6015\;
      \$15476_modulo6685895_arg%next\ <= \$15476_modulo6685895_arg\;
      \$17470%next\ <= \$17470\;
      \$12520_loop666_id%next\ <= \$12520_loop666_id\;
      \$18815%next\ <= \$18815\;
      \$v6559%next\ <= \$v6559\;
      \$18565%next\ <= \$18565\;
      \$16551_compbranch6505926_id%next\ <= \$16551_compbranch6505926_id\;
      \$15397_modulo6685888_result%next\ <= \$15397_modulo6685888_result\;
      \$12877%next\ <= \$12877\;
      \$18698%next\ <= \$18698\;
      \$18480%next\ <= \$18480\;
      \$v7300%next\ <= \$v7300\;
      \$15389_modulo6685895_result%next\ <= \$15389_modulo6685895_result\;
      \$v7144%next\ <= \$v7144\;
      \$v6780%next\ <= \$v6780\;
      \$19256_hd%next\ <= \$19256_hd\;
      \$15823_res%next\ <= \$15823_res\;
      \$15124_binop_int6435907_id%next\ <= \$15124_binop_int6435907_id\;
      \$v6218%next\ <= \$v6218\;
      \$v7406%next\ <= \$v7406\;
      \$16963_compbranch6505935_arg%next\ <= \$16963_compbranch6505935_arg\;
      \$v7132%next\ <= \$v7132\;
      \$v7200%next\ <= \$v7200\;
      \$18633_loop665_id%next\ <= \$18633_loop665_id\;
      \$17888%next\ <= \$17888\;
      \$19145%next\ <= \$19145\;
      \$15625_binop_compare6455916_id%next\ <= \$15625_binop_compare6455916_id\;
      \$19337%next\ <= \$19337\;
      \$15893%next\ <= \$15893\;
      \$14364_v%next\ <= \$14364_v\;
      \$16893_compbranch6505933_result%next\ <= \$16893_compbranch6505933_result\;
      \$v6406%next\ <= \$v6406\;
      \$v6489%next\ <= \$v6489\;
      \$14837_modulo6685888_result%next\ <= \$14837_modulo6685888_result\;
      \$14677_modulo6685888_arg%next\ <= \$14677_modulo6685888_arg\;
      \$v6667%next\ <= \$v6667\;
      \$v7413%next\ <= \$v7413\;
      \$v6508%next\ <= \$v6508\;
      \$v6591%next\ <= \$v6591\;
      \$16284_v%next\ <= \$16284_v\;
      \$12808_aux664_result%next\ <= \$12808_aux664_result\;
      \$13816%next\ <= \$13816\;
      \$v6211%next\ <= \$v6211\;
      \$15874%next\ <= \$15874\;
      \$14829_modulo6685895_id%next\ <= \$14829_modulo6685895_id\;
      \$v7027%next\ <= \$v7027\;
      \$v6596%next\ <= \$v6596\;
      \$17746%next\ <= \$17746\;
      \$13950%next\ <= \$13950\;
      \$v5963%next\ <= \$v5963\;
      \$v5944%next\ <= \$v5944\;
      \$14597_modulo6685888_result%next\ <= \$14597_modulo6685888_result\;
      \$14582_res%next\ <= \$14582_res\;
      \$17891%next\ <= \$17891\;
      \$15397_modulo6685888_arg%next\ <= \$15397_modulo6685888_arg\;
      \$13927_branch_if648_result%next\ <= \$13927_branch_if648_result\;
      \$v7306%next\ <= \$v7306\;
      \$v7074%next\ <= \$v7074\;
      \$15021_modulo6685888_result%next\ <= \$15021_modulo6685888_result\;
      \$12707%next\ <= \$12707\;
      \$16881_compare6445898_result%next\ <= \$16881_compare6445898_result\;
      \$13679_w%next\ <= \$13679_w\;
      \$13663%next\ <= \$13663\;
      \$18447%next\ <= \$18447\;
      \$v6732%next\ <= \$v6732\;
      \$v6298%next\ <= \$v6298\;
      \$v6518%next\ <= \$v6518\;
      \$18278%next\ <= \$18278\;
      \$12544%next\ <= \$12544\;
      \$13218_w%next\ <= \$13218_w\;
      \$15932%next\ <= \$15932\;
      \$v7402%next\ <= \$v7402\;
      \$v7085%next\ <= \$v7085\;
      \$18731%next\ <= \$18731\;
      \$13519_w%next\ <= \$13519_w\;
      \$13606%next\ <= \$13606\;
      \$17776%next\ <= \$17776\;
      \$18644%next\ <= \$18644\;
      \$16327%next\ <= \$16327\;
      \$16169_v%next\ <= \$16169_v\;
      \$16551_compbranch6505926_arg%next\ <= \$16551_compbranch6505926_arg\;
      \$15229_modulo6685895_arg%next\ <= \$15229_modulo6685895_arg\;
      \$17457_aux664_result%next\ <= \$17457_aux664_result\;
      \$v6633%next\ <= \$v6633\;
      \$17665_hd%next\ <= \$17665_hd\;
      \$18159%next\ <= \$18159\;
      \$v6058%next\ <= \$v6058\;
      \$14122%next\ <= \$14122\;
      \$18563%next\ <= \$18563\;
      \$13310%next\ <= \$13310\;
      \$14012%next\ <= \$14012\;
      \$14677_modulo6685888_id%next\ <= \$14677_modulo6685888_id\;
      \$14181_sp%next\ <= \$14181_sp\;
      \$v6235%next\ <= \$v6235\;
      \$15961%next\ <= \$15961\;
      \$15476_modulo6685895_result%next\ <= \$15476_modulo6685895_result\;
      \$15237_modulo6685888_id%next\ <= \$15237_modulo6685888_id\;
      \$17505_forever6705894_arg%next\ <= \$17505_forever6705894_arg\;
      \$13388%next\ <= \$13388\;
      \$v6480%next\ <= \$v6480\;
      \$17001%next\ <= \$17001\;
      \$17963%next\ <= \$17963\;
      \$17803%next\ <= \$17803\;
      \$19142%next\ <= \$19142\;
      \$18679_forever6705881_id%next\ <= \$18679_forever6705881_id\;
      \$v6291%next\ <= \$v6291\;
      \$v6532%next\ <= \$v6532\;
      \$v7293%next\ <= \$v7293\;
      \$18919%next\ <= \$18919\;
      \$12685%next\ <= \$12685\;
      \$v6501%next\ <= \$v6501\;
      \$17238_sp%next\ <= \$17238_sp\;
      \$18186%next\ <= \$18186\;
      \$v7279%next\ <= \$v7279\;
      \$v6460%next\ <= \$v6460\;
      \$14431%next\ <= \$14431\;
      \$13667%next\ <= \$13667\;
      \$17455_loop666_arg%next\ <= \$17455_loop666_arg\;
      \$12851%next\ <= \$12851\;
      \$18188%next\ <= \$18188\;
      \$v6172%next\ <= \$v6172\;
      \$v7403%next\ <= \$v7403\;
      \$v7216%next\ <= \$v7216\;
      \$v7035%next\ <= \$v7035\;
      \$v6397%next\ <= \$v6397\;
      \$18709%next\ <= \$18709\;
      \$15720_compare6445897_id%next\ <= \$15720_compare6445897_id\;
      \$13823%next\ <= \$13823\;
      \$14177_hd%next\ <= \$14177_hd\;
      \result6503%next\ <= result6503;
      \$13395%next\ <= \$13395\;
      \$16353%next\ <= \$16353\;
      \$v6239%next\ <= \$v6239\;
      \$17559%next\ <= \$17559\;
      \$14351_v%next\ <= \$14351_v\;
      \$12808_aux664_id%next\ <= \$12808_aux664_id\;
      \$19269%next\ <= \$19269\;
      \$17412%next\ <= \$17412\;
      \$v7007%next\ <= \$v7007\;
      \$v6941%next\ <= \$v6941\;
      \$v6746%next\ <= \$v6746\;
      \$18925%next\ <= \$18925\;
      \$v6838%next\ <= \$v6838\;
      \$18733%next\ <= \$18733\;
      \$v5957%next\ <= \$v5957\;
      \$v6953%next\ <= \$v6953\;
      \$15783_v%next\ <= \$15783_v\;
      \$18279%next\ <= \$18279\;
      \$14207_loop_push6495899_result%next\ <= \$14207_loop_push6495899_result\;
      \$v6108%next\ <= \$v6108\;
      \$v7025%next\ <= \$v7025\;
      \$18120%next\ <= \$18120\;
      \$18566%next\ <= \$18566\;
      \$13016%next\ <= \$13016\;
      \$v6304%next\ <= \$v6304\;
      \$12692%next\ <= \$12692\;
      \$16037_v%next\ <= \$16037_v\;
      \$12935%next\ <= \$12935\;
      \$13625%next\ <= \$13625\;
      \$v7434%next\ <= \$v7434\;
      \$v6739%next\ <= \$v6739\;
      \$17509_forever6705890_arg%next\ <= \$17509_forever6705890_arg\;
      \$v6274%next\ <= \$v6274\;
      \$19001%next\ <= \$19001\;
      \$v7290%next\ <= \$v7290\;
      \$17498%next\ <= \$17498\;
      \$16945_b%next\ <= \$16945_b\;
      \$15298_v%next\ <= \$15298_v\;
      \$18346%next\ <= \$18346\;
      \$16589_compbranch6505927_id%next\ <= \$16589_compbranch6505927_id\;
      \$v6708%next\ <= \$v6708\;
      \$13157%next\ <= \$13157\;
      \$18909_hd%next\ <= \$18909_hd\;
      \$17674%next\ <= \$17674\;
      \$12712%next\ <= \$12712\;
      \$12945%next\ <= \$12945\;
      \$17354%next\ <= \$17354\;
      \$16574_compare6445898_result%next\ <= \$16574_compare6445898_result\;
      \$16365%next\ <= \$16365\;
      \$12715%next\ <= \$12715\;
      \$16510_forever6705925_id%next\ <= \$16510_forever6705925_id\;
      \$15218_v%next\ <= \$15218_v\;
      \$18699%next\ <= \$18699\;
      \$17591%next\ <= \$17591\;
      \$v6627%next\ <= \$v6627\;
      \$12915%next\ <= \$12915\;
      \$v6136%next\ <= \$v6136\;
      \$18045%next\ <= \$18045\;
      \$17460_aux664_id%next\ <= \$17460_aux664_id\;
      \$12807_loop665_id%next\ <= \$12807_loop665_id\;
      \$15069_modulo6685895_id%next\ <= \$15069_modulo6685895_id\;
      \$v6492%next\ <= \$v6492\;
      \$17487%next\ <= \$17487\;
      \$v6892%next\ <= \$v6892\;
      \$17387%next\ <= \$17387\;
      \$15386_r%next\ <= \$15386_r\;
      \$v6729%next\ <= \$v6729\;
      \$v6914%next\ <= \$v6914\;
      \$18915%next\ <= \$18915\;
      \$17105_w06555936_id%next\ <= \$17105_w06555936_id\;
      \$16589_compbranch6505927_arg%next\ <= \$16589_compbranch6505927_arg\;
      \$13890%next\ <= \$13890\;
      \$19144%next\ <= \$19144\;
      \$16677%next\ <= \$16677\;
      \$v7034%next\ <= \$v7034\;
      \$17678%next\ <= \$17678\;
      \$16875_b%next\ <= \$16875_b\;
      \$13927_branch_if648_arg%next\ <= \$13927_branch_if648_arg\;
      \$v6883%next\ <= \$v6883\;
      \$16438_v%next\ <= \$16438_v\;
      \$15612%next\ <= \$15612\;
      \$14773_modulo6685896_arg%next\ <= \$14773_modulo6685896_arg\;
      \$19140%next\ <= \$19140\;
      \$19071%next\ <= \$19071\;
      \$12848%next\ <= \$12848\;
      \$18831_hd%next\ <= \$18831_hd\;
      \$v6710%next\ <= \$v6710\;
      \$13468%next\ <= \$13468\;
      \$v6856%next\ <= \$v6856\;
      \$15317_modulo6685888_result%next\ <= \$15317_modulo6685888_result\;
      \$18570%next\ <= \$18570\;
      \$13623%next\ <= \$13623\;
      \$18128_next%next\ <= \$18128_next\;
      \$v7248%next\ <= \$v7248\;
      \$14644_binop_int6435901_result%next\ <= \$14644_binop_int6435901_result\;
      \$12679_loop666_id%next\ <= \$12679_loop666_id\;
      \$16399%next\ <= \$16399\;
      \$19263%next\ <= \$19263\;
      \$14749_modulo6685895_id%next\ <= \$14749_modulo6685895_id\;
      \$17794_w%next\ <= \$17794_w\;
      \result6468%next\ <= result6468;
      \$v7045%next\ <= \$v7045\;
      \$18816%next\ <= \$18816\;
      \$17885%next\ <= \$17885\;
      \$v7164%next\ <= \$v7164\;
      \$15101_modulo6685888_result%next\ <= \$15101_modulo6685888_result\;
      \$v7042%next\ <= \$v7042\;
      \$15500_modulo6685896_arg%next\ <= \$15500_modulo6685896_arg\;
      \$15333_modulo6685896_result%next\ <= \$15333_modulo6685896_result\;
      \$17761_copy_root_in_ram6635891_result%next\ <= \$17761_copy_root_in_ram6635891_result\;
      \$15720_compare6445897_arg%next\ <= \$15720_compare6445897_arg\;
      \$16713_v%next\ <= \$16713_v\;
      \$15697_binop_compare6455918_arg%next\ <= \$15697_binop_compare6455918_arg\;
      \$17250_v%next\ <= \$17250_v\;
      \$12887%next\ <= \$12887\;
      \$v6826%next\ <= \$v6826\;
      \$17394%next\ <= \$17394\;
      \$v6695%next\ <= \$v6695\;
      \$17333_sp%next\ <= \$17333_sp\;
      \$v7017%next\ <= \$v7017\;
      \$16158_forever6705923_arg%next\ <= \$16158_forever6705923_arg\;
      \$v6874%next\ <= \$v6874\;
      \$v6574%next\ <= \$v6574\;
      \$15853_v%next\ <= \$15853_v\;
      \$v7372%next\ <= \$v7372\;
      \$v6651%next\ <= \$v6651\;
      \$v7013%next\ <= \$v7013\;
      \$15181_modulo6685888_result%next\ <= \$15181_modulo6685888_result\;
      \$12691%next\ <= \$12691\;
      \$17962%next\ <= \$17962\;
      \$v6367%next\ <= \$v6367\;
      \$v6200%next\ <= \$v6200\;
      \$16612_compare6445898_result%next\ <= \$16612_compare6445898_result\;
      \$v6688%next\ <= \$v6688\;
      \$14330_v%next\ <= \$14330_v\;
      \$v7361%next\ <= \$v7361\;
      \$17319%next\ <= \$17319\;
      \$13941%next\ <= \$13941\;
      \$16078%next\ <= \$16078\;
      \$16165%next\ <= \$16165\;
      \$v7299%next\ <= \$v7299\;
      \$17012_sp%next\ <= \$17012_sp\;
      \$15261_modulo6685888_arg%next\ <= \$15261_modulo6685888_arg\;
      \$v6342%next\ <= \$v6342\;
      \$v5954%next\ <= \$v5954\;
      \$16606_b%next\ <= \$16606_b\;
      \$14986_r%next\ <= \$14986_r\;
      \$13301_hd%next\ <= \$13301_hd\;
      \$15847%next\ <= \$15847\;
      \$v7179%next\ <= \$v7179\;
      \$15021_modulo6685888_arg%next\ <= \$15021_modulo6685888_arg\;
      \$13127%next\ <= \$13127\;
      \$v7004%next\ <= \$v7004\;
      \$v7090%next\ <= \$v7090\;
      \$v6709%next\ <= \$v6709\;
      \$17321%next\ <= \$17321\;
      \$13530%next\ <= \$13530\;
      \$14222%next\ <= \$14222\;
      \$v6868%next\ <= \$v6868\;
      \$v6203%next\ <= \$v6203\;
      \$v5866%next\ <= \$v5866\;
      \$v5951%next\ <= \$v5951\;
      \$18450%next\ <= \$18450\;
      \$13296_w%next\ <= \$13296_w\;
      \$14724_binop_int6435902_id%next\ <= \$14724_binop_int6435902_id\;
      \$v7400%next\ <= \$v7400\;
      \$13013%next\ <= \$13013\;
      \$17349%next\ <= \$17349\;
      \$16192%next\ <= \$16192\;
      \$12834%next\ <= \$12834\;
      \$16441%next\ <= \$16441\;
      \$17167%next\ <= \$17167\;
      \$16042_v%next\ <= \$16042_v\;
      \$15697_binop_compare6455918_result%next\ <= \$15697_binop_compare6455918_result\;
      \$12679_loop666_result%next\ <= \$12679_loop666_result\;
      \$16234%next\ <= \$16234\;
      \$15625_binop_compare6455916_result%next\ <= \$15625_binop_compare6455916_result\;
      \$v7140%next\ <= \$v7140\;
      \$18163%next\ <= \$18163\;
      \$v6007%next\ <= \$v6007\;
      \$14933_modulo6685896_result%next\ <= \$14933_modulo6685896_result\;
      \$v7066%next\ <= \$v7066\;
      \$14818_v%next\ <= \$14818_v\;
      \$v6750%next\ <= \$v6750\;
      \$15976_v%next\ <= \$15976_v\;
      \$v6935%next\ <= \$v6935\;
      \$14338_v%next\ <= \$14338_v\;
      \$v6986%next\ <= \$v6986\;
      \$16805_b%next\ <= \$16805_b\;
      \$17961%next\ <= \$17961\;
      \$16439_v%next\ <= \$16439_v\;
      \$14933_modulo6685896_id%next\ <= \$14933_modulo6685896_id\;
      \$17681%next\ <= \$17681\;
      \$12910%next\ <= \$12910\;
      \$v6445%next\ <= \$v6445\;
      \$12741%next\ <= \$12741\;
      \$v7455%next\ <= \$v7455\;
      \$v6277%next\ <= \$v6277\;
      \$v6962%next\ <= \$v6962\;
      \$v7441%next\ <= \$v7441\;
      \$13962%next\ <= \$13962\;
      \$15010_r%next\ <= \$15010_r\;
      \$14829_modulo6685895_result%next\ <= \$14829_modulo6685895_result\;
      \$12521_loop665_arg%next\ <= \$12521_loop665_arg\;
      \$14161%next\ <= \$14161\;
      \$15805_binop_compare6455921_arg%next\ <= \$15805_binop_compare6455921_arg\;
      \$12843%next\ <= \$12843\;
      \$15413_modulo6685896_result%next\ <= \$15413_modulo6685896_result\;
      \$v7064%next\ <= \$v7064\;
      \$15484_modulo6685888_arg%next\ <= \$15484_modulo6685888_arg\;
      \$v7368%next\ <= \$v7368\;
      \$v6117%next\ <= \$v6117\;
      \$18634_aux664_result%next\ <= \$18634_aux664_result\;
      \$12943%next\ <= \$12943\;
      \$v6995%next\ <= \$v6995\;
      \$v6657%next\ <= \$v6657\;
      \$17600%next\ <= \$17600\;
      \$v6214%next\ <= \$v6214\;
      \$13957%next\ <= \$13957\;
      \$v7016%next\ <= \$v7016\;
      \$v6307%next\ <= \$v6307\;
      \$v6268%next\ <= \$v6268\;
      \$18982_w%next\ <= \$18982_w\;
      \$13103%next\ <= \$13103\;
      \$14517_v%next\ <= \$14517_v\;
      \$v7023%next\ <= \$v7023\;
      \$13692%next\ <= \$13692\;
      \$18479%next\ <= \$18479\;
      \$v7358%next\ <= \$v7358\;
      \$v6271%next\ <= \$v6271\;
      \$v6681%next\ <= \$v6681\;
      \$12806_loop666_result%next\ <= \$12806_loop666_result\;
      \$12680_loop665_result%next\ <= \$12680_loop665_result\;
      \$18734%next\ <= \$18734\;
      \$15484_modulo6685888_id%next\ <= \$15484_modulo6685888_id\;
      \$v6055%next\ <= \$v6055\;
      \$14746_r%next\ <= \$14746_r\;
      \$17327%next\ <= \$17327\;
      \$13153%next\ <= \$13153\;
      \$v6701%next\ <= \$v6701\;
      \$v7453%next\ <= \$v7453\;
      \$v6950%next\ <= \$v6950\;
      \$15733_binop_compare6455919_arg%next\ <= \$15733_binop_compare6455919_arg\;
      \$16436_v%next\ <= \$16436_v\;
      \$v7335%next\ <= \$v7335\;
      \$14837_modulo6685888_arg%next\ <= \$14837_modulo6685888_arg\;
      \$14558%next\ <= \$14558\;
      \$v6609%next\ <= \$v6609\;
      \$v6102%next\ <= \$v6102\;
      \$v6865%next\ <= \$v6865\;
      \$v7121%next\ <= \$v7121\;
      \$v6175%next\ <= \$v6175\;
      \$17520_copy_root_in_ram6635893_id%next\ <= \$17520_copy_root_in_ram6635893_id\;
      \$18818%next\ <= \$18818\;
      \$17018_w36575938_id%next\ <= \$17018_w36575938_id\;
      \$13946%next\ <= \$13946\;
      \$v7354%next\ <= \$v7354\;
      \$17315%next\ <= \$17315\;
      \$15204_binop_int6435908_id%next\ <= \$15204_binop_int6435908_id\;
      \$14658_v%next\ <= \$14658_v\;
      \$13307%next\ <= \$13307\;
      \$14042%next\ <= \$14042\;
      \$12939%next\ <= \$12939\;
      \$12891_copy_root_in_ram6635884_arg%next\ <= \$12891_copy_root_in_ram6635884_arg\;
      \$v7416%next\ <= \$v7416\;
      \$18166%next\ <= \$18166\;
      \$15556_modulo6685895_result%next\ <= \$15556_modulo6685895_result\;
      \$16035%next\ <= \$16035\;
      \$14853_modulo6685896_arg%next\ <= \$14853_modulo6685896_arg\;
      \$15124_binop_int6435907_arg%next\ <= \$15124_binop_int6435907_arg\;
      \$13928_w652_result%next\ <= \$13928_w652_result\;
      \$15317_modulo6685888_arg%next\ <= \$15317_modulo6685888_arg\;
      \$17377%next\ <= \$17377\;
      \$16126%next\ <= \$16126\;
      \$v7133%next\ <= \$v7133\;
      \$16127_v%next\ <= \$16127_v\;
      \$12878%next\ <= \$12878\;
      \$16031%next\ <= \$16031\;
      \$18836%next\ <= \$18836\;
      \$12857_forever6705883_arg%next\ <= \$12857_forever6705883_arg\;
      \$v7219%next\ <= \$v7219\;
      \$v6773%next\ <= \$v6773\;
      \$14114%next\ <= \$14114\;
      \$v7086%next\ <= \$v7086\;
      \$18999%next\ <= \$18999\;
      \$18637%next\ <= \$18637\;
      \$v6301%next\ <= \$v6301\;
      \$17734_copy_root_in_ram6635892_arg%next\ <= \$17734_copy_root_in_ram6635892_arg\;
      \$v5874%next\ <= \$v5874\;
      \$v7185%next\ <= \$v7185\;
      \$13693%next\ <= \$13693\;
      \$v6229%next\ <= \$v6229\;
      \$14285_v%next\ <= \$14285_v\;
      \$12734%next\ <= \$12734\;
      \$15341_modulo6685888_arg%next\ <= \$15341_modulo6685888_arg\;
      \$12904%next\ <= \$12904\;
      \$v7077%next\ <= \$v7077\;
      \$17513_forever6705889_id%next\ <= \$17513_forever6705889_id\;
      \$v6853%next\ <= \$v6853\;
      \$13466%next\ <= \$13466\;
      \$v7322%next\ <= \$v7322\;
      \$14804_binop_int6435903_arg%next\ <= \$14804_binop_int6435903_arg\;
      \$17463%next\ <= \$17463\;
      \$19115%next\ <= \$19115\;
      \$18904_w%next\ <= \$18904_w\;
      \$12818%next\ <= \$12818\;
      \$v6751%next\ <= \$v6751\;
      \$16292%next\ <= \$16292\;
      \$12844_next%next\ <= \$12844_next\;
      \$16395_v%next\ <= \$16395_v\;
      \$14964_binop_int6435905_id%next\ <= \$14964_binop_int6435905_id\;
      \$16767%next\ <= \$16767\;
      \$15093_modulo6685896_arg%next\ <= \$15093_modulo6685896_arg\;
      \$v6103%next\ <= \$v6103\;
      \$15648_compare6445897_id%next\ <= \$15648_compare6445897_id\;
      \$v6165%next\ <= \$v6165\;
      \$18104%next\ <= \$18104\;
      \$v7030%next\ <= \$v7030\;
      \$14613_modulo6685896_id%next\ <= \$14613_modulo6685896_id\;
      \$v6738%next\ <= \$v6738\;
      \$v6678%next\ <= \$v6678\;
      \$17491%next\ <= \$17491\;
      \$13078_copy_root_in_ram6635885_id%next\ <= \$13078_copy_root_in_ram6635885_id\;
      \$15981_v%next\ <= \$15981_v\;
      \$12560%next\ <= \$12560\;
      \$v7057%next\ <= \$v7057\;
      \$v6364%next\ <= \$v6364\;
      \$12702%next\ <= \$12702\;
      \$13312%next\ <= \$13312\;
      \$12520_loop666_arg%next\ <= \$12520_loop666_arg\;
      \$15792_compare6445897_result%next\ <= \$15792_compare6445897_result\;
      \$15341_modulo6685888_result%next\ <= \$15341_modulo6685888_result\;
      \$v7076%next\ <= \$v7076\;
      \$14669_modulo6685895_id%next\ <= \$14669_modulo6685895_id\;
      \$v5878%next\ <= \$v5878\;
      \$18711%next\ <= \$18711\;
      \$15828_compare6445897_id%next\ <= \$15828_compare6445897_id\;
      \$15237_modulo6685888_arg%next\ <= \$15237_modulo6685888_arg\;
      \$v6183%next\ <= \$v6183\;
      \$v5992%next\ <= \$v5992\;
      \$v6314%next\ <= \$v6314\;
      \$12522_wait662_result%next\ <= \$12522_wait662_result\;
      \$v6947%next\ <= \$v6947\;
      \$v6595%next\ <= \$v6595\;
      \$17455_loop666_result%next\ <= \$17455_loop666_result\;
      \$v7458%next\ <= \$v7458\;
      \$v6162%next\ <= \$v6162\;
      \$12838_next%next\ <= \$12838_next\;
      \$v6012%next\ <= \$v6012\;
      \$18472%next\ <= \$18472\;
      \$16036_sp%next\ <= \$16036_sp\;
      \$18185%next\ <= \$18185\;
      \$14424_v%next\ <= \$14424_v\;
      \$14254%next\ <= \$14254\;
      \$13389%next\ <= \$13389\;
      \$18677%next\ <= \$18677\;
      \$17348%next\ <= \$17348\;
      \$13393%next\ <= \$13393\;
      \$15769_binop_compare6455920_id%next\ <= \$15769_binop_compare6455920_id\;
      \$13387%next\ <= \$13387\;
      \$17590%next\ <= \$17590\;
      \$v7398%next\ <= \$v7398\;
      \$16823_compbranch6505931_id%next\ <= \$16823_compbranch6505931_id\;
      \$17495%next\ <= \$17495\;
      \$16379_v%next\ <= \$16379_v\;
      \$16881_compare6445898_arg%next\ <= \$16881_compare6445898_arg\;
      \$18679_forever6705881_arg%next\ <= \$18679_forever6705881_arg\;
      \$v6048%next\ <= \$v6048\;
      \$14677_modulo6685888_result%next\ <= \$14677_modulo6685888_result\;
      \$18288_next%next\ <= \$18288_next\;
      \$12538_cy%next\ <= \$12538_cy\;
      \$15378_v%next\ <= \$15378_v\;
      \$12941%next\ <= \$12941\;
      \$17783%next\ <= \$17783\;
      \$13794%next\ <= \$13794\;
      \$14693_modulo6685896_arg%next\ <= \$14693_modulo6685896_arg\;
      \$12914%next\ <= \$12914\;
      \$19262%next\ <= \$19262\;
      \$v6847%next\ <= \$v6847\;
      \$15382_res%next\ <= \$15382_res\;
      \$12521_loop665_result%next\ <= \$12521_loop665_result\;
      \$13238%next\ <= \$13238\;
      \$v6286%next\ <= \$v6286\;
      \$19070%next\ <= \$19070\;
      \$17254%next\ <= \$17254\;
      \$13694%next\ <= \$13694\;
      \$14941_modulo6685888_arg%next\ <= \$14941_modulo6685888_arg\;
      \$v7328%next\ <= \$v7328\;
      \$18356%next\ <= \$18356\;
      \$v7054%next\ <= \$v7054\;
      \$17761_copy_root_in_ram6635891_id%next\ <= \$17761_copy_root_in_ram6635891_id\;
      \$12695%next\ <= \$12695\;
      \$v6089%next\ <= \$v6089\;
      \$17774%next\ <= \$17774\;
      \$16231%next\ <= \$16231\;
      \$v7015%next\ <= \$v7015\;
      \$16202_ofs%next\ <= \$16202_ofs\;
      \$v7091%next\ <= \$v7091\;
      \$16217_hd%next\ <= \$16217_hd\;
      \$v6400%next\ <= \$v6400\;
      \$v6388%next\ <= \$v6388\;
      \$16024%next\ <= \$16024\;
      \$12913%next\ <= \$12913\;
      \$17048_w16565937_arg%next\ <= \$17048_w16565937_arg\;
      \$15476_modulo6685895_id%next\ <= \$15476_modulo6685895_id\;
      \$16823_compbranch6505931_result%next\ <= \$16823_compbranch6505931_result\;
      \$16928_compbranch6505934_result%next\ <= \$16928_compbranch6505934_result\;
      \$18475%next\ <= \$18475\;
      \$17890%next\ <= \$17890\;
      \$15580_modulo6685896_id%next\ <= \$15580_modulo6685896_id\;
      \$15828_compare6445897_result%next\ <= \$15828_compare6445897_result\;
      \$12936%next\ <= \$12936\;
      \$17165%next\ <= \$17165\;
      \$12660%next\ <= \$12660\;
      \$v7232%next\ <= \$v7232\;
      \$12736%next\ <= \$12736\;
      \$v6724%next\ <= \$v6724\;
      \$18724_hd%next\ <= \$18724_hd\;
      \$17775%next\ <= \$17775\;
      \$16630%next\ <= \$16630\;
      \$15341_modulo6685888_id%next\ <= \$15341_modulo6685888_id\;
      \$18187%next\ <= \$18187\;
      \$v6998%next\ <= \$v6998\;
      \$17580_w%next\ <= \$17580_w\;
      \$17785%next\ <= \$17785\;
      \$12716%next\ <= \$12716\;
      \$15253_modulo6685896_id%next\ <= \$15253_modulo6685896_id\;
      \$14135%next\ <= \$14135\;
      \$15828_compare6445897_arg%next\ <= \$15828_compare6445897_arg\;
      \$13129%next\ <= \$13129\;
      \$18194%next\ <= \$18194\;
      \$18193%next\ <= \$18193\;
      \$16916_compare6445898_arg%next\ <= \$16916_compare6445898_arg\;
      \$17812%next\ <= \$17812\;
      \$12806_loop666_id%next\ <= \$12806_loop666_id\;
      \$15204_binop_int6435908_result%next\ <= \$15204_binop_int6435908_result\;
      \$v7210%next\ <= \$v7210\;
      \$17457_aux664_arg%next\ <= \$17457_aux664_arg\;
      \$14453_next_acc%next\ <= \$14453_next_acc\;
      \$18571%next\ <= \$18571\;
      \$15309_modulo6685895_result%next\ <= \$15309_modulo6685895_result\;
      \$17879_hd%next\ <= \$17879_hd\;
      \$13138_w%next\ <= \$13138_w\;
      \$v6624%next\ <= \$v6624\;
      \$v6992%next\ <= \$v6992\;
      \$14644_binop_int6435901_arg%next\ <= \$14644_binop_int6435901_arg\;
      \$v6515%next\ <= \$v6515\;
      \$13507%next\ <= \$13507\;
      \$19235%next\ <= \$19235\;
      \$17593%next\ <= \$17593\;
      \$17460_aux664_result%next\ <= \$17460_aux664_result\;
      \$v7283%next\ <= \$v7283\;
      \$16986_compare6445898_result%next\ <= \$16986_compare6445898_result\;
      \$14930_r%next\ <= \$14930_r\;
      \$v6898%next\ <= \$v6898\;
      \$v6003%next\ <= \$v6003\;
      \$17466%next\ <= \$17466\;
      \$v6579%next\ <= \$v6579\;
      \$v6121%next\ <= \$v6121\;
      \$14621_modulo6685888_result%next\ <= \$14621_modulo6685888_result\;
      \$13689%next\ <= \$13689\;
      \$14804_binop_int6435903_result%next\ <= \$14804_binop_int6435903_result\;
      \$12782%next\ <= \$12782\;
      \$18995%next\ <= \$18995\;
      \$v6110%next\ <= \$v6110\;
      \$v6179%next\ <= \$v6179\;
      \$18043%next\ <= \$18043\;
      \$19251_w%next\ <= \$19251_w\;
      \$14381%next\ <= \$14381\;
      \$v6066%next\ <= \$v6066\;
      \$12546_dur%next\ <= \$12546_dur\;
      \$v6911%next\ <= \$v6911\;
      \$v6207%next\ <= \$v6207\;
      \$15253_modulo6685896_result%next\ <= \$15253_modulo6685896_result\;
      \$17889%next\ <= \$17889\;
      \$14311%next\ <= \$14311\;
      \$v6971%next\ <= \$v6971\;
      \$v5999%next\ <= \$v5999\;
      \$12906%next\ <= \$12906\;
      \$v7206%next\ <= \$v7206\;
      \$14917_modulo6685888_id%next\ <= \$14917_modulo6685888_id\;
      \$18661%next\ <= \$18661\;
      \$17957_hd%next\ <= \$17957_hd\;
      \$12924_w%next\ <= \$12924_w\;
      \$v6546%next\ <= \$v6546\;
      \$18280%next\ <= \$18280\;
      \$13148%next\ <= \$13148\;
      \$v6232%next\ <= \$v6232\;
      \$18633_loop665_arg%next\ <= \$18633_loop665_arg\;
      \$14757_modulo6685888_result%next\ <= \$14757_modulo6685888_result\;
      \$13922_wait662_result%next\ <= \$13922_wait662_result\;
      \$v7364%next\ <= \$v7364\;
      \$15580_modulo6685896_result%next\ <= \$15580_modulo6685896_result\;
      \$15421_modulo6685888_id%next\ <= \$15421_modulo6685888_id\;
      \$14610_r%next\ <= \$14610_r\;
      \$16916_compare6445898_id%next\ <= \$16916_compare6445898_id\;
      \$12886%next\ <= \$12886\;
      \$16195_forever6705924_id%next\ <= \$16195_forever6705924_id\;
      \$v6670%next\ <= \$v6670\;
      \$13817%next\ <= \$13817\;
      \$v6817%next\ <= \$v6817\;
      \$14221%next\ <= \$14221\;
      \$v6062%next\ <= \$v6062\;
      \$17389%next\ <= \$17389\;
      \$v6563%next\ <= \$v6563\;
      \$v6080%next\ <= \$v6080\;
      \$v6799%next\ <= \$v6799\;
      \$v7092%next\ <= \$v7092\;
      \$14296%next\ <= \$14296\;
      \$17815%next\ <= \$17815\;
      \$v6463%next\ <= \$v6463\;
      \$13100%next\ <= \$13100\;
      \$v6097%next\ <= \$v6097\;
      \$v7203%next\ <= \$v7203\;
      \$13808_hd%next\ <= \$13808_hd\;
      \$13822%next\ <= \$13822\;
      \$16121_v%next\ <= \$16121_v\;
      \$v6403%next\ <= \$v6403\;
      \$17000_sp%next\ <= \$17000_sp\;
      \$12735%next\ <= \$12735\;
      \$v6424%next\ <= \$v6424\;
      \$15261_modulo6685888_result%next\ <= \$15261_modulo6685888_result\;
      \$17500%next\ <= \$17500\;
      \$17805%next\ <= \$17805\;
      \$v6421%next\ <= \$v6421\;
      \$13510%next\ <= \$13510\;
      \$13940%next\ <= \$13940\;
      \$v7433%next\ <= \$v7433\;
      \$15309_modulo6685895_arg%next\ <= \$15309_modulo6685895_arg\;
      \$18657%next\ <= \$18657\;
      \$16574_compare6445898_arg%next\ <= \$16574_compare6445898_arg\;
      \$13317%next\ <= \$13317\;
      \$v6287%next\ <= \$v6287\;
      \$12903%next\ <= \$12903\;
      \$16382%next\ <= \$16382\;
      \$15897%next\ <= \$15897\;
      \$14941_modulo6685888_result%next\ <= \$14941_modulo6685888_result\;
      \$14909_modulo6685895_result%next\ <= \$14909_modulo6685895_result\;
      \$v7135%next\ <= \$v7135\;
      \$18806%next\ <= \$18806\;
      \$17458_loop666_arg%next\ <= \$17458_loop666_arg\;
      \$12938%next\ <= \$12938\;
      \$15531_binop_int6435913_id%next\ <= \$15531_binop_int6435913_id\;
      \$15284_binop_int6435909_id%next\ <= \$15284_binop_int6435909_id\;
      \$13700%next\ <= \$13700\;
      \$18843%next\ <= \$18843\;
      \$15364_binop_int6435910_id%next\ <= \$15364_binop_int6435910_id\;
      \$12523_make_block579_arg%next\ <= \$12523_make_block579_arg\;
      \$v7245%next\ <= \$v7245\;
      \$16317%next\ <= \$16317\;
      \$18348%next\ <= \$18348\;
      \$13101%next\ <= \$13101\;
      \$v6069%next\ <= \$v6069\;
      \$16063_w6515922_result%next\ <= \$16063_w6515922_result\;
      \$v6096%next\ <= \$v6096\;
      \$12864_copy_root_in_ram6635886_arg%next\ <= \$12864_copy_root_in_ram6635886_arg\;
      \$14669_modulo6685895_arg%next\ <= \$14669_modulo6685895_arg\;
      \$17561%next\ <= \$17561\;
      \$19118%next\ <= \$19118\;
      \$14837_modulo6685888_id%next\ <= \$14837_modulo6685888_id\;
      \$12694%next\ <= \$12694\;
      \$15284_binop_int6435909_arg%next\ <= \$15284_binop_int6435909_arg\;
      \$12701%next\ <= \$12701\;
      \$v7450%next\ <= \$v7450\;
      \$16158_forever6705923_id%next\ <= \$16158_forever6705923_id\;
      \$15101_modulo6685888_id%next\ <= \$15101_modulo6685888_id\;
      \$v7145%next\ <= \$v7145\;
      \$v6654%next\ <= \$v6654\;
      \$v6042%next\ <= \$v6042\;
      \$13234%next\ <= \$13234\;
      \$v6717%next\ <= \$v6717\;
      \$15580_modulo6685896_arg%next\ <= \$15580_modulo6685896_arg\;
      \$15500_modulo6685896_result%next\ <= \$15500_modulo6685896_result\;
      \$15447_forever6705911_arg%next\ <= \$15447_forever6705911_arg\;
      \$18189%next\ <= \$18189\;
      \rdy6469%next\ <= rdy6469;
      \$17964%next\ <= \$17964\;
      \$18319%next\ <= \$18319\;
      \$v6920%next\ <= \$v6920\;
      \$v6989%next\ <= \$v6989\;
      \$14315_v%next\ <= \$14315_v\;
      \$18124%next\ <= \$18124\;
      \$16321%next\ <= \$16321\;
      \$v5986%next\ <= \$v5986\;
      \$13384%next\ <= \$13384\;
      \$13379_hd%next\ <= \$13379_hd\;
      \$15421_modulo6685888_arg%next\ <= \$15421_modulo6685888_arg\;
      \$v7365%next\ <= \$v7365\;
      \$13922_wait662_id%next\ <= \$13922_wait662_id\;
      \$12549%next\ <= \$12549\;
      \$v6832%next\ <= \$v6832\;
      \$v6765%next\ <= \$v6765\;
      \$v6104%next\ <= \$v6104\;
      \$18730%next\ <= \$18730\;
      \$18184%next\ <= \$18184\;
      \$17892%next\ <= \$17892\;
      \$v6543%next\ <= \$v6543\;
      \$v6585%next\ <= \$v6585\;
      \$17671%next\ <= \$17671\;
      \$v6106%next\ <= \$v6106\;
      \$12704%next\ <= \$12704\;
      \$v7399%next\ <= \$v7399\;
      \$v7110%next\ <= \$v7110\;
      \$18118%next\ <= \$18118\;
      \$13540%next\ <= \$13540\;
      \$v6862%next\ <= \$v6862\;
      \$15508_modulo6685888_result%next\ <= \$15508_modulo6685888_result\;
      \$v7100%next\ <= \$v7100\;
      \$17513_forever6705889_arg%next\ <= \$17513_forever6705889_arg\;
      \$v6835%next\ <= \$v6835\;
      \$16203%next\ <= \$16203\;
      \$15229_modulo6685895_result%next\ <= \$15229_modulo6685895_result\;
      \$15910%next\ <= \$15910\;
      \$17456_loop665_result%next\ <= \$17456_loop665_result\;
      \$v5995%next\ <= \$v5995\;
      \$13765%next\ <= \$13765\;
      \$12807_loop665_result%next\ <= \$12807_loop665_result\;
      \$v6373%next\ <= \$v6373\;
      \$v6171%next\ <= \$v6171\;
      \$18473%next\ <= \$18473\;
      \$v6758%next\ <= \$v6758\;
      \$v7332%next\ <= \$v7332\;
      \$v6646%next\ <= \$v6646\;
      \$v6692%next\ <= \$v6692\;
      \$v7188%next\ <= \$v7188\;
      \$16063_w6515922_id%next\ <= \$16063_w6515922_id\;
      \$v6562%next\ <= \$v6562\;
      \$v6743%next\ <= \$v6743\;
      \$v7426%next\ <= \$v7426\;
      \$13463%next\ <= \$13463\;
      \$18686_copy_root_in_ram6635880_id%next\ <= \$18686_copy_root_in_ram6635880_id\;
      \$v7378%next\ <= \$v7378\;
      \$v6742%next\ <= \$v6742\;
      \$14989_modulo6685895_result%next\ <= \$14989_modulo6685895_result\;
      \$v7375%next\ <= \$v7375\;
      \$15204_binop_int6435908_arg%next\ <= \$15204_binop_int6435908_arg\;
      \$18845%next\ <= \$18845\;
      \$14008%next\ <= \$14008\;
      \$v6328%next\ <= \$v6328\;
      \$v7355%next\ <= \$v7355\;
      \$v7044%next\ <= \$v7044\;
      \$v6319%next\ <= \$v6319\;
      \$15364_binop_int6435910_arg%next\ <= \$15364_binop_int6435910_arg\;
      \$v6965%next\ <= \$v6965\;
      \$12879%next\ <= \$12879\;
      \$15284_binop_int6435909_result%next\ <= \$15284_binop_int6435909_result\;
      \$12804_loop665_result%next\ <= \$12804_loop665_result\;
      \$18546%next\ <= \$18546\;
      \$v7020%next\ <= \$v7020\;
      \$15564_modulo6685888_result%next\ <= \$15564_modulo6685888_result\;
      \$v7081%next\ <= \$v7081\;
      \$v5872%next\ <= \$v5872\;
      \$v7393%next\ <= \$v7393\;
      \$14152%next\ <= \$14152\;
      \$v6766%next\ <= \$v6766\;
      \$18841%next\ <= \$18841\;
      \$15661_binop_compare6455917_result%next\ <= \$15661_binop_compare6455917_result\;
      \$13316%next\ <= \$13316\;
      \$13009_hd%next\ <= \$13009_hd\;
      \$14909_modulo6685895_arg%next\ <= \$14909_modulo6685895_arg\;
      \$12682_make_block579_result%next\ <= \$12682_make_block579_result\;
      \$18738%next\ <= \$18738\;
      \$16509%next\ <= \$16509\;
      \$12688%next\ <= \$12688\;
      \$15577_r%next\ <= \$15577_r\;
      \$v6093%next\ <= \$v6093\;
      \$v6109%next\ <= \$v6109\;
      \$15564_modulo6685888_arg%next\ <= \$15564_modulo6685888_arg\;
      \$16928_compbranch6505934_id%next\ <= \$16928_compbranch6505934_id\;
      \$14884_binop_int6435904_arg%next\ <= \$14884_binop_int6435904_arg\;
      \$v6553%next\ <= \$v6553\;
      \$14092%next\ <= \$14092\;
      \$v6535%next\ <= \$v6535\;
      \$18732%next\ <= \$18732\;
      \$17066%next\ <= \$17066\;
      \$15389_modulo6685895_id%next\ <= \$15389_modulo6685895_id\;
      \$v6660%next\ <= \$v6660\;
      \$17337%next\ <= \$17337\;
      \$18826_w%next\ <= \$18826_w\;
      \$v6036%next\ <= \$v6036\;
      \$17374_v%next\ <= \$17374_v\;
      \$17502%next\ <= \$17502\;
      \$12942%next\ <= \$12942\;
      \$14773_modulo6685896_id%next\ <= \$14773_modulo6685896_id\;
      \$14757_modulo6685888_id%next\ <= \$14757_modulo6685888_id\;
      \$18041%next\ <= \$18041\;
      \$v6547%next\ <= \$v6547\;
      \$v6184%next\ <= \$v6184\;
      \$12864_copy_root_in_ram6635886_id%next\ <= \$12864_copy_root_in_ram6635886_id\;
      \$18470%next\ <= \$18470\;
      \$12835%next\ <= \$12835\;
      \$15909%next\ <= \$15909\;
      \$v6902%next\ <= \$v6902\;
      \$17009_sp%next\ <= \$17009_sp\;
      \$18476%next\ <= \$18476\;
      \$16626%next\ <= \$16626\;
      \$17804%next\ <= \$17804\;
      \$18443%next\ <= \$18443\;
      \$14701_modulo6685888_result%next\ <= \$14701_modulo6685888_result\;
      \$v7167%next\ <= \$v7167\;
      \$14902_res%next\ <= \$14902_res\;
      \$12717%next\ <= \$12717\;
      \$v6908%next\ <= \$v6908\;
      \$13917%next\ <= \$13917\;
      \$16749_sp%next\ <= \$16749_sp\;
      \$v6155%next\ <= \$v6155\;
      \$17243%next\ <= \$17243\;
      \$v6442%next\ <= \$v6442\;
      \$13923_make_block579_result%next\ <= \$13923_make_block579_result\;
      \$v7445%next\ <= \$v7445\;
      \$v6354%next\ <= \$v6354\;
      \$14508_v%next\ <= \$14508_v\;
      \$15157_modulo6685888_arg%next\ <= \$15157_modulo6685888_arg\;
      \$19267%next\ <= \$19267\;
      \$16846_compare6445898_id%next\ <= \$16846_compare6445898_id\;
      \$15170_r%next\ <= \$15170_r\;
      \$v6616%next\ <= \$v6616\;
      \$13926_make_block_n646_id%next\ <= \$13926_make_block_n646_id\;
      \$18478%next\ <= \$18478\;
      \$16440%next\ <= \$16440\;
      \$15451_binop_int6435912_arg%next\ <= \$15451_binop_int6435912_arg\;
      \$15980_v%next\ <= \$15980_v\;
      \$v6623%next\ <= \$v6623\;
      \$14909_modulo6685895_id%next\ <= \$14909_modulo6685895_id\;
      \$12830%next\ <= \$12830\;
      \$13149%next\ <= \$13149\;
      \$17164%next\ <= \$17164\;
      \$14463_v%next\ <= \$14463_v\;
      \$13019%next\ <= \$13019\;
      \$15613%next\ <= \$15613\;
      \$17535%next\ <= \$17535\;
      \$13818%next\ <= \$13818\;
      \$v6521%next\ <= \$v6521\;
      \$16763_v%next\ <= \$16763_v\;
      \$18669%next\ <= \$18669\;
      \$18660%next\ <= \$18660\;
      \$v6137%next\ <= \$v6137\;
      \$v6790%next\ <= \$v6790\;
      \$v7117%next\ <= \$v7117\;
      \$v6223%next\ <= \$v6223\;
      \$13105_copy_root_in_ram6635884_arg%next\ <= \$13105_copy_root_in_ram6635884_arg\;
      \$v7387%next\ <= \$v7387\;
      \$17547_copy_root_in_ram6635891_id%next\ <= \$17547_copy_root_in_ram6635891_id\;
      \$15157_modulo6685888_id%next\ <= \$15157_modulo6685888_id\;
      \$18632_loop666_arg%next\ <= \$18632_loop666_arg\;
      \$17173%next\ <= \$17173\;
      \$15447_forever6705911_id%next\ <= \$15447_forever6705911_id\;
      \$15861_v%next\ <= \$15861_v\;
      \$13223_hd%next\ <= \$13223_hd\;
      \$13524_hd%next\ <= \$13524_hd\;
      \$16336%next\ <= \$16336\;
      \$v6899%next\ <= \$v6899\;
      \$v7156%next\ <= \$v7156\;
      \$15302_res%next\ <= \$15302_res\;
      \$19268%next\ <= \$19268\;
      \$18572%next\ <= \$18572\;
      \$v7459%next\ <= \$v7459\;
      \$v7229%next\ <= \$v7229\;
      \$17883%next\ <= \$17883\;
      \$18048%next\ <= \$18048\;
      \$13385%next\ <= \$13385\;
      \$17239_v%next\ <= \$17239_v\;
      \$14773_modulo6685896_result%next\ <= \$14773_modulo6685896_result\;
      \$17592%next\ <= \$17592\;
      \$13926_make_block_n646_result%next\ <= \$13926_make_block_n646_result\;
      \$17749%next\ <= \$17749\;
      \$18668%next\ <= \$18668\;
      \$v7093%next\ <= \$v7093\;
      \$v6176%next\ <= \$v6176\;
      \$12710%next\ <= \$12710\;
      \$18913%next\ <= \$18913\;
      \$v7107%next\ <= \$v7107\;
      \$v6075%next\ <= \$v6075\;
      \$v6031%next\ <= \$v6031\;
      \$14861_modulo6685888_arg%next\ <= \$14861_modulo6685888_arg\;
      \$v6352%next\ <= \$v6352\;
      \$13924_apply638_result%next\ <= \$13924_apply638_result\;
      \$15883%next\ <= \$15883\;
      \$v6684%next\ <= \$v6684\;
      \$13309%next\ <= \$13309\;
      \$12829%next\ <= \$12829\;
      \$14273%next\ <= \$14273\;
      \rdy6504%next\ <= rdy6504;
      \$v6938%next\ <= \$v6938\;
      \$17371_v%next\ <= \$17371_v\;
      \$v6880%next\ <= \$v6880\;
      \$v7011%next\ <= \$v7011\;
      \$17232%next\ <= \$17232\;
      \$12864_copy_root_in_ram6635886_result%next\ <= \$12864_copy_root_in_ram6635886_result\;
      \$v6829%next\ <= \$v6829\;
      \$v7056%next\ <= \$v7056\;
      \$14139%next\ <= \$14139\;
      \$v6379%next\ <= \$v6379\;
      \$17332_sp%next\ <= \$17332_sp\;
      \$17048_w16565937_result%next\ <= \$17048_w16565937_result\;
      \$19266%next\ <= \$19266\;
      \$15588_modulo6685888_result%next\ <= \$15588_modulo6685888_result\;
      \$v7260%next\ <= \$v7260\;
      \$14621_modulo6685888_arg%next\ <= \$14621_modulo6685888_arg\;
      \$13924_apply638_arg%next\ <= \$13924_apply638_arg\;
      \$v6643%next\ <= \$v6643\;
      \$v6152%next\ <= \$v6152\;
      \$18994%next\ <= \$18994\;
      \$15250_r%next\ <= \$15250_r\;
      \$15044_binop_int6435906_result%next\ <= \$15044_binop_int6435906_result\;
      \$16650_sp%next\ <= \$16650_sp\;
      \$v7350%next\ <= \$v7350\;
      \$18633_loop665_result%next\ <= \$18633_loop665_result\;
      \$12553%next\ <= \$12553\;
      \$18044%next\ <= \$18044\;
      \$12720%next\ <= \$12720\;
      \$17594%next\ <= \$17594\;
      \$v6190%next\ <= \$v6190\;
      \$v5964%next\ <= \$v5964\;
      \$13926_make_block_n646_arg%next\ <= \$13926_make_block_n646_arg\;
      \$15077_modulo6685888_id%next\ <= \$15077_modulo6685888_id\;
      \$v7021%next\ <= \$v7021\;
      \$17018_w36575938_result%next\ <= \$17018_w36575938_result\;
      \$v6180%next\ <= \$v6180\;
      \$v6889%next\ <= \$v6889\;
      \$15715_res%next\ <= \$15715_res\;
      \$16349_v%next\ <= \$16349_v\;
      \$14964_binop_int6435905_arg%next\ <= \$14964_binop_int6435905_arg\;
      \$18998%next\ <= \$18998\;
      \$13158%next\ <= \$13158\;
      \$v6283%next\ <= \$v6283\;
      \$17393%next\ <= \$17393\;
      \$v5948%next\ <= \$v5948\;
      \$13092%next\ <= \$13092\;
      \$v6714%next\ <= \$v6714\;
      \$v6325%next\ <= \$v6325\;
      \$14997_modulo6685888_result%next\ <= \$14997_modulo6685888_result\;
      \$v6550%next\ <= \$v6550\;
      \$v6236%next\ <= \$v6236\;
      \$12934%next\ <= \$12934\;
      \$v6588%next\ <= \$v6588\;
      \$v6256%next\ <= \$v6256\;
      \$17458_loop666_id%next\ <= \$17458_loop666_id\;
      \$17032%next\ <= \$17032\;
      \$12706%next\ <= \$12706\;
      \$16673_v%next\ <= \$16673_v\;
      \$13688%next\ <= \$13688\;
      \$v7427%next\ <= \$v7427\;
      \$17458_loop666_result%next\ <= \$17458_loop666_result\;
      \$12681_wait662_arg%next\ <= \$12681_wait662_arg\;
      \$18673%next\ <= \$18673\;
      \$17324%next\ <= \$17324\;
      \$14070_v%next\ <= \$14070_v\;
      \$12737%next\ <= \$12737\;
      \$19214%next\ <= \$19214\;
      \$15787_res%next\ <= \$15787_res\;
      \$14589_modulo6685895_arg%next\ <= \$14589_modulo6685895_arg\;
      \$v5967%next\ <= \$v5967\;
      \$17968%next\ <= \$17968\;
      \$14738_v%next\ <= \$14738_v\;
      \$v5998%next\ <= \$v5998\;
      \$18639%next\ <= \$18639\;
      \$13766%next\ <= \$13766\;
      \$15413_modulo6685896_arg%next\ <= \$15413_modulo6685896_arg\;
      \$15860%next\ <= \$15860\;
      \$v7010%next\ <= \$v7010\;
      \$18564%next\ <= \$18564\;
      \$v7449%next\ <= \$v7449\;
      \$v7046%next\ <= \$v7046\;
      \$17532%next\ <= \$17532\;
      \$v6243%next\ <= \$v6243\;
      \$19213%next\ <= \$19213\;
      \$13529%next\ <= \$13529\;
      \$v6493%next\ <= \$v6493\;
      \$15421_modulo6685888_result%next\ <= \$15421_modulo6685888_result\;
      \$18191%next\ <= \$18191\;
      \$14564_binop_int6435900_id%next\ <= \$14564_binop_int6435900_id\;
      \$12679_loop666_arg%next\ <= \$12679_loop666_arg\;
      \$14406_v%next\ <= \$14406_v\;
      \$15619%next\ <= \$15619\;
      \$v6917%next\ <= \$v6917\;
      \$16507%next\ <= \$16507\;
      \$v7116%next\ <= \$v7116\;
      \$v7273%next\ <= \$v7273\;
      \$14165%next\ <= \$14165\;
      \$13920_loop666_id%next\ <= \$13920_loop666_id\;
      \$15618%next\ <= \$15618\;
      \$16403%next\ <= \$16403\;
      \$17476%next\ <= \$17476\;
      \$13626%next\ <= \$13626\;
      \$17967%next\ <= \$17967\;
      \$12709%next\ <= \$12709\;
      \$v7213%next\ <= \$v7213\;
      \$14861_modulo6685888_id%next\ <= \$14861_modulo6685888_id\;
      \$v6844%next\ <= \$v6844\;
      \$12804_loop665_arg%next\ <= \$12804_loop665_arg\;
      \$14281%next\ <= \$14281\;
      \$16272%next\ <= \$16272\;
      \$17572%next\ <= \$17572\;
      \$12705%next\ <= \$12705\;
      \$12696%next\ <= \$12696\;
      \$13117%next\ <= \$13117\;
      \$13605%next\ <= \$13605\;
      \$16288%next\ <= \$16288\;
      \$12853_forever6705887_id%next\ <= \$12853_forever6705887_id\;
      \$17734_copy_root_in_ram6635892_result%next\ <= \$17734_copy_root_in_ram6635892_result\;
      \$17759%next\ <= \$17759\;
      \$v6247%next\ <= \$v6247\;
      \$16986_compare6445898_id%next\ <= \$16986_compare6445898_id\;
      \$17314%next\ <= \$17314\;
      \$v7197%next\ <= \$v7197\;
      \$12680_loop665_arg%next\ <= \$12680_loop665_arg\;
      \$18119%next\ <= \$18119\;
      \$v6072%next\ <= \$v6072\;
      \$12760%next\ <= \$12760\;
      \$12548_dis%next\ <= \$12548_dis\;
      \$15077_modulo6685888_arg%next\ <= \$15077_modulo6685888_arg\;
      \$14853_modulo6685896_result%next\ <= \$14853_modulo6685896_result\;
      \$18737%next\ <= \$18737\;
      \$18918%next\ <= \$18918\;
      \$17237_sp%next\ <= \$17237_sp\;
      \$15173_modulo6685896_arg%next\ <= \$15173_modulo6685896_arg\;
      \$17595%next\ <= \$17595\;
      \$17008%next\ <= \$17008\;
      \$17761_copy_root_in_ram6635891_arg%next\ <= \$17761_copy_root_in_ram6635891_arg\;
      \$v7101%next\ <= \$v7101\;
      \$12847%next\ <= \$12847\;
      \$v6859%next\ <= \$v6859\;
      \$12889%next\ <= \$12889\;
      \$18051%next\ <= \$18051\;
      \$v6219%next\ <= \$v6219\;
      \$14826_r%next\ <= \$14826_r\;
      \$14033%next\ <= \$14033\;
      \$v6606%next\ <= \$v6606\;
      \$18326%next\ <= \$18326\;
      \$18921%next\ <= \$18921\;
      \$13691%next\ <= \$13691\;
      \$v7083%next\ <= \$v7083\;
      \$v6956%next\ <= \$v6956\;
      \$15679_res%next\ <= \$15679_res\;
      \$v6666%next\ <= \$v6666\;
      \$19239%next\ <= \$19239\;
      \$14024%next\ <= \$14024\;
      \$v7442%next\ <= \$v7442\;
      \$16811_compare6445898_result%next\ <= \$16811_compare6445898_result\;
      \$14781_modulo6685888_arg%next\ <= \$14781_modulo6685888_arg\;
      \$v6335%next\ <= \$v6335\;
      \$19260%next\ <= \$19260\;
      \$17347%next\ <= \$17347\;
      \$15333_modulo6685896_id%next\ <= \$15333_modulo6685896_id\;
      \$18196%next\ <= \$18196\;
      \$v6752%next\ <= \$v6752\;
      \$16300%next\ <= \$16300\;
      \$17673%next\ <= \$17673\;
      \$13227%next\ <= \$13227\;
      \$16612_compare6445898_arg%next\ <= \$16612_compare6445898_arg\;
      \$13925_offsetclosure_n639_result%next\ <= \$13925_offsetclosure_n639_result\;
      \$v6409%next\ <= \$v6409\;
      \$17814%next\ <= \$17814\;
      \$17585_hd%next\ <= \$17585_hd\;
      \$17509_forever6705890_id%next\ <= \$17509_forever6705890_id\;
      \$17566%next\ <= \$17566\;
      \$12814%next\ <= \$12814\;
      \$19242%next\ <= \$19242\;
      \$17497%next\ <= \$17497\;
      \$13695%next\ <= \$13695\;
      \$v6394%next\ <= \$v6394\;
      \$v7397%next\ <= \$v7397\;
      \$v7289%next\ <= \$v7289\;
      \$v7194%next\ <= \$v7194\;
      \$17874_w%next\ <= \$17874_w\;
      \$18844%next\ <= \$18844\;
      \$15181_modulo6685888_arg%next\ <= \$15181_modulo6685888_arg\;
      \$18175_w%next\ <= \$18175_w\;
      \$v5876%next\ <= \$v5876\;
      \$18676%next\ <= \$18676\;
      \$17539%next\ <= \$17539\;
      \$v7115%next\ <= \$v7115\;
      \$v6263%next\ <= \$v6263\;
      \$v6353%next\ <= \$v6353\;
      \$18335_w%next\ <= \$18335_w\;
      \$18993%next\ <= \$18993\;
      \$13928_w652_id%next\ <= \$13928_w652_id\;
      \$17504%next\ <= \$17504\;
      \$18046%next\ <= \$18046\;
      \$12670%next\ <= \$12670\;
      \$v5972%next\ <= \$v5972\;
      \$v6133%next\ <= \$v6133\;
      \$12743%next\ <= \$12743\;
      \$13539%next\ <= \$13539\;
      \$v5947%next\ <= \$v5947\;
      \$17117_v%next\ <= \$17117_v\;
      \$15173_modulo6685896_result%next\ <= \$15173_modulo6685896_result\;
      \$15819_v%next\ <= \$15819_v\;
      \$17547_copy_root_in_ram6635891_arg%next\ <= \$17547_copy_root_in_ram6635891_arg\;
      \$12681_wait662_id%next\ <= \$12681_wait662_id\;
      \$14043_v%next\ <= \$14043_v\;
      \$13814%next\ <= \$13814\;
      \$12803_loop666_arg%next\ <= \$12803_loop666_arg\;
      \$v6436%next\ <= \$v6436\;
      \$19136%next\ <= \$19136\;
      \$18674%next\ <= \$18674\;
      \$v6784%next\ <= \$v6784\;
      \$v7296%next\ <= \$v7296\;
      \$17395%next\ <= \$17395\;
      \$13236%next\ <= \$13236\;
      \$13464%next\ <= \$13464\;
      \$14051%next\ <= \$14051\;
      \$v7014%next\ <= \$v7014\;
      \$17320%next\ <= \$17320\;
      \$v7095%next\ <= \$v7095\;
      \$v6433%next\ <= \$v6433\;
      \$12681_wait662_result%next\ <= \$12681_wait662_result\;
      \$13383%next\ <= \$13383\;
      \$14578_v%next\ <= \$14578_v\;
      \$v7112%next\ <= \$v7112\;
      \$17675%next\ <= \$17675\;
      \$19127_w%next\ <= \$19127_w\;
      \$18808%next\ <= \$18808\;
      \$14148%next\ <= \$14148\;
      \$18705%next\ <= \$18705\;
      \$14804_binop_int6435903_id%next\ <= \$14804_binop_int6435903_id\;
      \$v6650%next\ <= \$v6650\;
      \$v7267%next\ <= \$v7267\;
      \$13624%next\ <= \$13624\;
      \$15588_modulo6685888_arg%next\ <= \$15588_modulo6685888_arg\;
      \$v7051%next\ <= \$v7051\;
      \$v5867%next\ <= \$v5867\;
      \$17388%next\ <= \$17388\;
      \$15173_modulo6685896_id%next\ <= \$15173_modulo6685896_id\;
      \$16589_compbranch6505927_result%next\ <= \$16589_compbranch6505927_result\;
      \$14069%next\ <= \$14069\;
      \$v6531%next\ <= \$v6531\;
      \$12713%next\ <= \$12713\;
      \$13021%next\ <= \$13021\;
      \$18666_next%next\ <= \$18666_next\;
      \$14446_v%next\ <= \$14446_v\;
      \$17677%next\ <= \$17677\;
      \$18740%next\ <= \$18740\;
      \$18842%next\ <= \$18842\;
      \$17972%next\ <= \$17972\;
      \$14989_modulo6685895_id%next\ <= \$14989_modulo6685895_id\;
      \$17598%next\ <= \$17598\;
      \$12522_wait662_id%next\ <= \$12522_wait662_id\;
      \$18701%next\ <= \$18701\;
      \$16662_fill6535928_arg%next\ <= \$16662_fill6535928_arg\;
      \$17490_next%next\ <= \$17490_next\;
      \$v6759%next\ <= \$v6759\;
      \$16928_compbranch6505934_arg%next\ <= \$16928_compbranch6505934_arg\;
      \$18922%next\ <= \$18922\;
      \$18464_hd%next\ <= \$18464_hd\;
      \$16963_compbranch6505935_result%next\ <= \$16963_compbranch6505935_result\;
      \$13992_v%next\ <= \$13992_v\;
      \$15508_modulo6685888_arg%next\ <= \$15508_modulo6685888_arg\;
      \$12929_hd%next\ <= \$12929_hd\;
      \$v7457%next\ <= \$v7457\;
      \$13538%next\ <= \$13538\;
      \$16457%next\ <= \$16457\;
      \$15306_r%next\ <= \$15306_r\;
      \$v6705%next\ <= \$v6705\;
      \$18122%next\ <= \$18122\;
      \$v7102%next\ <= \$v7102\;
      \$19143%next\ <= \$19143\;
      \$18670_next%next\ <= \$18670_next\;
      \$18634_aux664_arg%next\ <= \$18634_aux664_arg\;
      \$18793_copy_root_in_ram6635879_id%next\ <= \$18793_copy_root_in_ram6635879_id\;
      \$15149_modulo6685895_id%next\ <= \$15149_modulo6685895_id\;
      \$16788_compbranch6505930_result%next\ <= \$16788_compbranch6505930_result\;
      \$13535%next\ <= \$13535\;
      \$15545_v%next\ <= \$15545_v\;
      \$17482%next\ <= \$17482\;
      \$v7061%next\ <= \$v7061\;
      \$v6253%next\ <= \$v6253\;
      \$13897%next\ <= \$13897\;
      \$18735%next\ <= \$18735\;
      \$v7126%next\ <= \$v7126\;
      \$18281%next\ <= \$18281\;
      \$16473%next\ <= \$16473\;
      \$14917_modulo6685888_result%next\ <= \$14917_modulo6685888_result\;
      \$16741%next\ <= \$16741\;
      \$16510_forever6705925_arg%next\ <= \$16510_forever6705925_arg\;
      \$v6536%next\ <= \$v6536\;
      \$12811%next\ <= \$12811\;
      \$v6796%next\ <= \$v6796\;
      \$18459_w%next\ <= \$18459_w\;
      \$14413_v%next\ <= \$14413_v\;
      \$12520_loop666_result%next\ <= \$12520_loop666_result\;
      \$16612_compare6445898_id%next\ <= \$16612_compare6445898_id\;
      \$17747%next\ <= \$17747\;
      \$v7104%next\ <= \$v7104\;
      \$13939%next\ <= \$13939\;
      \$15661_binop_compare6455917_id%next\ <= \$15661_binop_compare6455917_id\;
      \$17973%next\ <= \$17973\;
      \$12804_loop665_id%next\ <= \$12804_loop665_id\;
      \$17758%next\ <= \$17758\;
      \$12719%next\ <= \$12719\;
      \$15397_modulo6685888_id%next\ <= \$15397_modulo6685888_id\;
      \$17105_w06555936_arg%next\ <= \$17105_w06555936_arg\;
      \$12792%next\ <= \$12792\;
      \$16194%next\ <= \$16194\;
      \$v7176%next\ <= \$v7176\;
      \$14829_modulo6685895_arg%next\ <= \$14829_modulo6685895_arg\;
      \$18049%next\ <= \$18049\;
      \$13536%next\ <= \$13536\;
      \$12842%next\ <= \$12842\;
      \$v7182%next\ <= \$v7182\;
      \$v6511%next\ <= \$v6511\;
      \$14693_modulo6685896_id%next\ <= \$14693_modulo6685896_id\;
      \$13023%next\ <= \$13023\;
      \$v6098%next\ <= \$v6098\;
      \$15792_compare6445897_arg%next\ <= \$15792_compare6445897_arg\;
      \$v6905%next\ <= \$v6905\;
      \$13313%next\ <= \$13313\;
      \$14552%next\ <= \$14552\;
      \$16840_b%next\ <= \$16840_b\;
      \$16568_b%next\ <= \$16568_b\;
      \$14423_v%next\ <= \$14423_v\;
      \$v6527%next\ <= \$v6527\;
      \$18262%next\ <= \$18262\;
      \$13078_copy_root_in_ram6635885_result%next\ <= \$13078_copy_root_in_ram6635885_result\;
      \$18351%next\ <= \$18351\;
      \$16232%next\ <= \$16232\;
      \$16133%next\ <= \$16133\;
      \$15711_v%next\ <= \$15711_v\;
      \$15614_forever6705914_id%next\ <= \$15614_forever6705914_id\;
      \$13004_w%next\ <= \$13004_w\;
      \$12803_loop666_id%next\ <= \$12803_loop666_id\;
      \$12744%next\ <= \$12744\;
      \$13311%next\ <= \$13311\;
      \$18664_next%next\ <= \$18664_next\;
      \$19264%next\ <= \$19264\;
      \$13472_next%next\ <= \$13472_next\;
      \$16858_compbranch6505932_id%next\ <= \$16858_compbranch6505932_id\;
      \$v7096%next\ <= \$v7096\;
      \$17966%next\ <= \$17966\;
      \$v6787%next\ <= \$v6787\;
      \$17459_loop665_result%next\ <= \$17459_loop665_result\;
      \$v7120%next\ <= \$v7120\;
      \$17310%next\ <= \$17310\;
      \$17492_next%next\ <= \$17492_next\;
      \$v6045%next\ <= \$v6045\;
      \$17748%next\ <= \$17748\;
      \$18638%next\ <= \$18638\;
      \$15792_compare6445897_id%next\ <= \$15792_compare6445897_id\;
      \$13963%next\ <= \$13963\;
      \$v6140%next\ <= \$v6140\;
      \$12933%next\ <= \$12933\;
      \$18640%next\ <= \$18640\;
      \$13528%next\ <= \$13528\;
      \$v7254%next\ <= \$v7254\;
      \$16881_compare6445898_id%next\ <= \$16881_compare6445898_id\;
      \$17460_aux664_arg%next\ <= \$17460_aux664_arg\;
      \$12523_make_block579_result%next\ <= \$12523_make_block579_result\;
      \$13922_wait662_arg%next\ <= \$13922_wait662_arg\;
      \$v6156%next\ <= \$v6156\;
      \$v6814%next\ <= \$v6814\;
      \$v7419%next\ <= \$v7419\;
      \$15451_binop_int6435912_result%next\ <= \$15451_binop_int6435912_result\;
      \$v6322%next\ <= \$v6322\;
      \$17331_sp%next\ <= \$17331_sp\;
      \$17894%next\ <= \$17894\;
      \$v6002%next\ <= \$v6002\;
      \$v6476%next\ <= \$v6476\;
      \$13239%next\ <= \$13239\;
      \$12708%next\ <= \$12708\;
      \$18812%next\ <= \$18812\;
      \$v6187%next\ <= \$v6187\;
      \$v7072%next\ <= \$v7072\;
      \rdy6148%next\ <= rdy6148;
      \$18047%next\ <= \$18047\;
      \$14644_binop_int6435901_id%next\ <= \$14644_binop_int6435901_id\;
      \$14597_modulo6685888_id%next\ <= \$14597_modulo6685888_id\;
      \$v7103%next\ <= \$v7103\;
      \$19261%next\ <= \$19261\;
      \$16893_compbranch6505933_arg%next\ <= \$16893_compbranch6505933_arg\;
      \$13390%next\ <= \$13390\;
      \$16534%next\ <= \$16534\;
      \$v7191%next\ <= \$v7191\;
      \$19002%next\ <= \$19002\;
      \$v7041%next\ <= \$v7041\;
      \$v6968%next\ <= \$v6968\;
      \$v7127%next\ <= \$v7127\;
      \$17520_copy_root_in_ram6635893_result%next\ <= \$17520_copy_root_in_ram6635893_result\;
      \$v6332%next\ <= \$v6332\;
      \$13229%next\ <= \$13229\;
      \$v6159%next\ <= \$v6159\;
      \$15684_compare6445897_id%next\ <= \$15684_compare6445897_id\;
      \$v7114%next\ <= \$v7114\;
      \$17544%next\ <= \$17544\;
      \$v6704%next\ <= \$v6704\;
      \$18040%next\ <= \$18040\;
      \$17786%next\ <= \$17786\;
      \$v7233%next\ <= \$v7233\;
      \$14207_loop_push6495899_arg%next\ <= \$14207_loop_push6495899_arg\;
      \$16709%next\ <= \$16709\;
      \$v7113%next\ <= \$v7113\;
      \$14724_binop_int6435902_arg%next\ <= \$14724_binop_int6435902_arg\;
      \$13232%next\ <= \$13232\;
      \$16986_compare6445898_arg%next\ <= \$16986_compare6445898_arg\;
      \$v6054%next\ <= \$v6054\;
      \$16074_v%next\ <= \$16074_v\;
      \$v6781%next\ <= \$v6781\;
      \$v7047%next\ <= \$v7047\;
      \$17503%next\ <= \$17503\;
      \$13147%next\ <= \$13147\;
      \$v6259%next\ <= \$v6259\;
      \$v6144%next\ <= \$v6144\;
      \$13018%next\ <= \$13018\;
      \$v6603%next\ <= \$v6603\;
      \$14016_v%next\ <= \$14016_v\;
      \$16752_fill6545929_id%next\ <= \$16752_fill6545929_id\;
      \$v5973%next\ <= \$v5973\;
      \$13815%next\ <= \$13815\;
      \$v7033%next\ <= \$v7033\;
      \$v5983%next\ <= \$v5983\;
      \$19271%next\ <= \$19271\;
      \$v6735%next\ <= \$v6735\;
      \$v6769%next\ <= \$v6769\;
      \$v7242%next\ <= \$v7242\;
      \$16508%next\ <= \$16508\;
      \$12808_aux664_arg%next\ <= \$12808_aux664_arg\;
      \$18708%next\ <= \$18708\;
      \$18991%next\ <= \$18991\;
      \$14471%next\ <= \$14471\;
      \$v7070%next\ <= \$v7070\;
      \$12547%next\ <= \$12547\;
      \$v7031%next\ <= \$v7031\;
      \$v6315%next\ <= \$v6315\;
      \$12674%next\ <= \$12674\;
      \$12846%next\ <= \$12846\;
      \$17010%next\ <= \$17010\;
      \$17560%next\ <= \$17560\;
      \$16156%next\ <= \$16156\;
      \$15021_modulo6685888_id%next\ <= \$15021_modulo6685888_id\;
      \$13925_offsetclosure_n639_arg%next\ <= \$13925_offsetclosure_n639_arg\;
      \$14898_v%next\ <= \$14898_v\;
      \$14693_modulo6685896_result%next\ <= \$14693_modulo6685896_result\;
      \$15497_r%next\ <= \$15497_r\;
      \$13105_copy_root_in_ram6635884_id%next\ <= \$13105_copy_root_in_ram6635884_id\;
      \$17434%next\ <= \$17434\;
      \$16515%next\ <= \$16515\;
      \$14512_v%next\ <= \$14512_v\;
      \$14300_v%next\ <= \$14300_v\;
      \$18261%next\ <= \$18261\;
      \$17207_arg%next\ <= \$17207_arg\;
      \$13315%next\ <= \$13315\;
      \$18992%next\ <= \$18992\;
      \$18344%next\ <= \$18344\;
      \$17183%next\ <= \$17183\;
      \$v7032%next\ <= \$v7032\;
      \result6112%next\ <= result6112;
      \$v5960%next\ <= \$v5960\;
      \$v7084%next\ <= \$v7084\;
      \$v6639%next\ <= \$v6639\;
      \$v7060%next\ <= \$v7060\;
      \$18030_w%next\ <= \$18030_w\;
      \$18190%next\ <= \$18190\;
      \$16380_v%next\ <= \$16380_v\;
      \$v6295%next\ <= \$v6295\;
      \$18924%next\ <= \$18924\;
      \$12659%next\ <= \$12659\;
      \$v6111%next\ <= \$v6111\;
      \$v6011%next\ <= \$v6011\;
      \$12891_copy_root_in_ram6635884_result%next\ <= \$12891_copy_root_in_ram6635884_result\;
      \$18621%next\ <= \$18621\;
      \$14185_next_env%next\ <= \$14185_next_env\;
      \$17166%next\ <= \$17166\;
      \$v6059%next\ <= \$v6059\;
      \$12703%next\ <= \$12703\;
      \$v6358%next\ <= \$v6358\;
      \$12832%next\ <= \$12832\;
      \$15684_compare6445897_result%next\ <= \$15684_compare6445897_result\;
      \$v7111%next\ <= \$v7111\;
      \$17895%next\ <= \$17895\;
      \$13812%next\ <= \$13812\;
      \$18632_loop666_id%next\ <= \$18632_loop666_id\;
      \$17952_w%next\ <= \$17952_w\;
      \$13820%next\ <= \$13820\;
      \$13533%next\ <= \$13533\;
      \$15805_binop_compare6455921_result%next\ <= \$15805_binop_compare6455921_result\;
      \$15413_modulo6685896_id%next\ <= \$15413_modulo6685896_id\;
      \$13977_v%next\ <= \$13977_v\;
      \$v6294%next\ <= \$v6294\;
      \$12857_forever6705883_id%next\ <= \$12857_forever6705883_id\;
      \$v7438%next\ <= \$v7438\;
      \$v7082%next\ <= \$v7082\;
      \$v6415%next\ <= \$v6415\;
      \$v5982%next\ <= \$v5982\;
      \$19265%next\ <= \$19265\;
      \$17011%next\ <= \$17011\;
      \$v7012%next\ <= \$v7012\;
      \$17505_forever6705894_id%next\ <= \$17505_forever6705894_id\;
      \$v7282%next\ <= \$v7282\;
      \$12813%next\ <= \$12813\;
      \$17499%next\ <= \$17499\;
      \$v6457%next\ <= \$v6457\;
      \$13150%next\ <= \$13150\;
      \$17808%next\ <= \$17808\;
      \$v6820%next\ <= \$v6820\;
      \$17970%next\ <= \$17970\;
      \$12803_loop666_result%next\ <= \$12803_loop666_result\;
      \$v7276%next\ <= \$v7276\;
      \$14964_binop_int6435905_result%next\ <= \$14964_binop_int6435905_result\;
      \$v7134%next\ <= \$v7134\;
      \$17809%next\ <= \$17809\;
      \$16404%next\ <= \$16404\;
      \$v7157%next\ <= \$v7157\;
      \$17969%next\ <= \$17969\;
      \$v6280%next\ <= \$v6280\;
      \$12845%next\ <= \$12845\;
      \$v6361%next\ <= \$v6361\;
      \$12561%next\ <= \$12561\;
      \$17545%next\ <= \$17545\;
      \$18634_aux664_id%next\ <= \$18634_aux664_id\;
      \$15410_r%next\ <= \$15410_r\;
      \$v6582%next\ <= \$v6582\;
      \$v6600%next\ <= \$v6600\;
      \$15062_res%next\ <= \$15062_res\;
      \$v6264%next\ <= \$v6264\;
      \$14342%next\ <= \$14342\;
      \$v6691%next\ <= \$v6691\;
      \$12562%next\ <= \$12562\;
      \result5939%next\ <= result5939;
      \$12657%next\ <= \$12657\;
      \$v7130%next\ <= \$v7130\;
      \$16193%next\ <= \$16193\;
      \$16916_compare6445898_result%next\ <= \$16916_compare6445898_result\;
      \$18839%next\ <= \$18839\;
      \$13787%next\ <= \$13787\;
      \$v7303%next\ <= \$v7303\;
      \$19146%next\ <= \$19146\;
      \$15684_compare6445897_arg%next\ <= \$15684_compare6445897_arg\;
      \$15142_res%next\ <= \$15142_res\;
      \$12905%next\ <= \$12905\;
      \$v6267%next\ <= \$v6267\;
      \$18658%next\ <= \$18658\;
      \$13386%next\ <= \$13386\;
      \$17465%next\ <= \$17465\;
      \$v6477%next\ <= \$v6477\;
      \$13025%next\ <= \$13025\;
      \$18678%next\ <= \$18678\;
      \$16461%next\ <= \$16461\;
      \$v6774%next\ <= \$v6774\;
      \$18180_hd%next\ <= \$18180_hd\;
      \$v6811%next\ <= \$v6811\;
      \$13791%next\ <= \$13791\;
      \$14464_v%next\ <= \$14464_v\;
      \$15851_argument1%next\ <= \$15851_argument1\;
      \$13022%next\ <= \$13022\;
      \$15101_modulo6685888_arg%next\ <= \$15101_modulo6685888_arg\;
      \$13124%next\ <= \$13124\;
      \$v6762%next\ <= \$v6762\;
      \$v6720%next\ <= \$v6720\;
      \$v6528%next\ <= \$v6528\;
      \$v6083%next\ <= \$v6083\;
      \$16724%next\ <= \$16724\;
      \$v6524%next\ <= \$v6524\;
      \$v6448%next\ <= \$v6448\;
      \$17184%next\ <= \$17184\;
      \$13228%next\ <= \$13228\;
      \$19139%next\ <= \$19139\;
      \$v7036%next\ <= \$v7036\;
      \$v6755%next\ <= \$v6755\;
      \$17533%next\ <= \$17533\;
      \result5974%next\ <= result5974;
      \$v7037%next\ <= \$v7037\;
      \$18589%next\ <= \$18589\;
      \$14669_modulo6685895_result%next\ <= \$14669_modulo6685895_result\;
      \$13813%next\ <= \$13813\;
      \$17105_w06555936_result%next\ <= \$17105_w06555936_result\;
      \$13921_loop665_arg%next\ <= \$13921_loop665_arg\;
      \$17599%next\ <= \$17599\;
      \$13921_loop665_result%next\ <= \$13921_loop665_result\;
      \$v7401%next\ <= \$v7401\;
      \$v6980%next\ <= \$v6980\;
      \$16337%next\ <= \$16337\;
      \$17534%next\ <= \$17534\;
      \$12558%next\ <= \$12558\;
      \$v6926%next\ <= \$v6926\;
      \$16811_compare6445898_id%next\ <= \$16811_compare6445898_id\;
      \$v5989%next\ <= \$v5989\;
      \$14103%next\ <= \$14103\;
      \$15556_modulo6685895_arg%next\ <= \$15556_modulo6685895_arg\;
      \$19147%next\ <= \$19147\;
      \$16383%next\ <= \$16383\;
      \$v7149%next\ <= \$v7149\;
      \$13314%next\ <= \$13314\;
      \$15639_v%next\ <= \$15639_v\;
      \$16624_argument2%next\ <= \$16624_argument2\;
      \$15069_modulo6685895_result%next\ <= \$15069_modulo6685895_result\;
      \$16662_fill6535928_id%next\ <= \$16662_fill6535928_id\;
      \rdy6113%next\ <= rdy6113;
      \$17542%next\ <= \$17542\;
      \$v6345%next\ <= \$v6345\;
      \$v6194%next\ <= \$v6194\;
      \$v6571%next\ <= \$v6571\;
      \$15531_binop_int6435913_result%next\ <= \$15531_binop_int6435913_result\;
      \$v6439%next\ <= \$v6439\;
      \$v6079%next\ <= \$v6079\;
      \$15621_forever6705915_arg%next\ <= \$15621_forever6705915_arg\;
      \$17884%next\ <= \$17884\;
      \$v7097%next\ <= \$v7097\;
      \$13927_branch_if648_id%next\ <= \$13927_branch_if648_id\;
      \$14982_res%next\ <= \$14982_res\;
      \$18353%next\ <= \$18353\;
      \$v7347%next\ <= \$v7347\;
      \$16846_compare6445898_arg%next\ <= \$16846_compare6445898_arg\;
      \$v6895%next\ <= \$v6895\;
      \$16195_forever6705924_arg%next\ <= \$16195_forever6705924_arg\;
      \$17589%next\ <= \$17589\;
      \$13017%next\ <= \$13017\;
      \$15747_v%next\ <= \$15747_v\;
      \$16662_fill6535928_result%next\ <= \$16662_fill6535928_result\;
      \$18345%next\ <= \$18345\;
      \$v7122%next\ <= \$v7122\;
      \$17048_w16565937_id%next\ <= \$17048_w16565937_id\;
      \$18686_copy_root_in_ram6635880_result%next\ <= \$18686_copy_root_in_ram6635880_result\;
      \$15093_modulo6685896_id%next\ <= \$15093_modulo6685896_id\;
      \$18736%next\ <= \$18736\;
      \$18671%next\ <= \$18671\;
      \$15500_modulo6685896_id%next\ <= \$15500_modulo6685896_id\;
      \$v7226%next\ <= \$v7226\;
      \$17459_loop665_id%next\ <= \$17459_loop665_id\;
      \$15333_modulo6685896_arg%next\ <= \$15333_modulo6685896_arg\;
      \$17807%next\ <= \$17807\;
      \$v6220%next\ <= \$v6220\;
      \$13821%next\ <= \$13821\;
      \$18035_hd%next\ <= \$18035_hd\;
      \$v6290%next\ <= \$v6290\;
      \$17172%next\ <= \$17172\;
      \$13394%next\ <= \$13394\;
      \$19338%next\ <= \$19338\;
      \$17368_v%next\ <= \$17368_v\;
      \$v5871%next\ <= \$v5871\;
      \$13958%next\ <= \$13958\;
      \$12824%next\ <= \$12824\;
      \$17562%next\ <= \$17562\;
      \$16322%next\ <= \$16322\;
      \$v7105%next\ <= \$v7105\;
      \$13698%next\ <= \$13698\;
      \$17520_copy_root_in_ram6635893_arg%next\ <= \$17520_copy_root_in_ram6635893_arg\;
      \$15556_modulo6685895_id%next\ <= \$15556_modulo6685895_id\;
      \$13105_copy_root_in_ram6635884_result%next\ <= \$13105_copy_root_in_ram6635884_result\;
      \$12891_copy_root_in_ram6635884_id%next\ <= \$12891_copy_root_in_ram6635884_id\;
      \$12806_loop666_arg%next\ <= \$12806_loop666_arg\;
      \$v6566%next\ <= \$v6566\;
      \$15181_modulo6685888_id%next\ <= \$15181_modulo6685888_id\;
      \$v7080%next\ <= \$v7080\;
      \$v6675%next\ <= \$v6675\;
      \$v6576%next\ <= \$v6576\;
      \$16998_argument3%next\ <= \$16998_argument3\;
      \$v7423%next\ <= \$v7423\;
      \$18728%next\ <= \$18728\;
      \$16157%next\ <= \$16157\;
      \$13684_hd%next\ <= \$13684_hd\;
      \$19111%next\ <= \$19111\;
      \$v6647%next\ <= \$v6647\;
      \$13091%next\ <= \$13091\;
      \$13143_hd%next\ <= \$13143_hd\;
      \$18793_copy_root_in_ram6635879_result%next\ <= \$18793_copy_root_in_ram6635879_result\;
      \$15769_binop_compare6455920_result%next\ <= \$15769_binop_compare6455920_result\;
      \$16462%next\ <= \$16462\;
      \$14265%next\ <= \$14265\;
      \$12916%next\ <= \$12916\;
      \$v6244%next\ <= \$v6244\;
      \$12742%next\ <= \$12742\;
      \$13119%next\ <= \$13119\;
      \$13972_v%next\ <= \$13972_v\;
      \$14884_binop_int6435904_result%next\ <= \$14884_binop_int6435904_result\;
      \$13951%next\ <= \$13951\;
      \$v7024%next\ <= \$v7024\;
      \$13923_make_block579_arg%next\ <= \$13923_make_block579_arg\;
      \$15648_compare6445897_result%next\ <= \$15648_compare6445897_result\;
      \$17330_sp%next\ <= \$17330_sp\;
      \$v6620%next\ <= \$v6620\;
      \$17353%next\ <= \$17353\;
      \$v6983%next\ <= \$v6983\;
      \$v7257%next\ <= \$v7257\;
      \$v6663%next\ <= \$v6663\;
      \$13118%next\ <= \$13118\;
      \$v6032%next\ <= \$v6032\;
      \$18672%next\ <= \$18672\;
      \$19074%next\ <= \$19074\;
      \$15309_modulo6685895_id%next\ <= \$15309_modulo6685895_id\;
      \$v6260%next\ <= \$v6260\;
      \$19076%next\ <= \$19076\;
      \rdy5975%next\ <= rdy5975;
      \$15124_binop_int6435907_result%next\ <= \$15124_binop_int6435907_result\;
      \$16334_v%next\ <= \$16334_v\;
      \$v7270%next\ <= \$v7270\;
      \$18042%next\ <= \$18042\;
      \$18611%next\ <= \$18611\;
      \$14377_v%next\ <= \$14377_v\;
      \$16381_v%next\ <= \$16381_v\;
      \$v6076%next\ <= \$v6076\;
      \$15908%next\ <= \$15908\;
      \$12563%next\ <= \$12563\;
      \$v7026%next\ <= \$v7026\;
      \$v6698%next\ <= \$v6698\;
      \$15013_modulo6685896_result%next\ <= \$15013_modulo6685896_result\;
      \$12805_aux664_arg%next\ <= \$12805_aux664_arg\;
      \$v7075%next\ <= \$v7075\;
      \$13024%next\ <= \$13024\;
      \$13965%next\ <= \$13965\;
      \$18573%next\ <= \$18573\;
      \$v6124%next\ <= \$v6124\;
      \$17481%next\ <= \$17481\;
      \$v6215%next\ <= \$v6215\;
      \$15720_compare6445897_result%next\ <= \$15720_compare6445897_result\;
      \$v7160%next\ <= \$v7160\;
      \$v6497%next\ <= \$v6497\;
      \$15044_binop_int6435906_arg%next\ <= \$15044_binop_int6435906_arg\;
      \$13097%next\ <= \$13097\;
      \$17456_loop665_arg%next\ <= \$17456_loop665_arg\;
      \$13952%next\ <= \$13952\;
      \$15093_modulo6685896_result%next\ <= \$15093_modulo6685896_result\;
      \$13924_apply638_id%next\ <= \$13924_apply638_id\;
      \$v6556%next\ <= \$v6556\;
      \$14701_modulo6685888_id%next\ <= \$14701_modulo6685888_id\;
      \$12687%next\ <= \$12687\;
      \$15473_r%next\ <= \$15473_r\;
      \$17061%next\ <= \$17061\;
      \$16725%next\ <= \$16725\;
      \$v6412%next\ <= \$v6412\;
      \$v7407%next\ <= \$v7407\;
      \$v6747%next\ <= \$v6747\;
      \$12831%next\ <= \$12831\;
      \$16651%next\ <= \$16651\;
      \$14781_modulo6685888_id%next\ <= \$14781_modulo6685888_id\;
      \$16658%next\ <= \$16658\;
      \$v7136%next\ <= \$v7136\;
      \$14589_modulo6685895_id%next\ <= \$14589_modulo6685895_id\;
      \$v5968%next\ <= \$v5968\;
      \$v6339%next\ <= \$v6339\;
      \$16788_compbranch6505930_id%next\ <= \$16788_compbranch6505930_id\;
      \$17486%next\ <= \$17486\;
      \$v6331%next\ <= \$v6331\;
      \$18553%next\ <= \$18553\;
      \$14034_v%next\ <= \$14034_v\;
      \$v7410%next\ <= \$v7410\;
      \$v7131%next\ <= \$v7131\;
      \$18284%next\ <= \$18284\;
      \$v7390%next\ <= \$v7390\;
      \$13306%next\ <= \$13306\;
      \$v6539%next\ <= \$v6539\;
      \$v7341%next\ <= \$v7341\;
      \$15090_r%next\ <= \$15090_r\;
      \$14906_r%next\ <= \$14906_r\;
      \$13462%next\ <= \$13462\;
      \$19270%next\ <= \$19270\;
      \$v6850%next\ <= \$v6850\;
      \$v7430%next\ <= \$v7430\;
      \$v6671%next\ <= \$v6671\;
      \$15149_modulo6685895_result%next\ <= \$15149_modulo6685895_result\;
      \$15756_compare6445897_id%next\ <= \$15756_compare6445897_id\;
      \$v6418%next\ <= \$v6418\;
      \$v6250%next\ <= \$v6250\;
      \$v6051%next\ <= \$v6051\;
      \$15621_forever6705915_id%next\ <= \$15621_forever6705915_id\;
      \$v6886%next\ <= \$v6886\;
      \$16858_compbranch6505932_result%next\ <= \$16858_compbranch6505932_result\;
      \$15222_res%next\ <= \$15222_res\;
      \$v6770%next\ <= \$v6770\;
      \$v7040%next\ <= \$v7040\;
      \$16301%next\ <= \$16301\;
      \$13911%next\ <= \$13911\;
      \$17680%next\ <= \$17680\;
      \$v6191%next\ <= \$v6191\;
      \$15138_v%next\ <= \$15138_v\;
      \$v6486%next\ <= \$v6486\;
      \$13152%next\ <= \$13152\;
      \$16155%next\ <= \$16155\;
      \$14933_modulo6685896_arg%next\ <= \$14933_modulo6685896_arg\;
      \$12693%next\ <= \$12693\;
      \$v7106%next\ <= \$v7106\;
      \$v7067%next\ <= \$v7067\;
      \$13920_loop666_result%next\ <= \$13920_loop666_result\;
      \$16293%next\ <= \$16293\;
      \$13159%next\ <= \$13159\;
      \$13953%next\ <= \$13953\;
      \$15625_binop_compare6455916_arg%next\ <= \$15625_binop_compare6455916_arg\;
      \$13015%next\ <= \$13015\;
      \$17799_hd%next\ <= \$17799_hd\;
      \$v6039%next\ <= \$v6039\;
      \$15611%next\ <= \$15611\;
      \$v6808%next\ <= \$v6808\;
      \$17444%next\ <= \$17444\;
      \$14853_modulo6685896_id%next\ <= \$14853_modulo6685896_id\;
      \$18665%next\ <= \$18665\;
      \$19132_hd%next\ <= \$19132_hd\;
      \$16313_v%next\ <= \$16313_v\;
      \$14757_modulo6685888_arg%next\ <= \$14757_modulo6685888_arg\;
      \$18710%next\ <= \$18710\;
      \$v5979%next\ <= \$v5979\;
      \$v6006%next\ <= \$v6006\;
      \$14621_modulo6685888_id%next\ <= \$14621_modulo6685888_id\;
      \$14941_modulo6685888_id%next\ <= \$14941_modulo6685888_id\;
      \$19073%next\ <= \$19073\;
      \$15733_binop_compare6455919_id%next\ <= \$15733_binop_compare6455919_id\;
      \$15620%next\ <= \$15620\;
      \$17596%next\ <= \$17596\;
      \$16413%next\ <= \$16413\;
      \$19141%next\ <= \$19141\;
      \$17753%next\ <= \$17753\;
      \$16706%next\ <= \$16706\;
      \$16296%next\ <= \$16296\;
      \$v7001%next\ <= \$v7001\;
      \$18468%next\ <= \$18468\;
      \$19000%next\ <= \$19000\;
      \$v5877%next\ <= \$v5877\;
      \$16951_compare6445898_id%next\ <= \$16951_compare6445898_id\;
      \$13231%next\ <= \$13231\;
      \$v6024%next\ <= \$v6024\;
      \$13130%next\ <= \$13130\;
      \$15469_res%next\ <= \$15469_res\;
      \$18471%next\ <= \$18471\;
      \$v6793%next\ <= \$v6793\;
      \$v7266%next\ <= \$v7266\;
      \$18350%next\ <= \$18350\;
      \$16357%next\ <= \$16357\;
      \$15149_modulo6685895_arg%next\ <= \$15149_modulo6685895_arg\;
      \$13987_v%next\ <= \$13987_v\;
      \$v7055%next\ <= \$v7055\;
      \$17483%next\ <= \$17483\;
      \$14260%next\ <= \$14260\;
      \$15588_modulo6685888_id%next\ <= \$15588_modulo6685888_id\;
      \$v7309%next\ <= \$v7309\;
      \$15643_res%next\ <= \$15643_res\;
      \$13078_copy_root_in_ram6635885_arg%next\ <= \$13078_copy_root_in_ram6635885_arg\;
      \$18914%next\ <= \$18914\;
      \$17660_w%next\ <= \$17660_w\;
      \$16846_compare6445898_result%next\ <= \$16846_compare6445898_result\;
      \$18817%next\ <= \$18817\;
      \$v6871%next\ <= \$v6871\;
      \$17672%next\ <= \$17672\;
      \$19148%next\ <= \$19148\;
      \$v7329%next\ <= \$v7329\;
      \$19072%next\ <= \$19072\;
      \$15733_binop_compare6455919_result%next\ <= \$15733_binop_compare6455919_result\;
      \$14081%next\ <= \$14081\;
      \$18545%next\ <= \$18545\;
      \$13889%next\ <= \$13889\;
      \$14015%next\ <= \$14015\;
      \$12840_next%next\ <= \$12840_next\;
      \$18686_copy_root_in_ram6635880_arg%next\ <= \$18686_copy_root_in_ram6635880_arg\;
      \$14742_res%next\ <= \$14742_res\;
      \$14586_r%next\ <= \$14586_r\;
      \$18195%next\ <= \$18195\;
      \$v6540%next\ <= \$v6540\;
      \$18793_copy_root_in_ram6635879_arg%next\ <= \$18793_copy_root_in_ram6635879_arg\;
      \$15317_modulo6685888_id%next\ <= \$15317_modulo6685888_id\;
      \$16551_compbranch6505926_result%next\ <= \$16551_compbranch6505926_result\;
      \$17811%next\ <= \$17811\;
      \$16980_b%next\ <= \$16980_b\;
      \$18349%next\ <= \$18349\;
      \$15451_binop_int6435912_id%next\ <= \$15451_binop_int6435912_id\;
      \$14002_v%next\ <= \$14002_v\;
      \$14997_modulo6685888_arg%next\ <= \$14997_modulo6685888_arg\;
      \$16335_v%next\ <= \$16335_v\;
      \$13014%next\ <= \$13014\;
      \$v6977%next\ <= \$v6977\;
      \$18039%next\ <= \$18039\;
      \$13448%next\ <= \$13448\;
      \$17571%next\ <= \$17571\;
      \$17757%next\ <= \$17757\;
      \$v6018%next\ <= \$v6018\;
      \$16358%next\ <= \$16358\;
      \$v7052%next\ <= \$v7052\;
      \$17352%next\ <= \$17352\;
      \$17756%next\ <= \$17756\;
      \$v6141%next\ <= \$v6141\;
      \$13391%next\ <= \$13391\;
      \$v6086%next\ <= \$v6086\;
      \$v6145%next\ <= \$v6145\;
      \$15066_r%next\ <= \$15066_r\;
      \result6147%next\ <= result6147;
      \$15446%next\ <= \$15446\;
      \$v6877%next\ <= \$v6877\;
      \$16041_v%next\ <= \$16041_v\;
      \$16063_w6515922_arg%next\ <= \$16063_w6515922_arg\;
      \$12700%next\ <= \$12700\;
      \$16951_compare6445898_result%next\ <= \$16951_compare6445898_result\;
      \$v6210%next\ <= \$v6210\;
      \$15564_modulo6685888_id%next\ <= \$15564_modulo6685888_id\;
      \$12721%next\ <= \$12721\;
      \$18920%next\ <= \$18920\;
      \$14393_hd%next\ <= \$14393_hd\;
      \$18282%next\ <= \$18282\;
      \$v7141%next\ <= \$v7141\;
      \$15157_modulo6685888_result%next\ <= \$15157_modulo6685888_result\;
      \$14850_r%next\ <= \$14850_r\;
      \$17601%next\ <= \$17601\;
      \$v6310%next\ <= \$v6310\;
      \$14493_v%next\ <= \$14493_v\;
      \$12711%next\ <= \$12711\;
      \$v5864%next\ <= \$v5864\;
      \$v6483%next\ <= \$v6483\;
      \$13819%next\ <= \$13819\;
      \$v7325%next\ <= \$v7325\;
      \$13120%next\ <= \$13120\;
      \$v7087%next\ <= \$v7087\;
      \$v6615%next\ <= \$v6615\;
      \$15146_r%next\ <= \$15146_r\;
      \$v7394%next\ <= \$v7394\;
      \$18347%next\ <= \$18347\;
      \$18700%next\ <= \$18700\;
      \$v6777%next\ <= \$v6777\;
      \$12940%next\ <= \$12940\;
      \$v7173%next\ <= \$v7173\;
      \$17062%next\ <= \$17062\;
      \$v7073%next\ <= \$v7073\;
      \$14025_v%next\ <= \$14025_v\;
      \$14561%next\ <= \$14561\;
      \$16437_v%next\ <= \$16437_v\;
      \$15549_res%next\ <= \$15549_res\;
      \$15253_modulo6685896_arg%next\ <= \$15253_modulo6685896_arg\;
      \$15013_modulo6685896_arg%next\ <= \$15013_modulo6685896_arg\;
      \$14822_res%next\ <= \$14822_res\;
      \$18847%next\ <= \$18847\;
      \$18840%next\ <= \$18840\;
      \$18340_hd%next\ <= \$18340_hd\;
      \$v7148%next\ <= \$v7148\;
      \$14884_binop_int6435904_id%next\ <= \$14884_binop_int6435904_id\;
      \$18632_loop666_result%next\ <= \$18632_loop666_result\;
      \$15226_r%next\ <= \$15226_r\;
      \$18422%next\ <= \$18422\;
      \$15444%next\ <= \$15444\;
      \$19137%next\ <= \$19137\;
      \$18923%next\ <= \$18923\;
      \$17161%next\ <= \$17161\;
      \$12662%next\ <= \$12662\;
      \$v7065%next\ <= \$v7065\;
      \$14662_res%next\ <= \$14662_res\;
      \$v6226%next\ <= \$v6226\;
      \$v7319%next\ <= \$v7319\;
      \$17396%next\ <= \$17396\;
      \$17806%next\ <= \$17806\;
      \$v6612%next\ <= \$v6612\;
      \$15805_binop_compare6455921_id%next\ <= \$15805_binop_compare6455921_id\;
      \$13305%next\ <= \$13305\;
      \$13230%next\ <= \$13230\;
      \$19056%next\ <= \$19056\;
      \$18469%next\ <= \$18469\;
      \$v7286%next\ <= \$v7286\;
      \$13534%next\ <= \$13534\;
      \$v7152%next\ <= \$v7152\;
      \$v6929%next\ <= \$v6929\;
      \$16910_b%next\ <= \$16910_b\;
      \$v7043%next\ <= \$v7043\;
      \$12850%next\ <= \$12850\;
      \$17456_loop665_id%next\ <= \$17456_loop665_id\;
      \$18477%next\ <= \$18477\;
      \$v7225%next\ <= \$v7225\;
      \$v6923%next\ <= \$v6923\;
      \$v6674%next\ <= \$v6674\;
      \$13699%next\ <= \$13699\;
      \$v6944%next\ <= \$v6944\;
      \$13923_make_block579_id%next\ <= \$13923_make_block579_id\;
      \$14207_loop_push6495899_id%next\ <= \$14207_loop_push6495899_id\;
      \$15648_compare6445897_arg%next\ <= \$15648_compare6445897_arg\;
      \$13803_w%next\ <= \$13803_w\;
      \$17780%next\ <= \$17780\;
      \$12876%next\ <= \$12876\;
      \$18656%next\ <= \$18656\;
      \$v6687%next\ <= \$v6687\;
      \$v6107%next\ <= \$v6107\;
      \$12661%next\ <= \$12661\;
      \$v6630%next\ <= \$v6630\;
      \$15697_binop_compare6455918_id%next\ <= \$15697_binop_compare6455918_id\;
      \$v7124%next\ <= \$v7124\;
      \$v7384%next\ <= \$v7384\;
      \$v7063%next\ <= \$v7063\;
      \$13928_w652_arg%next\ <= \$13928_w652_arg\;
      \$15465_v%next\ <= \$15465_v\;
      \$13622%next\ <= \$13622\;
      \$14355%next\ <= \$14355\;
      \$v7312%next\ <= \$v7312\;
      \$v6636%next\ <= \$v6636\;
      \$14770_r%next\ <= \$14770_r\;
      \$v6063%next\ <= \$v6063\;
      \$15013_modulo6685896_id%next\ <= \$15013_modulo6685896_id\;
      \$14690_r%next\ <= \$14690_r\;
      \$12807_loop665_arg%next\ <= \$12807_loop665_arg\;
      \$v6120%next\ <= \$v6120\;
      \$17810%next\ <= \$17810\;
      \$v6168%next\ <= \$v6168\;
      \$v7053%next\ <= \$v7053\;
      \$v7239%next\ <= \$v7239\;
      \$17236%next\ <= \$17236\;
      \$v7209%next\ <= \$v7209\;
      \$13128%next\ <= \$13128\;
      \$15229_modulo6685895_id%next\ <= \$15229_modulo6685895_id\;
      \$v7316%next\ <= \$v7316\;
      \$12690%next\ <= \$12690\;
      \$13925_offsetclosure_n639_id%next\ <= \$13925_offsetclosure_n639_id\;
      \$13020%next\ <= \$13020\;
      \$v6932%next\ <= \$v6932\;
      \$12539%next\ <= \$12539\;
      \$v6592%next\ <= \$v6592\;
      \$v6010%next\ <= \$v6010\;
      \$13093%next\ <= \$13093\;
      \$18323%next\ <= \$18323\;
      \$17965%next\ <= \$17965\;
      \$v5971%next\ <= \$v5971\;
      \$16659_sp%next\ <= \$16659_sp\;
      \$17547_copy_root_in_ram6635891_result%next\ <= \$17547_copy_root_in_ram6635891_result\;
      \$13690%next\ <= \$13690\;
      \$13628%next\ <= \$13628\;
      \$v6349%next\ <= \$v6349\;
      \$13465%next\ <= \$13465\;
      \$12812%next\ <= \$12812\;
      \$v6028%next\ <= \$v6028\;
      \$13374_w%next\ <= \$13374_w\;
      \$14368%next\ <= \$14368\;
      \$12718%next\ <= \$12718\;
      \$17784%next\ <= \$17784\;
      \$15508_modulo6685888_id%next\ <= \$15508_modulo6685888_id\;
      \$15364_binop_int6435910_result%next\ <= \$15364_binop_int6435910_result\;
      \$14613_modulo6685896_arg%next\ <= \$14613_modulo6685896_arg\;
      \$15751_res%next\ <= \$15751_res\;
      \$13537%next\ <= \$13537\;
      \$12654%next\ <= \$12654\;
      \$v7071%next\ <= \$v7071\;
      \$v6311%next\ <= \$v6311\;
      \$ram_lock%next\ <= \$ram_lock\;
      \$global_end_lock%next\ <= \$global_end_lock\;
      \$code_lock%next\ <= \$code_lock\;
      
      
      result <= result5939;
      end process;
  end architecture;
