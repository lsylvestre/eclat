-- code generated from the following source code:
--   ../ocaml-vm/vm/mlvalue.ecl
--   ../ocaml-vm/vm/fail.ecl
--   ../ocaml-vm/vm/ram.ecl
--   ../ocaml-vm/vm/runtime.ecl
--   ../ocaml-vm/vm/debug.ecl
--   ../ocaml-vm/vm/alloc.ecl
--   ../ocaml-vm/vm/prims.ecl
--   ../ocaml-vm/bytecode.ecl
--   ../ocaml-vm/vm/vm.ecl
--   ../ocaml-vm/vm/target-specific/intel-max10/IOs.ecl
--   ../ocaml-vm/vm/target-specific/intel-max10/main.ecl
--
-- with the following command:
--
--    ./eclat -arg ((true,true,true,true,true,true,true,true,true,true),(true,false)) ../ocaml-vm/vm/mlvalue.ecl ../ocaml-vm/vm/fail.ecl ../ocaml-vm/vm/ram.ecl ../ocaml-vm/vm/runtime.ecl ../ocaml-vm/vm/debug.ecl ../ocaml-vm/vm/alloc.ecl ../ocaml-vm/vm/prims.ecl ../ocaml-vm/bytecode.ecl ../ocaml-vm/vm/vm.ecl ../ocaml-vm/vm/target-specific/intel-max10/IOs.ecl ../ocaml-vm/vm/target-specific/intel-max10/main.ecl

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.runtime.all;


entity main is
  
  port(signal clk    : in std_logic;
       signal reset  : in std_logic;
       signal run    : in std_logic;
       signal rdy    : out value(0 to 0);
       signal argument : in value(0 to 11);
       signal result : out value(0 to 57));
       
end entity;
architecture rtl of main is

  type t_state is (compute5551);
  signal state: t_state;
  type t_state_var6680 is (compute6667);
  signal state_var6680: t_state_var6680;
  type t_state_var6679 is (compute5565, pause_setI5566, pause_setI5570, pause_setI5574, pause_setI5578, pause_setI5582, pause_setI5586, pause_setI5590, pause_setI5594, pause_setI5598, pause_setI5602, pause_setI5606, pause_setI5610, pause_setI5614, pause_setI5618, pause_setI5622, pause_setI5626, pause_setI5630, pause_setI5634, pause_setI5638, pause_setI5642, pause_setI5646, pause_setI5650, pause_setI5654, pause_setI5658, pause_setI5662, pause_setI5666, pause_setI5670, pause_setI5674, pause_setI5678, pause_setI5682, pause_setI5686, pause_setI5690, pause_setI5694, pause_setI5698, pause_setI5702, pause_setI5706, pause_setII5567, pause_setII5571, pause_setII5575, pause_setII5579, pause_setII5583, pause_setII5587, pause_setII5591, pause_setII5595, pause_setII5599, pause_setII5603, pause_setII5607, pause_setII5611, pause_setII5615, pause_setII5619, pause_setII5623, pause_setII5627, pause_setII5631, pause_setII5635, pause_setII5639, pause_setII5643, pause_setII5647, pause_setII5651, pause_setII5655, pause_setII5659, pause_setII5663, pause_setII5667, pause_setII5671, pause_setII5675, pause_setII5679, pause_setII5683, pause_setII5687, pause_setII5691, pause_setII5695, pause_setII5699, pause_setII5703, pause_setII5707, q_wait5568, q_wait5572, q_wait5576, q_wait5580, q_wait5584, q_wait5588, q_wait5592, q_wait5596, q_wait5600, q_wait5604, q_wait5608, q_wait5612, q_wait5616, q_wait5620, q_wait5624, q_wait5628, q_wait5632, q_wait5636, q_wait5640, q_wait5644, q_wait5648, q_wait5652, q_wait5656, q_wait5660, q_wait5664, q_wait5668, q_wait5672, q_wait5676, q_wait5680, q_wait5684, q_wait5688, q_wait5692, q_wait5696, q_wait5700, q_wait5704, q_wait5708);
  signal state_var6679: t_state_var6679;
  type t_state_var6678 is (compute5560);
  signal state_var6678: t_state_var6678;
  type t_state_var6677 is (compute5726, \$14343_copy_root_in_ram604\, \$14350_aux605\, \$14360_forever611\, \$14386_loop606\, \$14453_loop607\, \$14580_loop607\, \$14676_loop607\, \$14772_loop607\, pause_getI5735, pause_getI5752, pause_getI5757, pause_getI5762, pause_getI5775, pause_getI5792, pause_getI5797, pause_getI5802, pause_getI5807, pause_getI5813, pause_getI5821, pause_getI5838, pause_getI5843, pause_getI5852, pause_getI5869, pause_getI5874, pause_getII5736, pause_getII5753, pause_getII5758, pause_getII5763, pause_getII5776, pause_getII5793, pause_getII5798, pause_getII5803, pause_getII5808, pause_getII5814, pause_getII5822, pause_getII5839, pause_getII5844, pause_getII5853, pause_getII5870, pause_getII5875, pause_setI5727, pause_setI5731, pause_setI5740, pause_setI5744, pause_setI5748, pause_setI5767, pause_setI5771, pause_setI5780, pause_setI5784, pause_setI5788, pause_setI5817, pause_setI5826, pause_setI5830, pause_setI5834, pause_setI5848, pause_setI5857, pause_setI5861, pause_setI5865, pause_setII5728, pause_setII5732, pause_setII5741, pause_setII5745, pause_setII5749, pause_setII5768, pause_setII5772, pause_setII5781, pause_setII5785, pause_setII5789, pause_setII5818, pause_setII5827, pause_setII5831, pause_setII5835, pause_setII5849, pause_setII5858, pause_setII5862, pause_setII5866, q_wait5729, q_wait5733, q_wait5737, q_wait5742, q_wait5746, q_wait5750, q_wait5754, q_wait5759, q_wait5764, q_wait5769, q_wait5773, q_wait5777, q_wait5782, q_wait5786, q_wait5790, q_wait5794, q_wait5799, q_wait5804, q_wait5809, q_wait5815, q_wait5819, q_wait5823, q_wait5828, q_wait5832, q_wait5836, q_wait5840, q_wait5845, q_wait5850, q_wait5854, q_wait5859, q_wait5863, q_wait5867, q_wait5871, q_wait5876);
  signal state_var6677: t_state_var6677;
  type t_state_var6676 is (compute5723);
  signal state_var6676: t_state_var6676;
  type t_state_var6675 is (compute5716, \$12199_make_block525\, \$12235_apply579\, \$12236_offsetclosure_n580\, \$12237_binop_int584\, \$12238_compare585\, \$12239_binop_compare586\, \$12240_make_block_n587\, \$12241_branch_if589\, \$12245_compbranch590\, \$12265_w0591\, \$12267_w1592\, \$12270_w3593\, \$12421_w594\, \$12474_fill595\, \$12564_fill596\, \$12782_w597\, \$12909_forever611\, \$12946_forever611\, \$13261_forever611\, \$13539_loop_push598\, \$13928_forever611\, \$13935_forever611\, \$13942_forever611\, \$14090_modulo609\, \$14105_modulo609\, \$14274_wait603\, pause_getI5884, pause_getI5916, pause_getI5921, pause_getI5926, pause_getI5937, pause_getI5942, pause_getI5950, pause_getI5959, pause_getI5969, pause_getI5974, pause_getI5978, pause_getI5982, pause_getI5986, pause_getI5990, pause_getI5994, pause_getI5998, pause_getI6002, pause_getI6014, pause_getI6022, pause_getI6030, pause_getI6038, pause_getI6046, pause_getI6054, pause_getI6062, pause_getI6070, pause_getI6074, pause_getI6078, pause_getI6082, pause_getI6086, pause_getI6094, pause_getI6102, pause_getI6110, pause_getI6122, pause_getI6127, pause_getI6131, pause_getI6151, pause_getI6155, pause_getI6159, pause_getI6163, pause_getI6171, pause_getI6179, pause_getI6187, pause_getI6195, pause_getI6199, pause_getI6203, pause_getI6207, pause_getI6215, pause_getI6219, pause_getI6223, pause_getI6227, pause_getI6235, pause_getI6239, pause_getI6243, pause_getI6247, pause_getI6251, pause_getI6255, pause_getI6259, pause_getI6279, pause_getI6283, pause_getI6295, pause_getI6299, pause_getI6319, pause_getI6323, pause_getI6327, pause_getI6331, pause_getI6335, pause_getI6344, pause_getI6349, pause_getI6353, pause_getI6357, pause_getI6374, pause_getI6378, pause_getI6394, pause_getI6402, pause_getI6406, pause_getI6410, pause_getI6431, pause_getI6440, pause_getI6449, pause_getI6453, pause_getI6462, pause_getI6466, pause_getI6470, pause_getI6479, pause_getI6483, pause_getI6487, pause_getI6491, pause_getI6500, pause_getI6504, pause_getI6508, pause_getI6512, pause_getI6524, pause_getI6532, pause_getI6537, pause_getI6545, pause_getI6559, pause_getI6563, pause_getI6567, pause_getI6571, pause_getI6583, pause_getI6596, pause_getI6605, pause_getI6632, pause_getI6637, pause_getI6642, pause_getI6647, pause_getI6652, pause_getII5885, pause_getII5917, pause_getII5922, pause_getII5927, pause_getII5938, pause_getII5943, pause_getII5951, pause_getII5960, pause_getII5970, pause_getII5975, pause_getII5979, pause_getII5983, pause_getII5987, pause_getII5991, pause_getII5995, pause_getII5999, pause_getII6003, pause_getII6015, pause_getII6023, pause_getII6031, pause_getII6039, pause_getII6047, pause_getII6055, pause_getII6063, pause_getII6071, pause_getII6075, pause_getII6079, pause_getII6083, pause_getII6087, pause_getII6095, pause_getII6103, pause_getII6111, pause_getII6123, pause_getII6128, pause_getII6132, pause_getII6152, pause_getII6156, pause_getII6160, pause_getII6164, pause_getII6172, pause_getII6180, pause_getII6188, pause_getII6196, pause_getII6200, pause_getII6204, pause_getII6208, pause_getII6216, pause_getII6220, pause_getII6224, pause_getII6228, pause_getII6236, pause_getII6240, pause_getII6244, pause_getII6248, pause_getII6252, pause_getII6256, pause_getII6260, pause_getII6280, pause_getII6284, pause_getII6296, pause_getII6300, pause_getII6320, pause_getII6324, pause_getII6328, pause_getII6332, pause_getII6336, pause_getII6345, pause_getII6350, pause_getII6354, pause_getII6358, pause_getII6375, pause_getII6379, pause_getII6395, pause_getII6403, pause_getII6407, pause_getII6411, pause_getII6432, pause_getII6441, pause_getII6450, pause_getII6454, pause_getII6463, pause_getII6467, pause_getII6471, pause_getII6480, pause_getII6484, pause_getII6488, pause_getII6492, pause_getII6501, pause_getII6505, pause_getII6509, pause_getII6513, pause_getII6525, pause_getII6533, pause_getII6538, pause_getII6546, pause_getII6560, pause_getII6564, pause_getII6568, pause_getII6572, pause_getII6584, pause_getII6597, pause_getII6606, pause_getII6633, pause_getII6638, pause_getII6643, pause_getII6648, pause_getII6653, pause_setI5717, pause_setI5888, pause_setI5893, pause_setI5898, pause_setI5903, pause_setI5907, pause_setI5911, pause_setI5946, pause_setI5955, pause_setI5964, pause_setI6006, pause_setI6010, pause_setI6018, pause_setI6026, pause_setI6034, pause_setI6042, pause_setI6050, pause_setI6058, pause_setI6066, pause_setI6090, pause_setI6098, pause_setI6106, pause_setI6114, pause_setI6118, pause_setI6135, pause_setI6139, pause_setI6143, pause_setI6147, pause_setI6167, pause_setI6175, pause_setI6183, pause_setI6191, pause_setI6211, pause_setI6231, pause_setI6263, pause_setI6267, pause_setI6271, pause_setI6275, pause_setI6287, pause_setI6291, pause_setI6303, pause_setI6307, pause_setI6311, pause_setI6315, pause_setI6340, pause_setI6361, pause_setI6365, pause_setI6370, pause_setI6382, pause_setI6386, pause_setI6390, pause_setI6398, pause_setI6415, pause_setI6419, pause_setI6423, pause_setI6427, pause_setI6436, pause_setI6445, pause_setI6458, pause_setI6475, pause_setI6496, pause_setI6516, pause_setI6520, pause_setI6528, pause_setI6541, pause_setI6550, pause_setI6554, pause_setI6575, pause_setI6579, pause_setI6588, pause_setI6592, pause_setI6601, pause_setI6609, pause_setI6614, pause_setI6619, pause_setI6623, pause_setI6627, pause_setII5718, pause_setII5889, pause_setII5894, pause_setII5899, pause_setII5904, pause_setII5908, pause_setII5912, pause_setII5947, pause_setII5956, pause_setII5965, pause_setII6007, pause_setII6011, pause_setII6019, pause_setII6027, pause_setII6035, pause_setII6043, pause_setII6051, pause_setII6059, pause_setII6067, pause_setII6091, pause_setII6099, pause_setII6107, pause_setII6115, pause_setII6119, pause_setII6136, pause_setII6140, pause_setII6144, pause_setII6148, pause_setII6168, pause_setII6176, pause_setII6184, pause_setII6192, pause_setII6212, pause_setII6232, pause_setII6264, pause_setII6268, pause_setII6272, pause_setII6276, pause_setII6288, pause_setII6292, pause_setII6304, pause_setII6308, pause_setII6312, pause_setII6316, pause_setII6341, pause_setII6362, pause_setII6366, pause_setII6371, pause_setII6383, pause_setII6387, pause_setII6391, pause_setII6399, pause_setII6416, pause_setII6420, pause_setII6424, pause_setII6428, pause_setII6437, pause_setII6446, pause_setII6459, pause_setII6476, pause_setII6497, pause_setII6517, pause_setII6521, pause_setII6529, pause_setII6542, pause_setII6551, pause_setII6555, pause_setII6576, pause_setII6580, pause_setII6589, pause_setII6593, pause_setII6602, pause_setII6610, pause_setII6615, pause_setII6620, pause_setII6624, pause_setII6628, q_wait5719, q_wait5886, q_wait5890, q_wait5895, q_wait5900, q_wait5905, q_wait5909, q_wait5913, q_wait5918, q_wait5923, q_wait5928, q_wait5939, q_wait5944, q_wait5948, q_wait5952, q_wait5957, q_wait5961, q_wait5966, q_wait5971, q_wait5976, q_wait5980, q_wait5984, q_wait5988, q_wait5992, q_wait5996, q_wait6000, q_wait6004, q_wait6008, q_wait6012, q_wait6016, q_wait6020, q_wait6024, q_wait6028, q_wait6032, q_wait6036, q_wait6040, q_wait6044, q_wait6048, q_wait6052, q_wait6056, q_wait6060, q_wait6064, q_wait6068, q_wait6072, q_wait6076, q_wait6080, q_wait6084, q_wait6088, q_wait6092, q_wait6096, q_wait6100, q_wait6104, q_wait6108, q_wait6112, q_wait6116, q_wait6120, q_wait6124, q_wait6129, q_wait6133, q_wait6137, q_wait6141, q_wait6145, q_wait6149, q_wait6153, q_wait6157, q_wait6161, q_wait6165, q_wait6169, q_wait6173, q_wait6177, q_wait6181, q_wait6185, q_wait6189, q_wait6193, q_wait6197, q_wait6201, q_wait6205, q_wait6209, q_wait6213, q_wait6217, q_wait6221, q_wait6225, q_wait6229, q_wait6233, q_wait6237, q_wait6241, q_wait6245, q_wait6249, q_wait6253, q_wait6257, q_wait6261, q_wait6265, q_wait6269, q_wait6273, q_wait6277, q_wait6281, q_wait6285, q_wait6289, q_wait6293, q_wait6297, q_wait6301, q_wait6305, q_wait6309, q_wait6313, q_wait6317, q_wait6321, q_wait6325, q_wait6329, q_wait6333, q_wait6337, q_wait6342, q_wait6346, q_wait6351, q_wait6355, q_wait6359, q_wait6363, q_wait6367, q_wait6372, q_wait6376, q_wait6380, q_wait6384, q_wait6388, q_wait6392, q_wait6396, q_wait6400, q_wait6404, q_wait6408, q_wait6412, q_wait6417, q_wait6421, q_wait6425, q_wait6429, q_wait6433, q_wait6438, q_wait6442, q_wait6447, q_wait6451, q_wait6455, q_wait6460, q_wait6464, q_wait6468, q_wait6472, q_wait6477, q_wait6481, q_wait6485, q_wait6489, q_wait6493, q_wait6498, q_wait6502, q_wait6506, q_wait6510, q_wait6514, q_wait6518, q_wait6522, q_wait6526, q_wait6530, q_wait6534, q_wait6539, q_wait6543, q_wait6547, q_wait6552, q_wait6556, q_wait6561, q_wait6565, q_wait6569, q_wait6573, q_wait6577, q_wait6581, q_wait6585, q_wait6590, q_wait6594, q_wait6598, q_wait6603, q_wait6607, q_wait6611, q_wait6616, q_wait6621, q_wait6625, q_wait6629, q_wait6634, q_wait6639, q_wait6644, q_wait6649, q_wait6654);
  signal state_var6675: t_state_var6675;
  type t_state_var6674 is (compute5713);
  signal state_var6674: t_state_var6674;
  type t_state_var6673 is (compute5558);
  signal state_var6673: t_state_var6673;
  type t_state_var6672 is (compute5553);
  signal state_var6672: t_state_var6672;
  type t_state_var6671 is (compute5553);
  signal state_var6671: t_state_var6671;
  type array_value_16 is array (natural range <>) of value(0 to 15);
  type array_value_31 is array (natural range <>) of value(0 to 30);
  type array_value_32 is array (natural range <>) of value(0 to 31);
  signal ram : array_value_32(0 to 16383) := (others => "000"& X"000000" & X"0" & eclat_true);
  signal \$ram_value\ : value(0 to 31);
  signal \$ram_ptr\ : natural range 0 to 16383;
  signal \$ram_ptr_write\ : natural range 0 to 16383;
  signal \$ram_write\ : value(0 to 31);
  signal \$ram_write_request\ : std_logic := '0';
  signal global_end : array_value_16(0 to 0) := (others => X"000" & X"0");
  signal \$global_end_value\ : value(0 to 15);
  signal \$global_end_ptr\ : natural range 0 to 0;
  signal \$global_end_ptr_write\ : natural range 0 to 0;
  signal \$global_end_write\ : value(0 to 15);
  signal \$global_end_write_request\ : std_logic := '0';
  signal code : array_value_31(0 to 34) := (others => "000"& X"000000" & X"0");
  signal \$code_value\ : value(0 to 30);
  signal \$code_ptr\ : natural range 0 to 34;
  signal \$code_ptr_write\ : natural range 0 to 34;
  signal \$code_write\ : value(0 to 30);
  signal \$code_write_request\ : std_logic := '0';
  
  begin
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$ram_write_request\ = '1' then
                    ram(\$ram_ptr_write\) <= \$ram_write\;
                  else
                   \$ram_value\ <= ram(\$ram_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$global_end_write_request\ = '1' then
                    global_end(\$global_end_ptr_write\) <= \$global_end_write\;
                  else
                   \$global_end_value\ <= global_end(\$global_end_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$code_write_request\ = '1' then
                    code(\$code_ptr_write\) <= \$code_write\;
                  else
                   \$code_value\ <= code(\$code_ptr\);
                  end if;
            end if;
        end process;
    
    process(clk)
      variable \$14855\ : value(0 to 1) := (others => '0');
      variable \$12257\, \$13996\, \$14386_loop606_arg\, \$12556\, 
               \$12199_make_block525_result\, \$12770\, \$12265_w0591_arg\, 
               \$12466\ : value(0 to 95) := (others => '0');
      variable \$12238_compare585_arg\ : value(0 to 93) := (others => '0');
      variable \$14186\, \$14323\, \$14340\, \$14180\, \$14422\, \$14547\, 
               \$14183\ : value(0 to 47) := (others => '0');
      variable \$14453_loop607_arg\, \$14676_loop607_arg\, 
               \$13539_loop_push598_arg\, \$12421_w594_arg\, 
               \$12782_w597_arg\, \$14772_loop607_arg\, \$14580_loop607_arg\, 
               \$14350_aux605_arg\ : value(0 to 63) := (others => '0');
      variable \$v6651\, \$v6636\, \$v6646\, \$v6641\ : value(0 to 7) := (others => '0');
      variable \$12176\, \$12241_branch_if589_arg\, \$12196\, \$12190\ : value(0 to 122) := (others => '0');
      variable \$14002_sp\, \$13543_sp\, \$14346_next\, 
               \$13539_loop_push598_result\, \$14189_sp\, 
               \$12564_fill596_result\, \$14343_copy_root_in_ram604_result\, 
               \$14345\, \$14344_next\, \$12270_w3593_result\, \$14190_sp\, 
               \$14351_next\, \$14386_loop606_result\, \$12265_w0591_result\, 
               \$14191_sp\, \$12782_w597_result\, \$12266_sp\, \$12953_ofs\, 
               \$12475_sp\, \$14001_sp\, \$12271_sp\, 
               \$12474_fill595_result\, \$12565_sp\, \$12783_sp\, 
               \$14387_next\, \$14350_aux605_result\, \$12256_sp\, 
               \$14192_sp\, \$12465_sp\ : value(0 to 15) := (others => '0');
      variable \$14105_modulo609_arg\, \$14090_modulo609_arg\ : value(0 to 61) := (others => '0');
      variable \$14274_wait603_arg\ : value(0 to 96) := (others => '0');
      variable result5549 : value(0 to 57) := (others => '0');
      variable \$12245_compbranch590_arg\ : value(0 to 215) := (others => '0');
      variable \$12143\, \$12168\ : value(0 to 3) := (others => '0');
      variable \$12199_make_block525_id\, \$14343_copy_root_in_ram604_id\, 
               \$12238_compare585_id\ : value(0 to 11) := (others => '0');
      variable \$v6435\, \$14106_r\, \$12321\, \$12243\, \$12954\, \$12253\, 
               \$v6444\, \$14090_modulo609_result\, \$12248_argument2\, 
               \$v6474\, \$12250_argument3\, \$13972_arg\, \$14086_res\, 
               \$v6495\, \$14091_r\, \$14105_modulo609_result\, \$v6457\, 
               \$12246_argument1\ : value(0 to 30) := (others => '0');
      variable \$12236_offsetclosure_n580_arg\ : value(0 to 137) := (others => '0');
      variable result5724 : value(0 to 127) := (others => '0');
      variable \$12199_make_block525_arg\ : value(0 to 103) := (others => '0');
      variable \$v6503\, \$v6294\, \$v6443\, \$12238_compare585_result\, 
               \$v5896\, \$v5806\, \$v5837\, \$v5770\, \$v5919\, \$v6659\, 
               \$v5954\, \$v6618\, \$v5661\, \$v5981\, \$v6655\, \$v6523\, 
               \$v5585\, \$v6660\, \$v6574\, \$v6535\, \$v6461\, \$v5738\, 
               \$v6553\, \$v5685\, \$v6109\, \$v5811\, \$v6093\, \$v6302\, 
               rdy5559, \$v5810\, \$v5915\, \$v5856\, \$v5633\, \$v6254\, 
               \$v6613\, \$v5881\, \$14858_rdy\, \$v5872\, \$v6630\, 
               \$v6278\, \$v5569\, \$v5973\, \$v6507\, \$v5860\, \$v6426\, 
               \$14676_loop607_result\, \$v5653\, \$v6258\, \$v6635\, 
               \$v5962\, \$v6562\, \$v6166\, \$v5791\, \$v6612\, \$v6360\, 
               \$v6373\, \$v5621\, rdy5712, \$v5779\, \$v6226\, \$v6544\, 
               \$v6381\, \$v6401\, \$v6413\, \$v5629\, \$v6494\, \$v5669\, 
               \$v6604\, \$v6270\, \$v5720\, \$v5556\, \$v5883\, \$v5787\, 
               \$v5555\, \$v5774\, \$v6322\, \$v6029\, 
               \$14580_loop607_result\, \$v6266\, \$v6586\, \$v5914\, 
               \$v6045\, \$v6274\, \$v5864\, \$v5930\, \$v6456\, \$v6310\, 
               rdy5552, \$v6125\, \$v6326\, \$v6210\, \$v5577\, \$v6101\, 
               \$v6113\, \$v6389\, \$v6665\, \$v6069\, \$v6202\, \$v6465\, 
               \$v6527\, \$v6049\, \$v5711\, \$v6558\, result5563, \$v6511\, 
               \$v6397\, \$v6222\, \$v6540\, \$v6041\, \$v5689\, \$v6097\, 
               \$v6452\, \$v6154\, \$v6548\, \$v6536\, \$v6001\, \$v5902\, 
               \$v5958\, \$v6670\, \$v5673\, \$v5910\, \$v5816\, \$v5842\, 
               \$v6025\, \$v5681\, \$v5625\, \$v5709\, \$v5901\, \$v6150\, 
               \$v5677\, \$v5877\, \$v6282\, \$v6081\, \$v6186\, \$v6531\, 
               \$v5657\, \$v5997\, \$v5609\, rdy5564, \$v6121\, \$v6298\, 
               \$v5925\, \$v6650\, rdy5550, \$v5641\, \$v5783\, \$v6142\, 
               \$v6138\, \$v6061\, \$v6242\, \$v6515\, \$v5963\, \$v5879\, 
               \$v6037\, \$v5665\, \$v5739\, \$v5873\, \$v6393\, \$v5993\, 
               \$v6238\, \$v5613\, rdy5725, \$v6622\, \$v6656\, \$v6591\, 
               \$v6486\, \$v5972\, \$v6414\, \$v5934\, \$v6057\, \$v6669\, 
               \$v5637\, \$v6250\, \$v6418\, \$v6218\, \$v6478\, \$v6347\, 
               \$v6198\, \$v6338\, \$v6640\, \$v5800\, \$v6339\, \$v5968\, 
               \$v5581\, \$v6409\, \$v6089\, \$v6631\, \$v5747\, \$v5605\, 
               \$v5891\, \$v5940\, \$v6599\, \$v6318\, \$v6430\, \$v6286\, 
               \$v5906\, \$14052_res\, \$v5924\, \$v6021\, rdy5722, \$v6578\, 
               \$v5929\, \$v5765\, \$v5833\, \$v5820\, \$v6519\, \$v5649\, 
               \$v5920\, \$v6234\, \$v6170\, \$v6146\, \$v6073\, \$v5597\, 
               \$v6230\, \$v6005\, \$v6013\, \$14453_loop607_result\, 
               \$v5949\, \$v6469\, \$v6162\, \$v5743\, \$v5766\, \$v6595\, 
               \$v6009\, \$v6663\, \$12421_w594_result\, \$v6617\, \$v5887\, 
               \$14772_loop607_result\, \$v6314\, \$v5693\, \$v5931\, 
               \$v6626\, \$v5801\, \$v5730\, \$v5760\, \$v5878\, \$v5935\, 
               \$v5705\, \$v5721\, \$v6364\, \$v5977\, \$v6085\, \$v6065\, 
               \$v5805\, \$v6566\, \$v5697\, \$v5847\, \$v5855\, \$v6343\, 
               \$v6182\, \$v6549\, \$v6645\, \$v5589\, \$v5933\, \$v5967\, 
               rdy6666, \$v5645\, \$v6290\, \$v6053\, \$v6369\, \$v5892\, 
               \$v5945\, \$v6306\, \$v6017\, \$v5573\, \$v6405\, \$v5593\, 
               \$v6482\, \$v6330\, \$v6439\, \$v5778\, \$v6194\, \$v5751\, 
               \$v5761\, \$v5824\, \$v6178\, \$v6385\, \$v6190\, \$v5601\, 
               \$v5841\, \$v5734\, \$v6348\, \$v5989\, \$v6662\, \$v5868\, 
               \$12267_w1592_result\, \$v6587\, \$v5825\, \$v6158\, \$v6105\, 
               rdy5715, \$v6077\, \$v5701\, \$v5953\, \$v6448\, \$v6206\, 
               \$v6352\, \$v6422\, \$v6262\, \$v6334\, rdy5557, \$v5829\, 
               \$v5851\, \$v6368\, \$v6126\, \$v6657\, \$v6214\, \$v6356\, 
               \$v6117\, \$v5932\, \$v5756\, \$v6174\, \$v6246\, \$v5795\, 
               \$v6473\, \$v6600\, \$v6582\, \$v5985\, \$v6434\, \$v5755\, 
               \$v5617\, \$v6377\, \$v5562\, \$v5796\, \$v6033\, \$14859\, 
               \$13322_b\, \$v5846\, \$v6490\, \$v6130\, \$v6134\, \$v6608\, 
               \$v5812\, \$v6499\, \$v6570\, \$v6557\, \$v5897\ : value(0 to 0) := (others => '0');
      variable \$12240_make_block_n587_arg\ : value(0 to 171) := (others => '0');
      variable \$12474_fill595_arg\, \$14274_wait603_result\, 
               \$12270_w3593_arg\, \$14250\, \$12267_w1592_arg\, \$14329\, 
               \$12564_fill596_arg\, \$14343_copy_root_in_ram604_arg\ : value(0 to 79) := (others => '0');
      variable \$12235_apply579_arg\ : value(0 to 165) := (others => '0');
      variable \$14302\, \$14292\ : value(0 to 128) := (others => '0');
      variable \$13192\, \$12239_binop_compare586_arg\, \$13134\, \$13023\, 
               \$13052\, \$12237_binop_int584_arg\, \$13088\ : value(0 to 153) := (others => '0');
      variable \$12709_v\, \$12426\, \$13413_v\, \$12920_v\, \$13869_v\, 
               \$13873_v\, \$12634\, \$14434_w\, \$13676_v\, \$14543\, 
               \$13358_v\, \$13774_v\, \$13725_v\, \$13333_v\, \$13475\, 
               \$14196\, \$12455\, \$12713_v\, \$12784_v\, \$12648\, 
               \$14907\, \$12878_v\, \$13691_v\, \$13854_v\, \$13538_hd\, 
               \$13487\, \$13338_v\, \$12528_v\, \$12376_v\, \$12820_v\, 
               \$12683\, \$13348_v\, \$14418\, \$14487\, \$13431_v\, 
               \$14758_hd\, \$13646_v\, \$v5936\, \$12965_hd\, \$13353_v\, 
               \$13878_v\, \$13877_v\, \$14082_v\, \$12580_v\, \$13712_v\, 
               \$12142_cy\, \$12544_v\, \$13377_v\, \$14439_hd\, \$13464\, 
               \$12490_v\, \$12788_v\, \$13661_v\, \$13754_hd\, \$13825_v\, 
               \$13824_v\, \$14382\, \$13422_v\, \$12789_v\, \$13785_v\, 
               \$12754\, \$13767_v\, \$12540\, \$14753_w\, \$13699_v\, 
               \$13363_v\, \$14662_hd\, \$14657_w\, \$14230_v\, \$12604_v\, 
               \$13442\, \$14614\, \$13807_v\, \$12160\, \$12524\, \$13453\, 
               \$12612_v\, \$13500\, \$14710\, \$14227_v\, \$13395_v\, 
               \$13146_v\, \$12872_v\, \$14561_w\, \$13035_v\, \$13784_v\, 
               \$13328_v\, \$13386_v\, \$13589\, \$v5941\, \$13814_next_acc\, 
               \$12149\, \$12714_v\, \$14014_v\, \$13343_v\, \$14233_v\, 
               \$13100_v\, \$14048_v\, \$13404_v\, \$13526\, \$13204_v\, 
               \$13738_v\, \$14566_hd\, \$14003_v\, \$13278_f0\, 
               \$13547_next_env\, \$12929_v\, \$13513\, \$14806\, \$13064_v\ : value(0 to 31) := (others => '0');
      variable \$12240_make_block_n587_result\, result5714, 
               \$12235_apply579_result\, \$12245_compbranch590_result\, 
               \$12241_branch_if589_result\, \$12237_binop_int584_result\, 
               \$12236_offsetclosure_n580_result\, 
               \$12239_binop_compare586_result\ : value(0 to 121) := (others => '0');
      variable \$ram_ptr_take\ : value(0 to 0) := "0";
      variable \$global_end_ptr_take\ : value(0 to 0) := "0";
      variable \$code_ptr_take\ : value(0 to 0) := "0";
      
    begin
      
      if rising_edge(clk) then
        if (reset = '1') then
          default_zero(\$14350_aux605_arg\); default_zero(\$v5897\); 
          default_zero(\$v6557\); default_zero(\$v6570\); 
          default_zero(\$v6499\); default_zero(\$v5812\); 
          default_zero(\$v6608\); default_zero(\$13064_v\); 
          default_zero(\$v6134\); default_zero(\$14806\); 
          default_zero(\$13513\); default_zero(\$v6130\); 
          default_zero(\$14183\); default_zero(\$14090_modulo609_arg\); 
          default_zero(\$12246_argument1\); 
          default_zero(\$12235_apply579_arg\); default_zero(\$v6457\); 
          default_zero(\$v6490\); default_zero(\$14580_loop607_arg\); 
          default_zero(\$v5846\); default_zero(\$13322_b\); 
          default_zero(\$12465_sp\); default_zero(\$14859\); 
          default_zero(\$v6033\); default_zero(\$12929_v\); 
          default_zero(\$13088\); default_zero(\$v5796\); 
          default_zero(\$v5562\); default_zero(\$v6377\); 
          default_zero(\$v5617\); default_zero(\$13547_next_env\); 
          default_zero(\$v5755\); default_zero(\$v6434\); 
          default_zero(\$13278_f0\); default_zero(\$14003_v\); 
          default_zero(\$14547\); default_zero(\$14566_hd\); 
          default_zero(\$v5985\); default_zero(\$v6582\); 
          default_zero(\$13738_v\); default_zero(\$14422\); 
          default_zero(\$v6600\); default_zero(\$v6473\); 
          default_zero(\$v5795\); 
          default_zero(\$12239_binop_compare586_result\); 
          default_zero(\$v6246\); default_zero(\$v6174\); 
          default_zero(\$14192_sp\); default_zero(\$14292\); 
          default_zero(\$14105_modulo609_result\); default_zero(\$v5756\); 
          default_zero(\$v5932\); default_zero(\$v6117\); 
          default_zero(\$v6356\); default_zero(\$12256_sp\); 
          default_zero(\$v6214\); default_zero(\$14772_loop607_arg\); 
          default_zero(\$v6657\); default_zero(\$v6126\); 
          default_zero(\$v6368\); default_zero(\$v5851\); 
          default_zero(\$v5829\); 
          default_zero(\$12236_offsetclosure_n580_result\); 
          default_zero(rdy5557); 
          default_zero(\$14343_copy_root_in_ram604_arg\); 
          default_zero(\$14274_wait603_arg\); default_zero(\$13204_v\); 
          default_zero(\$13526\); default_zero(\$v6334\); 
          default_zero(\$13404_v\); default_zero(\$v6262\); 
          default_zero(\$14048_v\); default_zero(\$v6422\); 
          default_zero(\$v6352\); default_zero(\$13100_v\); 
          default_zero(\$v6206\); default_zero(\$12564_fill596_arg\); 
          default_zero(\$v6448\); default_zero(\$14350_aux605_result\); 
          default_zero(\$v5953\); default_zero(\$v5701\); 
          default_zero(\$14329\); default_zero(\$v6077\); 
          default_zero(rdy5715); default_zero(\$v6105\); 
          default_zero(\$v6158\); default_zero(\$14233_v\); 
          default_zero(\$14180\); default_zero(\$12190\); 
          default_zero(\$v5825\); default_zero(\$v6587\); 
          default_zero(\$13343_v\); default_zero(\$14091_r\); 
          default_zero(\$12267_w1592_result\); default_zero(\$v5868\); 
          default_zero(\$v6662\); default_zero(\$v5989\); 
          default_zero(\$v6348\); default_zero(\$14014_v\); 
          default_zero(\$v5734\); default_zero(\$v5841\); 
          default_zero(\$v5601\); default_zero(\$12714_v\); 
          default_zero(\$v6190\); default_zero(\$v6385\); 
          default_zero(\$v6178\); default_zero(\$v5824\); 
          default_zero(\$12149\); default_zero(\$v5761\); 
          default_zero(\$v5751\); default_zero(\$12466\); 
          default_zero(\$12240_make_block_n587_arg\); default_zero(\$v6194\); 
          default_zero(\$v5778\); default_zero(\$v6439\); 
          default_zero(\$13814_next_acc\); default_zero(\$v5941\); 
          default_zero(\$12267_w1592_arg\); default_zero(\$13589\); 
          default_zero(\$13386_v\); default_zero(\$v6330\); 
          default_zero(\$13328_v\); default_zero(\$14387_next\); 
          default_zero(\$13784_v\); default_zero(\$12783_sp\); 
          default_zero(\$v6482\); default_zero(\$v5593\); 
          default_zero(\$13035_v\); default_zero(\$14561_w\); 
          default_zero(\$12872_v\); default_zero(\$v6405\); 
          default_zero(\$v5573\); default_zero(\$12237_binop_int584_result\); 
          default_zero(\$v6017\); default_zero(\$v6306\); 
          default_zero(\$v5945\); default_zero(\$v5892\); 
          default_zero(\$v6369\); default_zero(\$13146_v\); 
          default_zero(\$v6053\); default_zero(\$v6495\); 
          default_zero(\$v6290\); default_zero(\$13395_v\); 
          default_zero(\$14086_res\); 
          default_zero(\$12236_offsetclosure_n580_arg\); 
          default_zero(\$v5645\); default_zero(\$14227_v\); 
          default_zero(rdy6666); default_zero(\$v5967\); 
          default_zero(\$14250\); default_zero(\$14710\); 
          default_zero(\$13500\); default_zero(\$12238_compare585_id\); 
          default_zero(\$12612_v\); default_zero(\$v5933\); 
          default_zero(\$v5589\); default_zero(\$v6645\); 
          default_zero(\$14855\); default_zero(\$v6549\); 
          default_zero(\$v6182\); default_zero(\$12782_w597_arg\); 
          default_zero(\$v6343\); default_zero(\$v5855\); 
          default_zero(\$v5847\); default_zero(\$v5697\); 
          default_zero(\$v6566\); default_zero(\$v5805\); 
          default_zero(\$13453\); default_zero(\$v6065\); 
          default_zero(\$v6085\); default_zero(\$v5977\); 
          default_zero(\$12565_sp\); default_zero(\$12524\); 
          default_zero(\$13972_arg\); default_zero(\$12160\); 
          default_zero(\$v6364\); default_zero(\$12421_w594_arg\); 
          default_zero(\$v5721\); default_zero(\$v5705\); 
          default_zero(\$13807_v\); default_zero(\$v5935\); 
          default_zero(\$v5878\); default_zero(\$v5760\); 
          default_zero(\$v5730\); default_zero(\$v5801\); 
          default_zero(\$v6626\); default_zero(\$v5931\); 
          default_zero(\$14614\); default_zero(\$v5693\); 
          default_zero(\$v6314\); default_zero(\$13442\); 
          default_zero(\$14772_loop607_result\); default_zero(\$v5887\); 
          default_zero(\$v6617\); default_zero(\$12421_w594_result\); 
          default_zero(\$12250_argument3\); default_zero(\$v6663\); 
          default_zero(\$v6009\); default_zero(\$v6595\); 
          default_zero(\$v5766\); default_zero(\$v5743\); 
          default_zero(\$12237_binop_int584_arg\); default_zero(\$v6162\); 
          default_zero(\$v6469\); default_zero(\$v5949\); 
          default_zero(\$14453_loop607_result\); default_zero(\$v6013\); 
          default_zero(\$v6005\); default_zero(\$12474_fill595_result\); 
          default_zero(\$v6474\); default_zero(\$12196\); 
          default_zero(\$v6230\); default_zero(\$v5597\); 
          default_zero(\$v6073\); default_zero(\$v6146\); 
          default_zero(\$v6170\); default_zero(\$12604_v\); 
          default_zero(\$v6234\); default_zero(\$v5920\); 
          default_zero(\$v5649\); default_zero(\$v6519\); 
          default_zero(\$v5820\); default_zero(\$v5833\); 
          default_zero(\$v5765\); default_zero(\$12271_sp\); 
          default_zero(\$v5929\); default_zero(\$v6578\); 
          default_zero(rdy5722); default_zero(\$12270_w3593_arg\); 
          default_zero(\$14230_v\); default_zero(\$14657_w\); 
          default_zero(\$v6021\); default_zero(\$14662_hd\); 
          default_zero(\$13363_v\); default_zero(\$v5924\); 
          default_zero(\$14052_res\); default_zero(\$v5906\); 
          default_zero(\$14001_sp\); default_zero(\$13699_v\); 
          default_zero(\$14302\); default_zero(\$12241_branch_if589_result\); 
          default_zero(\$14753_w\); default_zero(\$v6286\); 
          default_zero(\$v6430\); default_zero(\$v6318\); 
          default_zero(\$v6599\); default_zero(\$12265_w0591_arg\); 
          default_zero(\$v5940\); default_zero(\$12199_make_block525_arg\); 
          default_zero(\$v5891\); default_zero(\$v5605\); 
          default_zero(\$v5747\); default_zero(\$v6631\); 
          default_zero(\$v6089\); default_zero(\$12540\); 
          default_zero(\$13767_v\); 
          default_zero(\$12245_compbranch590_result\); 
          default_zero(\$v6409\); default_zero(\$12754\); 
          default_zero(result5724); default_zero(\$v5581\); 
          default_zero(\$v5968\); default_zero(\$v6339\); 
          default_zero(\$13785_v\); default_zero(\$12789_v\); 
          default_zero(\$v5800\); default_zero(\$v6640\); 
          default_zero(\$13539_loop_push598_arg\); default_zero(\$12475_sp\); 
          default_zero(\$v6338\); default_zero(\$v6198\); 
          default_zero(\$v6347\); default_zero(\$v6478\); 
          default_zero(\$v6218\); default_zero(\$13422_v\); 
          default_zero(\$v6418\); default_zero(\$v6250\); 
          default_zero(\$v5637\); default_zero(\$v6669\); 
          default_zero(\$v6057\); default_zero(\$14382\); 
          default_zero(\$v5934\); default_zero(\$v6414\); 
          default_zero(\$13824_v\); default_zero(\$12770\); 
          default_zero(\$12235_apply579_result\); default_zero(\$13825_v\); 
          default_zero(\$v5972\); default_zero(\$v6486\); 
          default_zero(\$13754_hd\); default_zero(\$12238_compare585_arg\); 
          default_zero(\$v6591\); default_zero(\$v6656\); 
          default_zero(\$v6622\); default_zero(\$13661_v\); 
          default_zero(rdy5725); default_zero(\$14676_loop607_arg\); 
          default_zero(\$v5613\); default_zero(\$v6238\); 
          default_zero(\$v5993\); default_zero(\$v6393\); 
          default_zero(\$12788_v\); default_zero(\$12490_v\); 
          default_zero(\$v5873\); default_zero(\$v5739\); 
          default_zero(\$v5665\); default_zero(\$v6037\); 
          default_zero(\$12953_ofs\); default_zero(\$13464\); 
          default_zero(\$v5879\); default_zero(\$v5963\); 
          default_zero(\$v6515\); default_zero(\$v6242\); 
          default_zero(\$14439_hd\); default_zero(\$12266_sp\); 
          default_zero(result5714); default_zero(\$v6061\); 
          default_zero(\$v6138\); default_zero(\$v6142\); 
          default_zero(\$13377_v\); default_zero(\$v5783\); 
          default_zero(\$v5641\); default_zero(rdy5550); 
          default_zero(\$13052\); default_zero(\$v6650\); 
          default_zero(\$v5925\); default_zero(\$v6298\); 
          default_zero(\$v6121\); default_zero(rdy5564); 
          default_zero(\$v5609\); default_zero(\$v5997\); 
          default_zero(\$12248_argument2\); default_zero(\$v5657\); 
          default_zero(\$12544_v\); default_zero(\$v6531\); 
          default_zero(\$v6186\); default_zero(\$v6081\); 
          default_zero(\$v6282\); default_zero(\$v5877\); 
          default_zero(\$v5677\); default_zero(\$v6150\); 
          default_zero(\$12782_w597_result\); default_zero(\$v5901\); 
          default_zero(\$v5709\); default_zero(\$12142_cy\); 
          default_zero(\$12199_make_block525_result\); 
          default_zero(\$v5625\); default_zero(\$v5681\); 
          default_zero(\$v6025\); default_zero(\$v5842\); 
          default_zero(\$13712_v\); default_zero(\$12168\); 
          default_zero(\$v5816\); default_zero(\$v5910\); 
          default_zero(\$v5673\); default_zero(\$v6670\); 
          default_zero(\$12580_v\); default_zero(\$v5958\); 
          default_zero(\$v5902\); default_zero(\$v6001\); 
          default_zero(\$v6536\); default_zero(\$v6548\); 
          default_zero(\$v6154\); default_zero(\$v6452\); 
          default_zero(\$14082_v\); default_zero(\$13877_v\); 
          default_zero(\$v6097\); default_zero(\$v5689\); 
          default_zero(\$v6041\); 
          default_zero(\$12240_make_block_n587_result\); 
          default_zero(\$13878_v\); default_zero(\$v6540\); 
          default_zero(\$14191_sp\); default_zero(\$v6222\); 
          default_zero(\$13353_v\); default_zero(\$v6397\); 
          default_zero(\$14340\); default_zero(\$12965_hd\); 
          default_zero(\$12265_w0591_result\); default_zero(\$v5936\); 
          default_zero(\$v6511\); default_zero(\$13646_v\); 
          default_zero(\$14758_hd\); default_zero(result5563); 
          default_zero(\$13023\); default_zero(\$13431_v\); 
          default_zero(\$14090_modulo609_result\); default_zero(\$14487\); 
          default_zero(\$14418\); default_zero(\$v6558\); 
          default_zero(\$v5711\); default_zero(\$v6049\); 
          default_zero(\$v6527\); default_zero(\$v6465\); 
          default_zero(\$v6444\); default_zero(\$14105_modulo609_arg\); 
          default_zero(\$v6202\); default_zero(\$v6069\); 
          default_zero(\$14386_loop606_result\); default_zero(\$v6665\); 
          default_zero(\$v6389\); default_zero(\$13348_v\); 
          default_zero(\$v6113\); default_zero(\$v6101\); 
          default_zero(\$12683\); default_zero(\$12820_v\); 
          default_zero(\$v5577\); default_zero(\$v6210\); 
          default_zero(\$v6326\); default_zero(\$v6125\); 
          default_zero(\$14351_next\); default_zero(rdy5552); 
          default_zero(\$v6310\); default_zero(\$v6456\); 
          default_zero(\$14323\); default_zero(\$v5930\); 
          default_zero(\$12376_v\); default_zero(\$v5864\); 
          default_zero(\$v6274\); default_zero(\$v6045\); 
          default_zero(\$12528_v\); default_zero(\$v5914\); 
          default_zero(\$v6586\); default_zero(\$v6266\); 
          default_zero(\$v6641\); default_zero(\$14580_loop607_result\); 
          default_zero(\$14190_sp\); default_zero(\$13338_v\); 
          default_zero(\$v6029\); default_zero(\$v6322\); 
          default_zero(\$v5774\); default_zero(\$13487\); 
          default_zero(\$12270_w3593_result\); default_zero(\$13538_hd\); 
          default_zero(\$v5555\); default_zero(\$v5787\); 
          default_zero(\$v5883\); default_zero(\$v5556\); 
          default_zero(\$v5720\); default_zero(\$14344_next\); 
          default_zero(\$v6270\); default_zero(\$13854_v\); 
          default_zero(\$14345\); default_zero(\$v6604\); 
          default_zero(\$14274_wait603_result\); default_zero(\$12253\); 
          default_zero(\$v5669\); default_zero(\$12241_branch_if589_arg\); 
          default_zero(\$v6494\); default_zero(\$v5629\); 
          default_zero(\$v6413\); default_zero(\$v6401\); 
          default_zero(\$v6381\); default_zero(\$v6544\); 
          default_zero(\$13691_v\); default_zero(\$12878_v\); 
          default_zero(\$v6226\); default_zero(\$v5779\); 
          default_zero(\$14907\); default_zero(\$12556\); 
          default_zero(\$14343_copy_root_in_ram604_id\); 
          default_zero(rdy5712); default_zero(\$12648\); 
          default_zero(\$v5621\); default_zero(\$12474_fill595_arg\); 
          default_zero(\$12199_make_block525_id\); default_zero(\$v6373\); 
          default_zero(\$v6360\); default_zero(\$v6612\); 
          default_zero(\$12784_v\); default_zero(\$v5791\); 
          default_zero(\$12713_v\); default_zero(\$14386_loop606_arg\); 
          default_zero(\$v6646\); 
          default_zero(\$14343_copy_root_in_ram604_result\); 
          default_zero(\$v6166\); default_zero(\$v6562\); 
          default_zero(\$12564_fill596_result\); default_zero(\$12954\); 
          default_zero(\$v5962\); default_zero(\$v6635\); 
          default_zero(\$v6258\); default_zero(\$v5653\); 
          default_zero(\$14676_loop607_result\); default_zero(\$v6426\); 
          default_zero(\$v5860\); default_zero(\$12455\); 
          default_zero(\$v6507\); default_zero(\$v5973\); 
          default_zero(\$14196\); default_zero(\$v5569\); 
          default_zero(\$13996\); default_zero(\$v6278\); 
          default_zero(\$14189_sp\); 
          default_zero(\$12245_compbranch590_arg\); default_zero(\$v6630\); 
          default_zero(\$v5872\); default_zero(\$14453_loop607_arg\); 
          default_zero(\$14858_rdy\); default_zero(\$v5881\); 
          default_zero(\$v6613\); default_zero(\$12257\); 
          default_zero(\$v6254\); default_zero(\$13539_loop_push598_result\); 
          default_zero(\$v5633\); default_zero(\$13475\); 
          default_zero(\$v5856\); default_zero(\$13333_v\); 
          default_zero(\$v6636\); default_zero(\$13725_v\); 
          default_zero(\$v5915\); default_zero(\$v5810\); 
          default_zero(\$13774_v\); default_zero(rdy5559); 
          default_zero(\$v6302\); default_zero(\$v6093\); 
          default_zero(\$13358_v\); default_zero(\$14543\); 
          default_zero(\$12243\); default_zero(\$v5811\); 
          default_zero(\$12176\); default_zero(\$v6109\); 
          default_zero(\$v5685\); default_zero(\$v6553\); 
          default_zero(\$v5738\); default_zero(\$v6461\); 
          default_zero(\$13676_v\); default_zero(\$v6535\); 
          default_zero(\$14186\); default_zero(\$v6574\); 
          default_zero(\$14434_w\); default_zero(\$v6660\); 
          default_zero(\$v5585\); default_zero(\$v6651\); 
          default_zero(\$v6523\); default_zero(\$v6655\); 
          default_zero(result5549); default_zero(\$v5981\); 
          default_zero(\$v5661\); default_zero(\$13134\); 
          default_zero(\$12634\); default_zero(\$14346_next\); 
          default_zero(\$12143\); default_zero(\$v6618\); 
          default_zero(\$12239_binop_compare586_arg\); 
          default_zero(\$v5954\); default_zero(\$v6659\); 
          default_zero(\$13873_v\); default_zero(\$12321\); 
          default_zero(\$v5919\); default_zero(\$13869_v\); 
          default_zero(\$13543_sp\); default_zero(\$12920_v\); 
          default_zero(\$14106_r\); default_zero(\$13192\); 
          default_zero(\$13413_v\); default_zero(\$v5770\); 
          default_zero(\$v5837\); default_zero(\$v5806\); 
          default_zero(\$v5896\); default_zero(\$12426\); 
          default_zero(\$12709_v\); default_zero(\$v6435\); 
          default_zero(\$12238_compare585_result\); default_zero(\$v6443\); 
          default_zero(\$14002_sp\); default_zero(\$v6294\); 
          default_zero(\$v6503\); 
          rdy <= "1";
          rdy5550 := "0";
          state <= compute5551;
          state_var6680 <= compute6667;
          state_var6679 <= compute5565;
          state_var6678 <= compute5560;
          state_var6677 <= compute5726;
          state_var6676 <= compute5723;
          state_var6675 <= compute5716;
          state_var6674 <= compute5713;
          state_var6673 <= compute5558;
          state_var6672 <= compute5553;
          state_var6671 <= compute5553;
          
        else if run = '1' then
          case state is
          when compute5551 =>
            rdy5550 := eclat_false;
            \$v6670\ := eclat_not(""&argument(10));
            if \$v6670\(0) = '1' then
              result5549 := ""&argument(11) & ""&argument(11) & ""&argument(11) & ""&argument(11) & ""&argument(11) & ""&argument(11) & ""&argument(11) & ""&argument(11) & ""&argument(11) & ""&argument(11) & "01100011" & "00000011" & "01110001" & "01110001" & "01100001" & "01100001";
              rdy5550 := eclat_true;
              state <= compute5551;
            else
              \$v6669\ := eclat_not(rdy6666);
              if \$v6669\(0) = '1' then
                \$14907\ := X"0000000" & X"0";
              end if;
              case state_var6680 is
              when compute6667 =>
                rdy6666 := eclat_false;
                \$14907\ := eclat_if(""&argument(11) & X"0000000" & X"0" & eclat_add(\$14907\ & X"0000000" & X"1"));
                rdy6666 := eclat_true;
                state_var6680 <= compute6667;
              end case;
              \$14907\ := \$14907\;
              \$12142_cy\ := \$14907\;
              \$v6665\ := eclat_not(rdy5557);
              if \$v6665\(0) = '1' then
                \$12168\ := eclat_false & eclat_false & eclat_false & eclat_false;
              end if;
              case state_var6673 is
              when compute5558 =>
                rdy5557 := eclat_false;
                \$v6663\ := eclat_not(""&\$12168\(2));
                if \$v6663\(0) = '1' then
                  case state_var6679 is
                  when pause_setI5566 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5567;
                  when pause_setI5570 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5571;
                  when pause_setI5574 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5575;
                  when pause_setI5578 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5579;
                  when pause_setI5582 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5583;
                  when pause_setI5586 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5587;
                  when pause_setI5590 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5591;
                  when pause_setI5594 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5595;
                  when pause_setI5598 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5599;
                  when pause_setI5602 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5603;
                  when pause_setI5606 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5607;
                  when pause_setI5610 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5611;
                  when pause_setI5614 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5615;
                  when pause_setI5618 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5619;
                  when pause_setI5622 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5623;
                  when pause_setI5626 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5627;
                  when pause_setI5630 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5631;
                  when pause_setI5634 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5635;
                  when pause_setI5638 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5639;
                  when pause_setI5642 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5643;
                  when pause_setI5646 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5647;
                  when pause_setI5650 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5651;
                  when pause_setI5654 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5655;
                  when pause_setI5658 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5659;
                  when pause_setI5662 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5663;
                  when pause_setI5666 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5667;
                  when pause_setI5670 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5671;
                  when pause_setI5674 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5675;
                  when pause_setI5678 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5679;
                  when pause_setI5682 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5683;
                  when pause_setI5686 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5687;
                  when pause_setI5690 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5691;
                  when pause_setI5694 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5695;
                  when pause_setI5698 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5699;
                  when pause_setI5702 =>
                    \$code_write_request\ <= '0';
                    state_var6679 <= pause_setII5703;
                  when pause_setI5706 =>
                    \$global_end_write_request\ <= '0';
                    state_var6679 <= pause_setII5707;
                  when pause_setII5567 =>
                    \$code_ptr_take\(0) := '0';
                    result5563 := eclat_unit;
                    rdy5564 := eclat_true;
                    state_var6679 <= compute5565;
                  when pause_setII5571 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5569\ := \$code_ptr_take\;
                    if \$v5569\(0) = '1' then
                      state_var6679 <= q_wait5568;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 34;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"8f";
                      state_var6679 <= pause_setI5566;
                    end if;
                  when pause_setII5575 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5573\ := \$code_ptr_take\;
                    if \$v5573\(0) = '1' then
                      state_var6679 <= q_wait5572;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 33;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"000000" & X"1";
                      state_var6679 <= pause_setI5570;
                    end if;
                  when pause_setII5579 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5577\ := \$code_ptr_take\;
                    if \$v5577\(0) = '1' then
                      state_var6679 <= q_wait5576;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 32;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"13";
                      state_var6679 <= pause_setI5574;
                    end if;
                  when pause_setII5583 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5581\ := \$code_ptr_take\;
                    if \$v5581\(0) = '1' then
                      state_var6679 <= q_wait5580;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 31;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"000000" & X"0";
                      state_var6679 <= pause_setI5578;
                    end if;
                  when pause_setII5587 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5585\ := \$code_ptr_take\;
                    if \$v5585\(0) = '1' then
                      state_var6679 <= q_wait5584;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 30;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"5d";
                      state_var6679 <= pause_setI5582;
                    end if;
                  when pause_setII5591 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5589\ := \$code_ptr_take\;
                    if \$v5589\(0) = '1' then
                      state_var6679 <= q_wait5588;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 29;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"21";
                      state_var6679 <= pause_setI5586;
                    end if;
                  when pause_setII5595 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5593\ := \$code_ptr_take\;
                    if \$v5593\(0) = '1' then
                      state_var6679 <= q_wait5592;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 28;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"000000" & X"b";
                      state_var6679 <= pause_setI5590;
                    end if;
                  when pause_setII5599 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5597\ := \$code_ptr_take\;
                    if \$v5597\(0) = '1' then
                      state_var6679 <= q_wait5596;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 27;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"000000" & X"b";
                      state_var6679 <= pause_setI5594;
                    end if;
                  when pause_setII5603 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5601\ := \$code_ptr_take\;
                    if \$v5601\(0) = '1' then
                      state_var6679 <= q_wait5600;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 26;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"67";
                      state_var6679 <= pause_setI5598;
                    end if;
                  when pause_setII5607 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5605\ := \$code_ptr_take\;
                    if \$v5605\(0) = '1' then
                      state_var6679 <= q_wait5604;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 25;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"00000" & X"17");
                      state_var6679 <= pause_setI5602;
                    end if;
                  when pause_setII5611 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5609\ := \$code_ptr_take\;
                    if \$v5609\(0) = '1' then
                      state_var6679 <= q_wait5608;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 24;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"000000" & X"0";
                      state_var6679 <= pause_setI5606;
                    end if;
                  when pause_setII5615 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5613\ := \$code_ptr_take\;
                    if \$v5613\(0) = '1' then
                      state_var6679 <= q_wait5612;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 23;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"000000" & X"1";
                      state_var6679 <= pause_setI5610;
                    end if;
                  when pause_setII5619 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5617\ := \$code_ptr_take\;
                    if \$v5617\(0) = '1' then
                      state_var6679 <= q_wait5616;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 22;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"2c";
                      state_var6679 <= pause_setI5614;
                    end if;
                  when pause_setII5623 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5621\ := \$code_ptr_take\;
                    if \$v5621\(0) = '1' then
                      state_var6679 <= q_wait5620;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 21;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"000000" & X"1";
                      state_var6679 <= pause_setI5618;
                    end if;
                  when pause_setII5627 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5625\ := \$code_ptr_take\;
                    if \$v5625\(0) = '1' then
                      state_var6679 <= q_wait5624;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 20;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"28";
                      state_var6679 <= pause_setI5622;
                    end if;
                  when pause_setII5631 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5629\ := \$code_ptr_take\;
                    if \$v5629\(0) = '1' then
                      state_var6679 <= q_wait5628;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 19;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"6e";
                      state_var6679 <= pause_setI5626;
                    end if;
                  when pause_setII5635 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5633\ := \$code_ptr_take\;
                    if \$v5633\(0) = '1' then
                      state_var6679 <= q_wait5632;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 18;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"21";
                      state_var6679 <= pause_setI5630;
                    end if;
                  when pause_setII5639 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5637\ := \$code_ptr_take\;
                    if \$v5637\(0) = '1' then
                      state_var6679 <= q_wait5636;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 17;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"32";
                      state_var6679 <= pause_setI5634;
                    end if;
                  when pause_setII5643 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5641\ := \$code_ptr_take\;
                    if \$v5641\(0) = '1' then
                      state_var6679 <= q_wait5640;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 16;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"000000" & X"1");
                      state_var6679 <= pause_setI5638;
                    end if;
                  when pause_setII5647 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5645\ := \$code_ptr_take\;
                    if \$v5645\(0) = '1' then
                      state_var6679 <= q_wait5644;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 15;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"7f";
                      state_var6679 <= pause_setI5642;
                    end if;
                  when pause_setII5651 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5649\ := \$code_ptr_take\;
                    if \$v5649\(0) = '1' then
                      state_var6679 <= q_wait5648;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 14;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"000000" & X"b";
                      state_var6679 <= pause_setI5646;
                    end if;
                  when pause_setII5655 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5653\ := \$code_ptr_take\;
                    if \$v5653\(0) = '1' then
                      state_var6679 <= q_wait5652;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 13;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"21";
                      state_var6679 <= pause_setI5650;
                    end if;
                  when pause_setII5659 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5657\ := \$code_ptr_take\;
                    if \$v5657\(0) = '1' then
                      state_var6679 <= q_wait5656;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 12;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"32";
                      state_var6679 <= pause_setI5654;
                    end if;
                  when pause_setII5663 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5661\ := \$code_ptr_take\;
                    if \$v5661\(0) = '1' then
                      state_var6679 <= q_wait5660;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 11;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"000000" & X"2");
                      state_var6679 <= pause_setI5658;
                    end if;
                  when pause_setII5667 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5665\ := \$code_ptr_take\;
                    if \$v5665\(0) = '1' then
                      state_var6679 <= q_wait5664;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 10;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"7f";
                      state_var6679 <= pause_setI5662;
                    end if;
                  when pause_setII5671 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5669\ := \$code_ptr_take\;
                    if \$v5669\(0) = '1' then
                      state_var6679 <= q_wait5668;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 9;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"000000" & X"0";
                      state_var6679 <= pause_setI5666;
                    end if;
                  when pause_setII5675 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5673\ := \$code_ptr_take\;
                    if \$v5673\(0) = '1' then
                      state_var6679 <= q_wait5672;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 8;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"000000" & X"1";
                      state_var6679 <= pause_setI5670;
                    end if;
                  when pause_setII5679 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5677\ := \$code_ptr_take\;
                    if \$v5677\(0) = '1' then
                      state_var6679 <= q_wait5676;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 7;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"28";
                      state_var6679 <= pause_setI5674;
                    end if;
                  when pause_setII5683 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5681\ := \$code_ptr_take\;
                    if \$v5681\(0) = '1' then
                      state_var6679 <= q_wait5680;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 6;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"64";
                      state_var6679 <= pause_setI5678;
                    end if;
                  when pause_setII5687 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5685\ := \$code_ptr_take\;
                    if \$v5685\(0) = '1' then
                      state_var6679 <= q_wait5684;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 5;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"000000" & X"4";
                      state_var6679 <= pause_setI5682;
                    end if;
                  when pause_setII5691 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5689\ := \$code_ptr_take\;
                    if \$v5689\(0) = '1' then
                      state_var6679 <= q_wait5688;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 4;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"000000" & X"2";
                      state_var6679 <= pause_setI5686;
                    end if;
                  when pause_setII5695 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5693\ := \$code_ptr_take\;
                    if \$v5693\(0) = '1' then
                      state_var6679 <= q_wait5692;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 3;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"86";
                      state_var6679 <= pause_setI5690;
                    end if;
                  when pause_setII5699 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5697\ := \$code_ptr_take\;
                    if \$v5697\(0) = '1' then
                      state_var6679 <= q_wait5696;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 2;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"000000" & X"0";
                      state_var6679 <= pause_setI5694;
                    end if;
                  when pause_setII5703 =>
                    \$code_ptr_take\(0) := '0';
                    \$v5701\ := \$code_ptr_take\;
                    if \$v5701\(0) = '1' then
                      state_var6679 <= q_wait5700;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 1;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"15";
                      state_var6679 <= pause_setI5698;
                    end if;
                  when pause_setII5707 =>
                    \$global_end_ptr_take\(0) := '0';
                    \$v5705\ := \$code_ptr_take\;
                    if \$v5705\(0) = '1' then
                      state_var6679 <= q_wait5704;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 0;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"54";
                      state_var6679 <= pause_setI5702;
                    end if;
                  when q_wait5568 =>
                    \$v5569\ := \$code_ptr_take\;
                    if \$v5569\(0) = '1' then
                      state_var6679 <= q_wait5568;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 34;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"8f";
                      state_var6679 <= pause_setI5566;
                    end if;
                  when q_wait5572 =>
                    \$v5573\ := \$code_ptr_take\;
                    if \$v5573\(0) = '1' then
                      state_var6679 <= q_wait5572;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 33;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"000000" & X"1";
                      state_var6679 <= pause_setI5570;
                    end if;
                  when q_wait5576 =>
                    \$v5577\ := \$code_ptr_take\;
                    if \$v5577\(0) = '1' then
                      state_var6679 <= q_wait5576;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 32;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"13";
                      state_var6679 <= pause_setI5574;
                    end if;
                  when q_wait5580 =>
                    \$v5581\ := \$code_ptr_take\;
                    if \$v5581\(0) = '1' then
                      state_var6679 <= q_wait5580;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 31;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"000000" & X"0";
                      state_var6679 <= pause_setI5578;
                    end if;
                  when q_wait5584 =>
                    \$v5585\ := \$code_ptr_take\;
                    if \$v5585\(0) = '1' then
                      state_var6679 <= q_wait5584;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 30;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"5d";
                      state_var6679 <= pause_setI5582;
                    end if;
                  when q_wait5588 =>
                    \$v5589\ := \$code_ptr_take\;
                    if \$v5589\(0) = '1' then
                      state_var6679 <= q_wait5588;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 29;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"21";
                      state_var6679 <= pause_setI5586;
                    end if;
                  when q_wait5592 =>
                    \$v5593\ := \$code_ptr_take\;
                    if \$v5593\(0) = '1' then
                      state_var6679 <= q_wait5592;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 28;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"000000" & X"b";
                      state_var6679 <= pause_setI5590;
                    end if;
                  when q_wait5596 =>
                    \$v5597\ := \$code_ptr_take\;
                    if \$v5597\(0) = '1' then
                      state_var6679 <= q_wait5596;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 27;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"000000" & X"b";
                      state_var6679 <= pause_setI5594;
                    end if;
                  when q_wait5600 =>
                    \$v5601\ := \$code_ptr_take\;
                    if \$v5601\(0) = '1' then
                      state_var6679 <= q_wait5600;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 26;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"67";
                      state_var6679 <= pause_setI5598;
                    end if;
                  when q_wait5604 =>
                    \$v5605\ := \$code_ptr_take\;
                    if \$v5605\(0) = '1' then
                      state_var6679 <= q_wait5604;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 25;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"00000" & X"17");
                      state_var6679 <= pause_setI5602;
                    end if;
                  when q_wait5608 =>
                    \$v5609\ := \$code_ptr_take\;
                    if \$v5609\(0) = '1' then
                      state_var6679 <= q_wait5608;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 24;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"000000" & X"0";
                      state_var6679 <= pause_setI5606;
                    end if;
                  when q_wait5612 =>
                    \$v5613\ := \$code_ptr_take\;
                    if \$v5613\(0) = '1' then
                      state_var6679 <= q_wait5612;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 23;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"000000" & X"1";
                      state_var6679 <= pause_setI5610;
                    end if;
                  when q_wait5616 =>
                    \$v5617\ := \$code_ptr_take\;
                    if \$v5617\(0) = '1' then
                      state_var6679 <= q_wait5616;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 22;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"2c";
                      state_var6679 <= pause_setI5614;
                    end if;
                  when q_wait5620 =>
                    \$v5621\ := \$code_ptr_take\;
                    if \$v5621\(0) = '1' then
                      state_var6679 <= q_wait5620;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 21;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"000000" & X"1";
                      state_var6679 <= pause_setI5618;
                    end if;
                  when q_wait5624 =>
                    \$v5625\ := \$code_ptr_take\;
                    if \$v5625\(0) = '1' then
                      state_var6679 <= q_wait5624;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 20;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"28";
                      state_var6679 <= pause_setI5622;
                    end if;
                  when q_wait5628 =>
                    \$v5629\ := \$code_ptr_take\;
                    if \$v5629\(0) = '1' then
                      state_var6679 <= q_wait5628;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 19;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"6e";
                      state_var6679 <= pause_setI5626;
                    end if;
                  when q_wait5632 =>
                    \$v5633\ := \$code_ptr_take\;
                    if \$v5633\(0) = '1' then
                      state_var6679 <= q_wait5632;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 18;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"21";
                      state_var6679 <= pause_setI5630;
                    end if;
                  when q_wait5636 =>
                    \$v5637\ := \$code_ptr_take\;
                    if \$v5637\(0) = '1' then
                      state_var6679 <= q_wait5636;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 17;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"32";
                      state_var6679 <= pause_setI5634;
                    end if;
                  when q_wait5640 =>
                    \$v5641\ := \$code_ptr_take\;
                    if \$v5641\(0) = '1' then
                      state_var6679 <= q_wait5640;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 16;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"000000" & X"1");
                      state_var6679 <= pause_setI5638;
                    end if;
                  when q_wait5644 =>
                    \$v5645\ := \$code_ptr_take\;
                    if \$v5645\(0) = '1' then
                      state_var6679 <= q_wait5644;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 15;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"7f";
                      state_var6679 <= pause_setI5642;
                    end if;
                  when q_wait5648 =>
                    \$v5649\ := \$code_ptr_take\;
                    if \$v5649\(0) = '1' then
                      state_var6679 <= q_wait5648;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 14;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"000000" & X"b";
                      state_var6679 <= pause_setI5646;
                    end if;
                  when q_wait5652 =>
                    \$v5653\ := \$code_ptr_take\;
                    if \$v5653\(0) = '1' then
                      state_var6679 <= q_wait5652;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 13;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"21";
                      state_var6679 <= pause_setI5650;
                    end if;
                  when q_wait5656 =>
                    \$v5657\ := \$code_ptr_take\;
                    if \$v5657\(0) = '1' then
                      state_var6679 <= q_wait5656;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 12;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"32";
                      state_var6679 <= pause_setI5654;
                    end if;
                  when q_wait5660 =>
                    \$v5661\ := \$code_ptr_take\;
                    if \$v5661\(0) = '1' then
                      state_var6679 <= q_wait5660;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 11;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"000000" & X"2");
                      state_var6679 <= pause_setI5658;
                    end if;
                  when q_wait5664 =>
                    \$v5665\ := \$code_ptr_take\;
                    if \$v5665\(0) = '1' then
                      state_var6679 <= q_wait5664;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 10;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"7f";
                      state_var6679 <= pause_setI5662;
                    end if;
                  when q_wait5668 =>
                    \$v5669\ := \$code_ptr_take\;
                    if \$v5669\(0) = '1' then
                      state_var6679 <= q_wait5668;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 9;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"000000" & X"0";
                      state_var6679 <= pause_setI5666;
                    end if;
                  when q_wait5672 =>
                    \$v5673\ := \$code_ptr_take\;
                    if \$v5673\(0) = '1' then
                      state_var6679 <= q_wait5672;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 8;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"000000" & X"1";
                      state_var6679 <= pause_setI5670;
                    end if;
                  when q_wait5676 =>
                    \$v5677\ := \$code_ptr_take\;
                    if \$v5677\(0) = '1' then
                      state_var6679 <= q_wait5676;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 7;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"28";
                      state_var6679 <= pause_setI5674;
                    end if;
                  when q_wait5680 =>
                    \$v5681\ := \$code_ptr_take\;
                    if \$v5681\(0) = '1' then
                      state_var6679 <= q_wait5680;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 6;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"64";
                      state_var6679 <= pause_setI5678;
                    end if;
                  when q_wait5684 =>
                    \$v5685\ := \$code_ptr_take\;
                    if \$v5685\(0) = '1' then
                      state_var6679 <= q_wait5684;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 5;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"000000" & X"4";
                      state_var6679 <= pause_setI5682;
                    end if;
                  when q_wait5688 =>
                    \$v5689\ := \$code_ptr_take\;
                    if \$v5689\(0) = '1' then
                      state_var6679 <= q_wait5688;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 4;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"000000" & X"2";
                      state_var6679 <= pause_setI5686;
                    end if;
                  when q_wait5692 =>
                    \$v5693\ := \$code_ptr_take\;
                    if \$v5693\(0) = '1' then
                      state_var6679 <= q_wait5692;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 3;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"86";
                      state_var6679 <= pause_setI5690;
                    end if;
                  when q_wait5696 =>
                    \$v5697\ := \$code_ptr_take\;
                    if \$v5697\(0) = '1' then
                      state_var6679 <= q_wait5696;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 2;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"000000" & X"0";
                      state_var6679 <= pause_setI5694;
                    end if;
                  when q_wait5700 =>
                    \$v5701\ := \$code_ptr_take\;
                    if \$v5701\(0) = '1' then
                      state_var6679 <= q_wait5700;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 1;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"15";
                      state_var6679 <= pause_setI5698;
                    end if;
                  when q_wait5704 =>
                    \$v5705\ := \$code_ptr_take\;
                    if \$v5705\(0) = '1' then
                      state_var6679 <= q_wait5704;
                    else
                      \$code_ptr_take\(0) := '1';
                      \$code_ptr_write\ <= 0;
                      \$code_write_request\ <= '1';
                      \$code_write\ <= "000"& X"00000" & X"54";
                      state_var6679 <= pause_setI5702;
                    end if;
                  when q_wait5708 =>
                    \$v5709\ := \$global_end_ptr_take\;
                    if \$v5709\(0) = '1' then
                      state_var6679 <= q_wait5708;
                    else
                      \$global_end_ptr_take\(0) := '1';
                      \$global_end_ptr_write\ <= 0;
                      \$global_end_write_request\ <= '1';
                      \$global_end_write\ <= eclat_add(X"3e80" & X"000" & X"c");
                      state_var6679 <= pause_setI5706;
                    end if;
                  when compute5565 =>
                    rdy5564 := eclat_false;
                    \$v5709\ := \$global_end_ptr_take\;
                    if \$v5709\(0) = '1' then
                      state_var6679 <= q_wait5708;
                    else
                      \$global_end_ptr_take\(0) := '1';
                      \$global_end_ptr_write\ <= 0;
                      \$global_end_write_request\ <= '1';
                      \$global_end_write\ <= eclat_add(X"3e80" & X"000" & X"c");
                      state_var6679 <= pause_setI5706;
                    end if;
                  end case;
                  \$v5711\ := eclat_not(rdy5564);
                  if \$v5711\(0) = '1' then
                    result5563 := eclat_unit;
                  end if;
                  \$14855\ := result5563 & rdy5564;
                  \$v5562\ := eclat_not(rdy5559);
                  if \$v5562\(0) = '1' then
                    \$14859\ := eclat_false;
                  end if;
                  case state_var6678 is
                  when compute5560 =>
                    rdy5559 := eclat_false;
                    \$14859\ := eclat_and(eclat_if(\$14859\ & eclat_true & ""&\$14855\(1)) & eclat_not(eclat_false));
                    rdy5559 := eclat_true;
                    state_var6678 <= compute5560;
                  end case;
                  \$14859\ := \$14859\;
                  \$14858_rdy\ := \$14859\;
                  \$12168\ := eclat_false & eclat_true & \$14858_rdy\ & ""&\$12168\(3);
                  rdy5557 := eclat_true;
                  state_var6673 <= compute5558;
                else
                  \$v6662\ := eclat_not(rdy5712);
                  if \$v6662\(0) = '1' then
                    \$12190\ := X"000" & X"0" & "000"& X"000000" & X"1" & eclat_true & X"0" & X"3e8" & "000"& X"000000" & X"1" & eclat_true & "00000000" & X"000" & X"0" & eclat_false & eclat_false & eclat_true;
                  end if;
                  case state_var6674 is
                  when compute5713 =>
                    rdy5712 := eclat_false;
                    \$v6660\ := eclat_not(""&\$12168\(2));
                    if \$v6660\(0) = '1' then
                      \$12190\ := \$12190\(0 to 121) & eclat_true;
                      rdy5712 := eclat_true;
                      state_var6674 <= compute5713;
                    else
                      case state_var6675 is
                      when \$12199_make_block525\ =>
                        eclat_print_string(of_string("GC-ALLOC:(size="));
                        
                        eclat_print_int(eclat_add(eclat_if(eclat_eq(\$12199_make_block525_arg\(88 to 103) & X"000" & X"0") & X"000" & X"1" & \$12199_make_block525_arg\(88 to 103)) & X"000" & X"1"));
                        
                        eclat_print_string(of_string(")"));
                        
                        eclat_print_newline(eclat_unit);
                        
                        \$14274_wait603_arg\ := eclat_unit & \$12199_make_block525_arg\(16 to 47) & \$12199_make_block525_arg\(48 to 79) & \$12199_make_block525_arg\(0 to 15) & eclat_add(
                        eclat_if(eclat_eq(\$12199_make_block525_arg\(88 to 103) & X"000" & X"0") & X"000" & X"1" & \$12199_make_block525_arg\(88 to 103)) & X"000" & X"1");
                        state_var6675 <= \$14274_wait603\;
                      when \$12235_apply579\ =>
                        eclat_print_string(of_string("ENV:"));
                        
                        eclat_print_int(\$12235_apply579_arg\(110 to 140));
                        
                        eclat_print_string(of_string("<"));
                        
                        \$v5931\ := ""&\$12235_apply579_arg\(141);
                        if \$v5931\(0) = '1' then
                          eclat_print_string(of_string("int"));
                          
                          eclat_print_string(of_string(">"));
                          
                          eclat_print_newline(eclat_unit);
                          
                          \$v5930\ := ""&\$12235_apply579_arg\(0);
                          if \$v5930\(0) = '1' then
                            \$v5929\ := \$ram_ptr_take\;
                            if \$v5929\(0) = '1' then
                              state_var6675 <= q_wait5928;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12235_apply579_arg\(92 to 107) & X"000" & X"1")));
                              state_var6675 <= pause_getI5926;
                            end if;
                          else
                            \$14180\ := "000"& X"000000" & X"1" & eclat_true & \$12235_apply579_arg\(92 to 107);
                            \$v5925\ := ""&\$12235_apply579_arg\(1);
                            if \$v5925\(0) = '1' then
                              \$v5924\ := \$ram_ptr_take\;
                              if \$v5924\(0) = '1' then
                                state_var6675 <= q_wait5923;
                              else
                                \$ram_ptr_take\(0) := '1';
                                \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$14180\(32 to 47) & X"000" & X"1")));
                                state_var6675 <= pause_getI5921;
                              end if;
                            else
                              \$14183\ := "000"& X"000000" & X"1" & eclat_true & \$14180\(32 to 47);
                              \$v5920\ := ""&\$12235_apply579_arg\(2);
                              if \$v5920\(0) = '1' then
                                \$v5919\ := \$ram_ptr_take\;
                                if \$v5919\(0) = '1' then
                                  state_var6675 <= q_wait5918;
                                else
                                  \$ram_ptr_take\(0) := '1';
                                  \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$14183\(32 to 47) & X"000" & X"1")));
                                  state_var6675 <= pause_getI5916;
                                end if;
                              else
                                \$14186\ := "000"& X"000000" & X"1" & eclat_true & \$14183\(32 to 47);
                                \$v5915\ := ""&\$12235_apply579_arg\(11);
                                if \$v5915\(0) = '1' then
                                  \$14189_sp\ := eclat_add(eclat_sub(\$14186\(32 to 47) & \$12235_apply579_arg\(12 to 27)) & \$12235_apply579_arg\(28 to 43));
                                  \$v5902\ := ""&\$12235_apply579_arg\(2);
                                  if \$v5902\(0) = '1' then
                                    \$v5901\ := \$ram_ptr_take\;
                                    if \$v5901\(0) = '1' then
                                      state_var6675 <= q_wait5900;
                                    else
                                      \$ram_ptr_take\(0) := '1';
                                      \$ram_ptr_write\ <= to_integer(unsigned(\$14189_sp\));
                                      \$ram_write_request\ <= '1';
                                      \$ram_write\ <= \$14186\(0 to 31);
                                      state_var6675 <= pause_setI5898;
                                    end if;
                                  else
                                    \$14190_sp\ := \$14189_sp\;
                                    \$v5897\ := ""&\$12235_apply579_arg\(1);
                                    if \$v5897\(0) = '1' then
                                      \$v5896\ := \$ram_ptr_take\;
                                      if \$v5896\(0) = '1' then
                                        state_var6675 <= q_wait5895;
                                      else
                                        \$ram_ptr_take\(0) := '1';
                                        \$ram_ptr_write\ <= to_integer(unsigned(\$14190_sp\));
                                        \$ram_write_request\ <= '1';
                                        \$ram_write\ <= \$14183\(0 to 31);
                                        state_var6675 <= pause_setI5893;
                                      end if;
                                    else
                                      \$14191_sp\ := \$14190_sp\;
                                      \$v5892\ := ""&\$12235_apply579_arg\(0);
                                      if \$v5892\(0) = '1' then
                                        \$v5891\ := \$ram_ptr_take\;
                                        if \$v5891\(0) = '1' then
                                          state_var6675 <= q_wait5890;
                                        else
                                          \$ram_ptr_take\(0) := '1';
                                          \$ram_ptr_write\ <= to_integer(unsigned(\$14191_sp\));
                                          \$ram_write_request\ <= '1';
                                          \$ram_write\ <= \$14180\(0 to 31);
                                          state_var6675 <= pause_setI5888;
                                        end if;
                                      else
                                        \$14192_sp\ := \$14191_sp\;
                                        \$v5887\ := \$ram_ptr_take\;
                                        if \$v5887\(0) = '1' then
                                          state_var6675 <= q_wait5886;
                                        else
                                          \$ram_ptr_take\(0) := '1';
                                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12235_apply579_arg\(60 to 90),16) & X"000" & X"0") & X"000" & X"1")));
                                          state_var6675 <= pause_getI5884;
                                        end if;
                                      end if;
                                    end if;
                                  end if;
                                else
                                  \$v5914\ := \$ram_ptr_take\;
                                  if \$v5914\(0) = '1' then
                                    state_var6675 <= q_wait5913;
                                  else
                                    \$ram_ptr_take\(0) := '1';
                                    \$ram_ptr_write\ <= to_integer(unsigned(\$14186\(32 to 47)));
                                    \$ram_write_request\ <= '1';
                                    \$ram_write\ <= eclat_resize(\$12235_apply579_arg\(142 to 149),31) & eclat_true;
                                    state_var6675 <= pause_setI5911;
                                  end if;
                                end if;
                              end if;
                            end if;
                          end if;
                        else
                          eclat_print_string(of_string("ptr"));
                          
                          eclat_print_string(of_string(">"));
                          
                          eclat_print_newline(eclat_unit);
                          
                          \$v5930\ := ""&\$12235_apply579_arg\(0);
                          if \$v5930\(0) = '1' then
                            \$v5929\ := \$ram_ptr_take\;
                            if \$v5929\(0) = '1' then
                              state_var6675 <= q_wait5928;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12235_apply579_arg\(92 to 107) & X"000" & X"1")));
                              state_var6675 <= pause_getI5926;
                            end if;
                          else
                            \$14180\ := "000"& X"000000" & X"1" & eclat_true & \$12235_apply579_arg\(92 to 107);
                            \$v5925\ := ""&\$12235_apply579_arg\(1);
                            if \$v5925\(0) = '1' then
                              \$v5924\ := \$ram_ptr_take\;
                              if \$v5924\(0) = '1' then
                                state_var6675 <= q_wait5923;
                              else
                                \$ram_ptr_take\(0) := '1';
                                \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$14180\(32 to 47) & X"000" & X"1")));
                                state_var6675 <= pause_getI5921;
                              end if;
                            else
                              \$14183\ := "000"& X"000000" & X"1" & eclat_true & \$14180\(32 to 47);
                              \$v5920\ := ""&\$12235_apply579_arg\(2);
                              if \$v5920\(0) = '1' then
                                \$v5919\ := \$ram_ptr_take\;
                                if \$v5919\(0) = '1' then
                                  state_var6675 <= q_wait5918;
                                else
                                  \$ram_ptr_take\(0) := '1';
                                  \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$14183\(32 to 47) & X"000" & X"1")));
                                  state_var6675 <= pause_getI5916;
                                end if;
                              else
                                \$14186\ := "000"& X"000000" & X"1" & eclat_true & \$14183\(32 to 47);
                                \$v5915\ := ""&\$12235_apply579_arg\(11);
                                if \$v5915\(0) = '1' then
                                  \$14189_sp\ := eclat_add(eclat_sub(\$14186\(32 to 47) & \$12235_apply579_arg\(12 to 27)) & \$12235_apply579_arg\(28 to 43));
                                  \$v5902\ := ""&\$12235_apply579_arg\(2);
                                  if \$v5902\(0) = '1' then
                                    \$v5901\ := \$ram_ptr_take\;
                                    if \$v5901\(0) = '1' then
                                      state_var6675 <= q_wait5900;
                                    else
                                      \$ram_ptr_take\(0) := '1';
                                      \$ram_ptr_write\ <= to_integer(unsigned(\$14189_sp\));
                                      \$ram_write_request\ <= '1';
                                      \$ram_write\ <= \$14186\(0 to 31);
                                      state_var6675 <= pause_setI5898;
                                    end if;
                                  else
                                    \$14190_sp\ := \$14189_sp\;
                                    \$v5897\ := ""&\$12235_apply579_arg\(1);
                                    if \$v5897\(0) = '1' then
                                      \$v5896\ := \$ram_ptr_take\;
                                      if \$v5896\(0) = '1' then
                                        state_var6675 <= q_wait5895;
                                      else
                                        \$ram_ptr_take\(0) := '1';
                                        \$ram_ptr_write\ <= to_integer(unsigned(\$14190_sp\));
                                        \$ram_write_request\ <= '1';
                                        \$ram_write\ <= \$14183\(0 to 31);
                                        state_var6675 <= pause_setI5893;
                                      end if;
                                    else
                                      \$14191_sp\ := \$14190_sp\;
                                      \$v5892\ := ""&\$12235_apply579_arg\(0);
                                      if \$v5892\(0) = '1' then
                                        \$v5891\ := \$ram_ptr_take\;
                                        if \$v5891\(0) = '1' then
                                          state_var6675 <= q_wait5890;
                                        else
                                          \$ram_ptr_take\(0) := '1';
                                          \$ram_ptr_write\ <= to_integer(unsigned(\$14191_sp\));
                                          \$ram_write_request\ <= '1';
                                          \$ram_write\ <= \$14180\(0 to 31);
                                          state_var6675 <= pause_setI5888;
                                        end if;
                                      else
                                        \$14192_sp\ := \$14191_sp\;
                                        \$v5887\ := \$ram_ptr_take\;
                                        if \$v5887\(0) = '1' then
                                          state_var6675 <= q_wait5886;
                                        else
                                          \$ram_ptr_take\(0) := '1';
                                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12235_apply579_arg\(60 to 90),16) & X"000" & X"0") & X"000" & X"1")));
                                          state_var6675 <= pause_getI5884;
                                        end if;
                                      end if;
                                    end if;
                                  end if;
                                else
                                  \$v5914\ := \$ram_ptr_take\;
                                  if \$v5914\(0) = '1' then
                                    state_var6675 <= q_wait5913;
                                  else
                                    \$ram_ptr_take\(0) := '1';
                                    \$ram_ptr_write\ <= to_integer(unsigned(\$14186\(32 to 47)));
                                    \$ram_write_request\ <= '1';
                                    \$ram_write\ <= eclat_resize(\$12235_apply579_arg\(142 to 149),31) & eclat_true;
                                    state_var6675 <= pause_setI5911;
                                  end if;
                                end if;
                              end if;
                            end if;
                          end if;
                        end if;
                      when \$12236_offsetclosure_n580\ =>
                        \$12236_offsetclosure_n580_result\ := \$12236_offsetclosure_n580_arg\(0 to 15) & eclat_resize(eclat_add(eclat_resize(\$12236_offsetclosure_n580_arg\(106 to 136),16) & \$12236_offsetclosure_n580_arg\(32 to 47)),31) & eclat_false & \$12236_offsetclosure_n580_arg\(16 to 31) & \$12236_offsetclosure_n580_arg\(48 to 103) & \$12236_offsetclosure_n580_arg\(104 to 105);
                        result5714 := \$12236_offsetclosure_n580_result\;
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when \$12237_binop_int584\ =>
                        \$v5940\ := \$ram_ptr_take\;
                        if \$v5940\(0) = '1' then
                          state_var6675 <= q_wait5939;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12237_binop_int584_arg\(80 to 95) & X"000" & X"1")));
                          state_var6675 <= pause_getI5937;
                        end if;
                      when \$12238_compare585\ =>
                        \$v5941\ := \$12238_compare585_arg\(0 to 31);
                        case \$v5941\ is
                        when X"0000000" & X"0" =>
                          \$12238_compare585_result\ := eclat_eq(\$12238_compare585_arg\(32 to 62) & \$12238_compare585_arg\(63 to 93));
                          case \$12238_compare585_id\ is
                          when "000000001101" =>
                            \$14052_res\ := \$12238_compare585_result\;
                            \$12239_binop_compare586_result\ := eclat_add(\$12239_binop_compare586_arg\(32 to 47) & X"000" & X"1") & 
                            eclat_if(\$14052_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & eclat_sub(\$12239_binop_compare586_arg\(80 to 95) & X"000" & X"1") & \$12239_binop_compare586_arg\(96 to 151) & \$12239_binop_compare586_arg\(152 to 153);
                            result5714 := \$12239_binop_compare586_result\;
                            rdy5715 := eclat_true;
                            state_var6675 <= compute5716;
                          when "000000110011" =>
                            \$13322_b\ := \$12238_compare585_result\;
                            \$12245_compbranch590_result\ := eclat_if(\$13322_b\ & eclat_add(eclat_add(\$12245_compbranch590_arg\(94 to 109) & X"000" & X"2") & eclat_resize(\$12245_compbranch590_arg\(63 to 93),16)) & \$12245_compbranch590_arg\(110 to 141) & \$12245_compbranch590_arg\(142 to 157) & \$12245_compbranch590_arg\(158 to 213) & \$12245_compbranch590_arg\(214 to 215) & eclat_add(\$12245_compbranch590_arg\(94 to 109) & X"000" & X"3") & \$12245_compbranch590_arg\(110 to 141) & \$12245_compbranch590_arg\(142 to 157) & \$12245_compbranch590_arg\(158 to 213) & \$12245_compbranch590_arg\(214 to 215));
                            result5714 := \$12245_compbranch590_result\;
                            rdy5715 := eclat_true;
                            state_var6675 <= compute5716;
                          when others =>
                            
                          end case;
                        when X"0000000" & X"1" =>
                          \$12238_compare585_result\ := eclat_not(eclat_eq(\$12238_compare585_arg\(32 to 62) & \$12238_compare585_arg\(63 to 93)));
                          case \$12238_compare585_id\ is
                          when "000000001101" =>
                            \$14052_res\ := \$12238_compare585_result\;
                            \$12239_binop_compare586_result\ := eclat_add(\$12239_binop_compare586_arg\(32 to 47) & X"000" & X"1") & 
                            eclat_if(\$14052_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & eclat_sub(\$12239_binop_compare586_arg\(80 to 95) & X"000" & X"1") & \$12239_binop_compare586_arg\(96 to 151) & \$12239_binop_compare586_arg\(152 to 153);
                            result5714 := \$12239_binop_compare586_result\;
                            rdy5715 := eclat_true;
                            state_var6675 <= compute5716;
                          when "000000110011" =>
                            \$13322_b\ := \$12238_compare585_result\;
                            \$12245_compbranch590_result\ := eclat_if(\$13322_b\ & eclat_add(eclat_add(\$12245_compbranch590_arg\(94 to 109) & X"000" & X"2") & eclat_resize(\$12245_compbranch590_arg\(63 to 93),16)) & \$12245_compbranch590_arg\(110 to 141) & \$12245_compbranch590_arg\(142 to 157) & \$12245_compbranch590_arg\(158 to 213) & \$12245_compbranch590_arg\(214 to 215) & eclat_add(\$12245_compbranch590_arg\(94 to 109) & X"000" & X"3") & \$12245_compbranch590_arg\(110 to 141) & \$12245_compbranch590_arg\(142 to 157) & \$12245_compbranch590_arg\(158 to 213) & \$12245_compbranch590_arg\(214 to 215));
                            result5714 := \$12245_compbranch590_result\;
                            rdy5715 := eclat_true;
                            state_var6675 <= compute5716;
                          when others =>
                            
                          end case;
                        when X"0000000" & X"2" =>
                          \$12238_compare585_result\ := eclat_lt(\$12238_compare585_arg\(32 to 62) & \$12238_compare585_arg\(63 to 93));
                          case \$12238_compare585_id\ is
                          when "000000001101" =>
                            \$14052_res\ := \$12238_compare585_result\;
                            \$12239_binop_compare586_result\ := eclat_add(\$12239_binop_compare586_arg\(32 to 47) & X"000" & X"1") & 
                            eclat_if(\$14052_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & eclat_sub(\$12239_binop_compare586_arg\(80 to 95) & X"000" & X"1") & \$12239_binop_compare586_arg\(96 to 151) & \$12239_binop_compare586_arg\(152 to 153);
                            result5714 := \$12239_binop_compare586_result\;
                            rdy5715 := eclat_true;
                            state_var6675 <= compute5716;
                          when "000000110011" =>
                            \$13322_b\ := \$12238_compare585_result\;
                            \$12245_compbranch590_result\ := eclat_if(\$13322_b\ & eclat_add(eclat_add(\$12245_compbranch590_arg\(94 to 109) & X"000" & X"2") & eclat_resize(\$12245_compbranch590_arg\(63 to 93),16)) & \$12245_compbranch590_arg\(110 to 141) & \$12245_compbranch590_arg\(142 to 157) & \$12245_compbranch590_arg\(158 to 213) & \$12245_compbranch590_arg\(214 to 215) & eclat_add(\$12245_compbranch590_arg\(94 to 109) & X"000" & X"3") & \$12245_compbranch590_arg\(110 to 141) & \$12245_compbranch590_arg\(142 to 157) & \$12245_compbranch590_arg\(158 to 213) & \$12245_compbranch590_arg\(214 to 215));
                            result5714 := \$12245_compbranch590_result\;
                            rdy5715 := eclat_true;
                            state_var6675 <= compute5716;
                          when others =>
                            
                          end case;
                        when X"0000000" & X"3" =>
                          \$12238_compare585_result\ := eclat_if(eclat_lt(\$12238_compare585_arg\(32 to 62) & \$12238_compare585_arg\(63 to 93)) & eclat_true & eclat_eq(\$12238_compare585_arg\(32 to 62) & \$12238_compare585_arg\(63 to 93)));
                          case \$12238_compare585_id\ is
                          when "000000001101" =>
                            \$14052_res\ := \$12238_compare585_result\;
                            \$12239_binop_compare586_result\ := eclat_add(\$12239_binop_compare586_arg\(32 to 47) & X"000" & X"1") & 
                            eclat_if(\$14052_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & eclat_sub(\$12239_binop_compare586_arg\(80 to 95) & X"000" & X"1") & \$12239_binop_compare586_arg\(96 to 151) & \$12239_binop_compare586_arg\(152 to 153);
                            result5714 := \$12239_binop_compare586_result\;
                            rdy5715 := eclat_true;
                            state_var6675 <= compute5716;
                          when "000000110011" =>
                            \$13322_b\ := \$12238_compare585_result\;
                            \$12245_compbranch590_result\ := eclat_if(\$13322_b\ & eclat_add(eclat_add(\$12245_compbranch590_arg\(94 to 109) & X"000" & X"2") & eclat_resize(\$12245_compbranch590_arg\(63 to 93),16)) & \$12245_compbranch590_arg\(110 to 141) & \$12245_compbranch590_arg\(142 to 157) & \$12245_compbranch590_arg\(158 to 213) & \$12245_compbranch590_arg\(214 to 215) & eclat_add(\$12245_compbranch590_arg\(94 to 109) & X"000" & X"3") & \$12245_compbranch590_arg\(110 to 141) & \$12245_compbranch590_arg\(142 to 157) & \$12245_compbranch590_arg\(158 to 213) & \$12245_compbranch590_arg\(214 to 215));
                            result5714 := \$12245_compbranch590_result\;
                            rdy5715 := eclat_true;
                            state_var6675 <= compute5716;
                          when others =>
                            
                          end case;
                        when X"0000000" & X"4" =>
                          \$12238_compare585_result\ := eclat_not(eclat_if(eclat_lt(\$12238_compare585_arg\(32 to 62) & \$12238_compare585_arg\(63 to 93)) & eclat_true & eclat_eq(\$12238_compare585_arg\(32 to 62) & \$12238_compare585_arg\(63 to 93))));
                          case \$12238_compare585_id\ is
                          when "000000001101" =>
                            \$14052_res\ := \$12238_compare585_result\;
                            \$12239_binop_compare586_result\ := eclat_add(\$12239_binop_compare586_arg\(32 to 47) & X"000" & X"1") & 
                            eclat_if(\$14052_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & eclat_sub(\$12239_binop_compare586_arg\(80 to 95) & X"000" & X"1") & \$12239_binop_compare586_arg\(96 to 151) & \$12239_binop_compare586_arg\(152 to 153);
                            result5714 := \$12239_binop_compare586_result\;
                            rdy5715 := eclat_true;
                            state_var6675 <= compute5716;
                          when "000000110011" =>
                            \$13322_b\ := \$12238_compare585_result\;
                            \$12245_compbranch590_result\ := eclat_if(\$13322_b\ & eclat_add(eclat_add(\$12245_compbranch590_arg\(94 to 109) & X"000" & X"2") & eclat_resize(\$12245_compbranch590_arg\(63 to 93),16)) & \$12245_compbranch590_arg\(110 to 141) & \$12245_compbranch590_arg\(142 to 157) & \$12245_compbranch590_arg\(158 to 213) & \$12245_compbranch590_arg\(214 to 215) & eclat_add(\$12245_compbranch590_arg\(94 to 109) & X"000" & X"3") & \$12245_compbranch590_arg\(110 to 141) & \$12245_compbranch590_arg\(142 to 157) & \$12245_compbranch590_arg\(158 to 213) & \$12245_compbranch590_arg\(214 to 215));
                            result5714 := \$12245_compbranch590_result\;
                            rdy5715 := eclat_true;
                            state_var6675 <= compute5716;
                          when others =>
                            
                          end case;
                        when X"0000000" & X"5" =>
                          \$12238_compare585_result\ := eclat_not(eclat_lt(\$12238_compare585_arg\(32 to 62) & \$12238_compare585_arg\(63 to 93)));
                          case \$12238_compare585_id\ is
                          when "000000001101" =>
                            \$14052_res\ := \$12238_compare585_result\;
                            \$12239_binop_compare586_result\ := eclat_add(\$12239_binop_compare586_arg\(32 to 47) & X"000" & X"1") & 
                            eclat_if(\$14052_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & eclat_sub(\$12239_binop_compare586_arg\(80 to 95) & X"000" & X"1") & \$12239_binop_compare586_arg\(96 to 151) & \$12239_binop_compare586_arg\(152 to 153);
                            result5714 := \$12239_binop_compare586_result\;
                            rdy5715 := eclat_true;
                            state_var6675 <= compute5716;
                          when "000000110011" =>
                            \$13322_b\ := \$12238_compare585_result\;
                            \$12245_compbranch590_result\ := eclat_if(\$13322_b\ & eclat_add(eclat_add(\$12245_compbranch590_arg\(94 to 109) & X"000" & X"2") & eclat_resize(\$12245_compbranch590_arg\(63 to 93),16)) & \$12245_compbranch590_arg\(110 to 141) & \$12245_compbranch590_arg\(142 to 157) & \$12245_compbranch590_arg\(158 to 213) & \$12245_compbranch590_arg\(214 to 215) & eclat_add(\$12245_compbranch590_arg\(94 to 109) & X"000" & X"3") & \$12245_compbranch590_arg\(110 to 141) & \$12245_compbranch590_arg\(142 to 157) & \$12245_compbranch590_arg\(158 to 213) & \$12245_compbranch590_arg\(214 to 215));
                            result5714 := \$12245_compbranch590_result\;
                            rdy5715 := eclat_true;
                            state_var6675 <= compute5716;
                          when others =>
                            
                          end case;
                        when others =>
                          \$12238_compare585_result\ := eclat_false;
                          case \$12238_compare585_id\ is
                          when "000000001101" =>
                            \$14052_res\ := \$12238_compare585_result\;
                            \$12239_binop_compare586_result\ := eclat_add(\$12239_binop_compare586_arg\(32 to 47) & X"000" & X"1") & 
                            eclat_if(\$14052_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & eclat_sub(\$12239_binop_compare586_arg\(80 to 95) & X"000" & X"1") & \$12239_binop_compare586_arg\(96 to 151) & \$12239_binop_compare586_arg\(152 to 153);
                            result5714 := \$12239_binop_compare586_result\;
                            rdy5715 := eclat_true;
                            state_var6675 <= compute5716;
                          when "000000110011" =>
                            \$13322_b\ := \$12238_compare585_result\;
                            \$12245_compbranch590_result\ := eclat_if(\$13322_b\ & eclat_add(eclat_add(\$12245_compbranch590_arg\(94 to 109) & X"000" & X"2") & eclat_resize(\$12245_compbranch590_arg\(63 to 93),16)) & \$12245_compbranch590_arg\(110 to 141) & \$12245_compbranch590_arg\(142 to 157) & \$12245_compbranch590_arg\(158 to 213) & \$12245_compbranch590_arg\(214 to 215) & eclat_add(\$12245_compbranch590_arg\(94 to 109) & X"000" & X"3") & \$12245_compbranch590_arg\(110 to 141) & \$12245_compbranch590_arg\(142 to 157) & \$12245_compbranch590_arg\(158 to 213) & \$12245_compbranch590_arg\(214 to 215));
                            result5714 := \$12245_compbranch590_result\;
                            rdy5715 := eclat_true;
                            state_var6675 <= compute5716;
                          when others =>
                            
                          end case;
                        end case;
                      when \$12239_binop_compare586\ =>
                        \$v5945\ := \$ram_ptr_take\;
                        if \$v5945\(0) = '1' then
                          state_var6675 <= q_wait5944;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12239_binop_compare586_arg\(80 to 95) & X"000" & X"1")));
                          state_var6675 <= pause_getI5942;
                        end if;
                      when \$12240_make_block_n587\ =>
                        \$12199_make_block525_id\ := "000000001110";
                        \$12199_make_block525_arg\ := \$12240_make_block_n587_arg\(16 to 31) & \$12240_make_block_n587_arg\(82 to 113) & \$12240_make_block_n587_arg\(116 to 147) & eclat_resize(\$12240_make_block_n587_arg\(35 to 65),8) & \$12240_make_block_n587_arg\(66 to 81);
                        state_var6675 <= \$12199_make_block525\;
                      when \$12241_branch_if589\ =>
                        \$v5973\ := eclat_if(""&\$12241_branch_if589_arg\(0) & eclat_not(eclat_neq(\$12241_branch_if589_arg\(17 to 47) & "000"& X"000000" & X"0")) & eclat_neq(\$12241_branch_if589_arg\(17 to 47) & "000"& X"000000" & X"0"));
                        if \$v5973\(0) = '1' then
                          \$v5972\ := \$code_ptr_take\;
                          if \$v5972\(0) = '1' then
                            state_var6675 <= q_wait5971;
                          else
                            \$code_ptr_take\(0) := '1';
                            \$code_ptr\ <= to_integer(unsigned(eclat_add(\$12241_branch_if589_arg\(1 to 16) & X"000" & X"1")));
                            state_var6675 <= pause_getI5969;
                          end if;
                        else
                          \$12241_branch_if589_result\ := eclat_add(\$12241_branch_if589_arg\(1 to 16) & X"000" & X"2") & \$12241_branch_if589_arg\(17 to 48) & \$12241_branch_if589_arg\(49 to 64) & \$12241_branch_if589_arg\(65 to 120) & \$12241_branch_if589_arg\(121 to 122);
                          result5714 := \$12241_branch_if589_result\;
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        end if;
                      when \$12245_compbranch590\ =>
                        \$12238_compare585_id\ := "000000110011";
                        \$12238_compare585_arg\ := \$12245_compbranch590_arg\(0 to 31) & \$12245_compbranch590_arg\(32 to 62) & \$12245_compbranch590_arg\(110 to 140);
                        state_var6675 <= \$12238_compare585\;
                      when \$12265_w0591\ =>
                        \$v6600\ := eclat_ge(\$12265_w0591_arg\(0 to 15) & \$12265_w0591_arg\(48 to 63));
                        if \$v6600\(0) = '1' then
                          \$12265_w0591_result\ := \$12265_w0591_arg\(16 to 31);
                          \$12266_sp\ := \$12265_w0591_result\;
                          \$12267_w1592_arg\ := X"000" & X"1" & \$12190\(0 to 15) & eclat_resize(\$12246_argument1\,16) & \$12257\(64 to 95);
                          state_var6675 <= \$12267_w1592\;
                        else
                          \$v6599\ := \$ram_ptr_take\;
                          if \$v6599\(0) = '1' then
                            state_var6675 <= q_wait6598;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12265_w0591_arg\(16 to 31) & X"000" & X"1")));
                            state_var6675 <= pause_getI6596;
                          end if;
                        end if;
                      when \$12267_w1592\ =>
                        \$v6613\ := eclat_ge(\$12267_w1592_arg\(0 to 15) & \$12267_w1592_arg\(32 to 47));
                        if \$v6613\(0) = '1' then
                          \$12267_w1592_result\ := eclat_unit;
                          \$v6622\ := \$ram_ptr_take\;
                          if \$v6622\(0) = '1' then
                            state_var6675 <= q_wait6621;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12266_sp\));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12257\(64 to 95);
                            state_var6675 <= pause_setI6619;
                          end if;
                        else
                          \$v6612\ := \$ram_ptr_take\;
                          if \$v6612\(0) = '1' then
                            state_var6675 <= q_wait6611;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12267_w1592_arg\(48 to 78),16) & eclat_sub(eclat_mult(X"000" & X"2" & \$12267_w1592_arg\(0 to 15)) & X"000" & X"1")) & X"000" & X"1")));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= eclat_lor(eclat_lsl(eclat_resize("11111001",31) & "000"& X"00000" & X"18") & eclat_lsl(eclat_resize(eclat_mult(X"000" & X"2" & \$12267_w1592_arg\(0 to 15)),31) & "000"& X"000000" & X"2")) & eclat_true;
                            state_var6675 <= pause_setI6609;
                          end if;
                        end if;
                      when \$12270_w3593\ =>
                        \$v6618\ := eclat_ge(\$12270_w3593_arg\(0 to 15) & \$12270_w3593_arg\(32 to 47));
                        if \$v6618\(0) = '1' then
                          \$12270_w3593_result\ := \$12270_w3593_arg\(16 to 31);
                          \$12271_sp\ := \$12270_w3593_result\;
                          result5714 := eclat_add(eclat_add(\$12190\(0 to 15) & X"000" & X"3") & eclat_resize(\$12246_argument1\,16)) & \$12257\(64 to 95) & \$12271_sp\ & \$12257\(32 to 63) & \$12190\(96 to 103) & \$12190\(104 to 119) & \$12190\(120 to 121);
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        else
                          \$v6617\ := \$ram_ptr_take\;
                          if \$v6617\(0) = '1' then
                            state_var6675 <= q_wait6616;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12270_w3593_arg\(16 to 31)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= eclat_resize(eclat_add(eclat_resize(\$12270_w3593_arg\(48 to 78),16) & eclat_mult(X"000" & X"2" & \$12270_w3593_arg\(0 to 15))),31) & eclat_true;
                            state_var6675 <= pause_setI6614;
                          end if;
                        end if;
                      when \$12421_w594\ =>
                        \$v6536\ := eclat_gt(\$12421_w594_arg\(0 to 15) & \$12421_w594_arg\(32 to 47));
                        if \$v6536\(0) = '1' then
                          \$12421_w594_result\ := eclat_unit;
                          \$v6540\ := \$ram_ptr_take\;
                          if \$v6540\(0) = '1' then
                            state_var6675 <= q_wait6539;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & X"000" & X"0") & X"000" & X"1")));
                            state_var6675 <= pause_getI6537;
                          end if;
                        else
                          \$v6535\ := \$ram_ptr_take\;
                          if \$v6535\(0) = '1' then
                            state_var6675 <= q_wait6534;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12421_w594_arg\(16 to 31) & \$12421_w594_arg\(0 to 15))));
                            state_var6675 <= pause_getI6532;
                          end if;
                        end if;
                      when \$12474_fill595\ =>
                        \$v6549\ := eclat_gt(\$12474_fill595_arg\(0 to 15) & \$12474_fill595_arg\(32 to 47));
                        if \$v6549\(0) = '1' then
                          \$12474_fill595_result\ := \$12474_fill595_arg\(16 to 31);
                          \$12475_sp\ := \$12474_fill595_result\;
                          result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"3") & \$12466\(64 to 95) & \$12475_sp\ & \$12466\(32 to 63) & \$12190\(96 to 103) & \$12190\(104 to 119) & \$12190\(120 to 121);
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        else
                          \$v6548\ := \$ram_ptr_take\;
                          if \$v6548\(0) = '1' then
                            state_var6675 <= q_wait6547;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12474_fill595_arg\(16 to 31) & X"000" & X"1")));
                            state_var6675 <= pause_getI6545;
                          end if;
                        end if;
                      when \$12564_fill596\ =>
                        \$v6587\ := eclat_ge(\$12564_fill596_arg\(0 to 15) & \$12564_fill596_arg\(32 to 47));
                        if \$v6587\(0) = '1' then
                          \$12564_fill596_result\ := \$12564_fill596_arg\(16 to 31);
                          \$12565_sp\ := \$12564_fill596_result\;
                          result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"3") & \$12556\(64 to 95) & \$12565_sp\ & \$12556\(32 to 63) & \$12190\(96 to 103) & \$12190\(104 to 119) & \$12190\(120 to 121);
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        else
                          \$v6586\ := \$ram_ptr_take\;
                          if \$v6586\(0) = '1' then
                            state_var6675 <= q_wait6585;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12564_fill596_arg\(16 to 31) & X"000" & X"1")));
                            state_var6675 <= pause_getI6583;
                          end if;
                        end if;
                      when \$12782_w597\ =>
                        \$v6348\ := eclat_gt(\$12782_w597_arg\(0 to 7) & \$12782_w597_arg\(24 to 31));
                        if \$v6348\(0) = '1' then
                          \$12782_w597_result\ := \$12782_w597_arg\(8 to 23);
                          \$12783_sp\ := \$12782_w597_result\;
                          \$v6360\ := \$ram_ptr_take\;
                          if \$v6360\(0) = '1' then
                            state_var6675 <= q_wait6359;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12783_sp\ & X"000" & X"1")));
                            state_var6675 <= pause_getI6357;
                          end if;
                        else
                          \$v6347\ := \$ram_ptr_take\;
                          if \$v6347\(0) = '1' then
                            state_var6675 <= q_wait6346;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12782_w597_arg\(8 to 23) & X"000" & X"1")));
                            state_var6675 <= pause_getI6344;
                          end if;
                        end if;
                      when \$12909_forever611\ =>
                        state_var6675 <= \$12909_forever611\;
                      when \$12946_forever611\ =>
                        state_var6675 <= \$12946_forever611\;
                      when \$13261_forever611\ =>
                        state_var6675 <= \$13261_forever611\;
                      when \$13539_loop_push598\ =>
                        \$v6126\ := eclat_ge(\$13539_loop_push598_arg\(16 to 23) & eclat_sub(\$13539_loop_push598_arg\(56 to 63) & "00000010"));
                        if \$v6126\(0) = '1' then
                          \$13539_loop_push598_result\ := \$13539_loop_push598_arg\(0 to 15);
                          \$13543_sp\ := \$13539_loop_push598_result\;
                          \$v6130\ := \$ram_ptr_take\;
                          if \$v6130\(0) = '1' then
                            state_var6675 <= q_wait6129;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(64 to 94),16) & X"000" & X"1") & X"000" & X"1")));
                            state_var6675 <= pause_getI6127;
                          end if;
                        else
                          \$v6125\ := \$ram_ptr_take\;
                          if \$v6125\(0) = '1' then
                            state_var6675 <= q_wait6124;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$13539_loop_push598_arg\(24 to 54),16) & eclat_resize(eclat_add(\$13539_loop_push598_arg\(16 to 23) & "00000010"),16)) & X"000" & X"1")));
                            state_var6675 <= pause_getI6122;
                          end if;
                        end if;
                      when \$13928_forever611\ =>
                        state_var6675 <= \$13928_forever611\;
                      when \$13935_forever611\ =>
                        state_var6675 <= \$13935_forever611\;
                      when \$13942_forever611\ =>
                        state_var6675 <= \$13942_forever611\;
                      when \$14090_modulo609\ =>
                        \$v5932\ := eclat_lt(\$14090_modulo609_arg\(0 to 30) & \$14090_modulo609_arg\(31 to 61));
                        if \$v5932\(0) = '1' then
                          \$14090_modulo609_result\ := \$14090_modulo609_arg\(0 to 30);
                          \$14091_r\ := \$14090_modulo609_result\;
                          \$14086_res\ := eclat_if(eclat_lt(\$12237_binop_int584_arg\(48 to 78) & "000"& X"000000" & X"0") & eclat_sub("000"& X"000000" & X"0" & \$14091_r\) & \$14091_r\);
                          \$12237_binop_int584_result\ := eclat_add(\$12237_binop_int584_arg\(32 to 47) & X"000" & X"1") & \$14086_res\ & eclat_true & eclat_sub(\$12237_binop_int584_arg\(80 to 95) & X"000" & X"1") & \$12237_binop_int584_arg\(96 to 151) & \$12237_binop_int584_arg\(152 to 153);
                          result5714 := \$12237_binop_int584_result\;
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        else
                          \$14090_modulo609_arg\ := eclat_sub(\$14090_modulo609_arg\(0 to 30) & \$14090_modulo609_arg\(31 to 61)) & \$14090_modulo609_arg\(31 to 61);
                          state_var6675 <= \$14090_modulo609\;
                        end if;
                      when \$14105_modulo609\ =>
                        \$v5934\ := eclat_lt(\$14105_modulo609_arg\(0 to 30) & \$14105_modulo609_arg\(31 to 61));
                        if \$v5934\(0) = '1' then
                          \$14105_modulo609_result\ := \$14105_modulo609_arg\(0 to 30);
                          \$14106_r\ := \$14105_modulo609_result\;
                          \$14086_res\ := eclat_if(eclat_lt(\$12237_binop_int584_arg\(48 to 78) & "000"& X"000000" & X"0") & eclat_sub("000"& X"000000" & X"0" & \$14106_r\) & \$14106_r\);
                          \$12237_binop_int584_result\ := eclat_add(\$12237_binop_int584_arg\(32 to 47) & X"000" & X"1") & \$14086_res\ & eclat_true & eclat_sub(\$12237_binop_int584_arg\(80 to 95) & X"000" & X"1") & \$12237_binop_int584_arg\(96 to 151) & \$12237_binop_int584_arg\(152 to 153);
                          result5714 := \$12237_binop_int584_result\;
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        else
                          \$14105_modulo609_arg\ := eclat_sub(\$14105_modulo609_arg\(0 to 30) & \$14105_modulo609_arg\(31 to 61)) & \$14105_modulo609_arg\(31 to 61);
                          state_var6675 <= \$14105_modulo609\;
                        end if;
                      when \$14274_wait603\ =>
                        \$v5883\ := eclat_not(rdy5722);
                        if \$v5883\(0) = '1' then
                          \$14302\ := \$14274_wait603_arg\(1 to 32) & \$14274_wait603_arg\(33 to 64) & X"0" & X"fa0" & X"0" & X"fa0" & X"0" & X"fa0" & eclat_add(X"0" & X"fa0" & X"1770") & eclat_false;
                        end if;
                        case state_var6676 is
                        when compute5723 =>
                          rdy5722 := eclat_false;
                          case state_var6677 is
                          when \$14343_copy_root_in_ram604\ =>
                            \$v5766\ := eclat_ge(\$14343_copy_root_in_ram604_arg\(0 to 15) & \$14343_copy_root_in_ram604_arg\(16 to 31));
                            if \$v5766\(0) = '1' then
                              \$14343_copy_root_in_ram604_result\ := \$14343_copy_root_in_ram604_arg\(32 to 47);
                              case \$14343_copy_root_in_ram604_id\ is
                              when "000000000110" =>
                                \$14346_next\ := \$14343_copy_root_in_ram604_result\;
                                eclat_print_string(of_string("======================================="));
                                
                                eclat_print_newline(eclat_unit);
                                
                                \$14350_aux605_arg\ := \$14302\(112 to 127) & \$14346_next\ & \$14302\(96 to 111) & \$14302\(112 to 127);
                                state_var6677 <= \$14350_aux605\;
                              when "000000000111" =>
                                \$14344_next\ := \$14343_copy_root_in_ram604_result\;
                                \$v5816\ := \$global_end_ptr_take\;
                                if \$v5816\(0) = '1' then
                                  state_var6677 <= q_wait5815;
                                else
                                  \$global_end_ptr_take\(0) := '1';
                                  \$global_end_ptr\ <= 0;
                                  state_var6677 <= pause_getI5813;
                                end if;
                              when others =>
                                
                              end case;
                            else
                              eclat_print_string(of_string("racine:"));
                              
                              eclat_print_int(\$14343_copy_root_in_ram604_arg\(0 to 15));
                              
                              eclat_print_newline(eclat_unit);
                              
                              \$v5765\ := \$ram_ptr_take\;
                              if \$v5765\(0) = '1' then
                                state_var6677 <= q_wait5764;
                              else
                                \$ram_ptr_take\(0) := '1';
                                \$ram_ptr\ <= to_integer(unsigned(\$14343_copy_root_in_ram604_arg\(0 to 15)));
                                state_var6677 <= pause_getI5762;
                              end if;
                            end if;
                          when \$14350_aux605\ =>
                            eclat_print_string(of_string("     scan="));
                            
                            eclat_print_int(\$14350_aux605_arg\(0 to 15));
                            
                            eclat_print_string(of_string(" | next="));
                            
                            eclat_print_int(\$14350_aux605_arg\(16 to 31));
                            
                            eclat_print_newline(eclat_unit);
                            
                            \$v5811\ := eclat_ge(\$14350_aux605_arg\(0 to 15) & \$14350_aux605_arg\(16 to 31));
                            if \$v5811\(0) = '1' then
                              \$14350_aux605_result\ := \$14350_aux605_arg\(16 to 31);
                              \$14351_next\ := \$14350_aux605_result\;
                              eclat_print_string(of_string("memory copied in to_space : "));
                              
                              eclat_print_int(eclat_sub(\$14351_next\ & \$14302\(112 to 127)));
                              
                              eclat_print_string(of_string(" words"));
                              
                              eclat_print_newline(eclat_unit);
                              
                              \$v5812\ := eclat_gt(eclat_sub(\$14351_next\ & \$14302\(112 to 127)) & X"1770");
                              if \$v5812\(0) = '1' then
                                eclat_print_string(of_string("fatal error: "));
                                
                                eclat_print_string(of_string("Out of memory"));
                                
                                eclat_print_newline(eclat_unit);
                                
                                state_var6677 <= \$14360_forever611\;
                              else
                                \$14329\ := \$14323\(0 to 31) & \$14340\(0 to 31) & \$14351_next\;
                                eclat_print_newline(eclat_unit);
                                
                                eclat_print_newline(eclat_unit);
                                
                                eclat_print_string(of_string("[================= GC END ======================]"));
                                
                                eclat_print_newline(eclat_unit);
                                
                                eclat_print_newline(eclat_unit);
                                
                                result5724 := \$14329\(0 to 31) & \$14329\(32 to 63) & \$14329\(64 to 79) & eclat_add(\$14329\(64 to 79) & \$14274_wait603_arg\(81 to 96)) & \$14302\(112 to 127) & \$14302\(96 to 111);
                                rdy5725 := eclat_true;
                                state_var6677 <= compute5726;
                              end if;
                            else
                              \$v5810\ := \$ram_ptr_take\;
                              if \$v5810\(0) = '1' then
                                state_var6677 <= q_wait5809;
                              else
                                \$ram_ptr_take\(0) := '1';
                                \$ram_ptr\ <= to_integer(unsigned(\$14350_aux605_arg\(0 to 15)));
                                state_var6677 <= pause_getI5807;
                              end if;
                            end if;
                          when \$14360_forever611\ =>
                            state_var6677 <= \$14360_forever611\;
                          when \$14386_loop606\ =>
                            \$v5806\ := eclat_ge(\$14386_loop606_arg\(0 to 15) & eclat_add(\$14386_loop606_arg\(80 to 95) & X"000" & X"1"));
                            if \$v5806\(0) = '1' then
                              \$14386_loop606_result\ := \$14386_loop606_arg\(16 to 31);
                              \$14387_next\ := \$14386_loop606_result\;
                              \$14350_aux605_arg\ := eclat_add(\$14350_aux605_arg\(0 to 15) & eclat_add(eclat_resize(eclat_lsr(eclat_resize(eclat_resize(\$14382\(0 to 30),16),31) & "000"& X"000000" & X"2"),16) & X"000" & X"1")) & \$14387_next\ & \$14350_aux605_arg\(32 to 47) & \$14350_aux605_arg\(48 to 63);
                              state_var6677 <= \$14350_aux605\;
                            else
                              \$v5805\ := \$ram_ptr_take\;
                              if \$v5805\(0) = '1' then
                                state_var6677 <= q_wait5804;
                              else
                                \$ram_ptr_take\(0) := '1';
                                \$ram_ptr\ <= to_integer(unsigned(eclat_add(\$14386_loop606_arg\(64 to 79) & \$14386_loop606_arg\(0 to 15))));
                                state_var6677 <= pause_getI5802;
                              end if;
                            end if;
                          when \$14453_loop607\ =>
                            \$v5779\ := eclat_ge(\$14453_loop607_arg\(0 to 15) & eclat_add(\$14453_loop607_arg\(48 to 63) & X"000" & X"1"));
                            if \$v5779\(0) = '1' then
                              \$14453_loop607_result\ := eclat_unit;
                              \$v5787\ := \$ram_ptr_take\;
                              if \$v5787\(0) = '1' then
                                state_var6677 <= q_wait5786;
                              else
                                \$ram_ptr_take\(0) := '1';
                                \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$14418\(0 to 30),16)));
                                \$ram_write_request\ <= '1';
                                \$ram_write\ <= eclat_resize(\$14386_loop606_arg\(16 to 31),31) & eclat_false;
                                state_var6677 <= pause_setI5784;
                              end if;
                            else
                              \$v5778\ := \$ram_ptr_take\;
                              if \$v5778\(0) = '1' then
                                state_var6677 <= q_wait5777;
                              else
                                \$ram_ptr_take\(0) := '1';
                                \$ram_ptr\ <= to_integer(unsigned(eclat_add(\$14453_loop607_arg\(32 to 47) & \$14453_loop607_arg\(0 to 15))));
                                state_var6677 <= pause_getI5775;
                              end if;
                            end if;
                          when \$14580_loop607\ =>
                            \$v5739\ := eclat_ge(\$14580_loop607_arg\(0 to 15) & eclat_add(\$14580_loop607_arg\(48 to 63) & X"000" & X"1"));
                            if \$v5739\(0) = '1' then
                              \$14580_loop607_result\ := eclat_unit;
                              \$v5747\ := \$ram_ptr_take\;
                              if \$v5747\(0) = '1' then
                                state_var6677 <= q_wait5746;
                              else
                                \$ram_ptr_take\(0) := '1';
                                \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$14543\(0 to 30),16)));
                                \$ram_write_request\ <= '1';
                                \$ram_write\ <= eclat_resize(\$14343_copy_root_in_ram604_arg\(32 to 47),31) & eclat_false;
                                state_var6677 <= pause_setI5744;
                              end if;
                            else
                              \$v5738\ := \$ram_ptr_take\;
                              if \$v5738\(0) = '1' then
                                state_var6677 <= q_wait5737;
                              else
                                \$ram_ptr_take\(0) := '1';
                                \$ram_ptr\ <= to_integer(unsigned(eclat_add(\$14580_loop607_arg\(32 to 47) & \$14580_loop607_arg\(0 to 15))));
                                state_var6677 <= pause_getI5735;
                              end if;
                            end if;
                          when \$14676_loop607\ =>
                            \$v5825\ := eclat_ge(\$14676_loop607_arg\(0 to 15) & eclat_add(\$14676_loop607_arg\(48 to 63) & X"000" & X"1"));
                            if \$v5825\(0) = '1' then
                              \$14676_loop607_result\ := eclat_unit;
                              \$v5833\ := \$ram_ptr_take\;
                              if \$v5833\(0) = '1' then
                                state_var6677 <= q_wait5832;
                              else
                                \$ram_ptr_take\(0) := '1';
                                \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$14274_wait603_arg\(33 to 63),16)));
                                \$ram_write_request\ <= '1';
                                \$ram_write\ <= eclat_resize(\$14323\(32 to 47),31) & eclat_false;
                                state_var6677 <= pause_setI5830;
                              end if;
                            else
                              \$v5824\ := \$ram_ptr_take\;
                              if \$v5824\(0) = '1' then
                                state_var6677 <= q_wait5823;
                              else
                                \$ram_ptr_take\(0) := '1';
                                \$ram_ptr\ <= to_integer(unsigned(eclat_add(\$14676_loop607_arg\(32 to 47) & \$14676_loop607_arg\(0 to 15))));
                                state_var6677 <= pause_getI5821;
                              end if;
                            end if;
                          when \$14772_loop607\ =>
                            \$v5856\ := eclat_ge(\$14772_loop607_arg\(0 to 15) & eclat_add(\$14772_loop607_arg\(48 to 63) & X"000" & X"1"));
                            if \$v5856\(0) = '1' then
                              \$14772_loop607_result\ := eclat_unit;
                              \$v5864\ := \$ram_ptr_take\;
                              if \$v5864\(0) = '1' then
                                state_var6677 <= q_wait5863;
                              else
                                \$ram_ptr_take\(0) := '1';
                                \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$14274_wait603_arg\(1 to 31),16)));
                                \$ram_write_request\ <= '1';
                                \$ram_write\ <= eclat_resize(\$14302\(112 to 127),31) & eclat_false;
                                state_var6677 <= pause_setI5861;
                              end if;
                            else
                              \$v5855\ := \$ram_ptr_take\;
                              if \$v5855\(0) = '1' then
                                state_var6677 <= q_wait5854;
                              else
                                \$ram_ptr_take\(0) := '1';
                                \$ram_ptr\ <= to_integer(unsigned(eclat_add(\$14772_loop607_arg\(32 to 47) & \$14772_loop607_arg\(0 to 15))));
                                state_var6677 <= pause_getI5852;
                              end if;
                            end if;
                          when pause_getI5735 =>
                            state_var6677 <= pause_getII5736;
                          when pause_getI5752 =>
                            state_var6677 <= pause_getII5753;
                          when pause_getI5757 =>
                            state_var6677 <= pause_getII5758;
                          when pause_getI5762 =>
                            state_var6677 <= pause_getII5763;
                          when pause_getI5775 =>
                            state_var6677 <= pause_getII5776;
                          when pause_getI5792 =>
                            state_var6677 <= pause_getII5793;
                          when pause_getI5797 =>
                            state_var6677 <= pause_getII5798;
                          when pause_getI5802 =>
                            state_var6677 <= pause_getII5803;
                          when pause_getI5807 =>
                            state_var6677 <= pause_getII5808;
                          when pause_getI5813 =>
                            state_var6677 <= pause_getII5814;
                          when pause_getI5821 =>
                            state_var6677 <= pause_getII5822;
                          when pause_getI5838 =>
                            state_var6677 <= pause_getII5839;
                          when pause_getI5843 =>
                            state_var6677 <= pause_getII5844;
                          when pause_getI5852 =>
                            state_var6677 <= pause_getII5853;
                          when pause_getI5869 =>
                            state_var6677 <= pause_getII5870;
                          when pause_getI5874 =>
                            state_var6677 <= pause_getII5875;
                          when pause_getII5736 =>
                            \$ram_ptr_take\(0) := '0';
                            \$14614\ := \$ram_value\;
                            \$v5734\ := \$ram_ptr_take\;
                            if \$v5734\(0) = '1' then
                              state_var6677 <= q_wait5733;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(\$14580_loop607_arg\(16 to 31) & \$14580_loop607_arg\(0 to 15))));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$14614\;
                              state_var6677 <= pause_setI5731;
                            end if;
                          when pause_getII5753 =>
                            \$ram_ptr_take\(0) := '0';
                            \$14566_hd\ := \$ram_value\;
                            eclat_print_string(of_string("bloc "));
                            
                            eclat_print_int(eclat_resize(\$14543\(0 to 30),16));
                            
                            eclat_print_string(of_string(" of size "));
                            
                            eclat_print_int(eclat_add(eclat_resize(eclat_lsr(\$14566_hd\(0 to 30) & "000"& X"000000" & X"2"),16) & X"000" & X"1"));
                            
                            eclat_print_string(of_string(" from "));
                            
                            eclat_print_int(eclat_resize(\$14543\(0 to 30),16));
                            
                            eclat_print_string(of_string(" to "));
                            
                            eclat_print_int(\$14343_copy_root_in_ram604_arg\(32 to 47));
                            
                            eclat_print_newline(eclat_unit);
                            
                            \$v5751\ := \$ram_ptr_take\;
                            if \$v5751\(0) = '1' then
                              state_var6677 <= q_wait5750;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(\$14343_copy_root_in_ram604_arg\(32 to 47)));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$14566_hd\;
                              state_var6677 <= pause_setI5748;
                            end if;
                          when pause_getII5758 =>
                            \$ram_ptr_take\(0) := '0';
                            \$14561_w\ := \$ram_value\;
                            \$v5756\ := eclat_if(eclat_not(""&\$14561_w\(31)) & 
                                        eclat_if(eclat_le(\$14343_copy_root_in_ram604_arg\(64 to 79) & eclat_resize(\$14561_w\(0 to 30),16)) & eclat_lt(eclat_resize(\$14561_w\(0 to 30),16) & eclat_add(\$14343_copy_root_in_ram604_arg\(64 to 79) & X"1770")) & eclat_false) & eclat_false);
                            if \$v5756\(0) = '1' then
                              \$14547\ := \$14561_w\ & \$14343_copy_root_in_ram604_arg\(32 to 47);
                              \$v5730\ := \$ram_ptr_take\;
                              if \$v5730\(0) = '1' then
                                state_var6677 <= q_wait5729;
                              else
                                \$ram_ptr_take\(0) := '1';
                                \$ram_ptr_write\ <= to_integer(unsigned(\$14343_copy_root_in_ram604_arg\(0 to 15)));
                                \$ram_write_request\ <= '1';
                                \$ram_write\ <= \$14547\(0 to 31);
                                state_var6677 <= pause_setI5727;
                              end if;
                            else
                              \$v5755\ := \$ram_ptr_take\;
                              if \$v5755\(0) = '1' then
                                state_var6677 <= q_wait5754;
                              else
                                \$ram_ptr_take\(0) := '1';
                                \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$14543\(0 to 30),16)));
                                state_var6677 <= pause_getI5752;
                              end if;
                            end if;
                          when pause_getII5763 =>
                            \$ram_ptr_take\(0) := '0';
                            \$14543\ := \$ram_value\;
                            \$v5761\ := eclat_not(eclat_if(eclat_not(""&\$14543\(31)) & 
                                                  eclat_if(eclat_le(\$14343_copy_root_in_ram604_arg\(48 to 63) & eclat_resize(\$14543\(0 to 30),16)) & eclat_lt(eclat_resize(\$14543\(0 to 30),16) & eclat_add(\$14343_copy_root_in_ram604_arg\(48 to 63) & X"1770")) & eclat_false) & eclat_false));
                            if \$v5761\(0) = '1' then
                              \$14547\ := \$14543\ & \$14343_copy_root_in_ram604_arg\(32 to 47);
                              \$v5730\ := \$ram_ptr_take\;
                              if \$v5730\(0) = '1' then
                                state_var6677 <= q_wait5729;
                              else
                                \$ram_ptr_take\(0) := '1';
                                \$ram_ptr_write\ <= to_integer(unsigned(\$14343_copy_root_in_ram604_arg\(0 to 15)));
                                \$ram_write_request\ <= '1';
                                \$ram_write\ <= \$14547\(0 to 31);
                                state_var6677 <= pause_setI5727;
                              end if;
                            else
                              \$v5760\ := \$ram_ptr_take\;
                              if \$v5760\(0) = '1' then
                                state_var6677 <= q_wait5759;
                              else
                                \$ram_ptr_take\(0) := '1';
                                \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_resize(\$14543\(0 to 30),16) & X"000" & X"1")));
                                state_var6677 <= pause_getI5757;
                              end if;
                            end if;
                          when pause_getII5776 =>
                            \$ram_ptr_take\(0) := '0';
                            \$14487\ := \$ram_value\;
                            \$v5774\ := \$ram_ptr_take\;
                            if \$v5774\(0) = '1' then
                              state_var6677 <= q_wait5773;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(\$14453_loop607_arg\(16 to 31) & \$14453_loop607_arg\(0 to 15))));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$14487\;
                              state_var6677 <= pause_setI5771;
                            end if;
                          when pause_getII5793 =>
                            \$ram_ptr_take\(0) := '0';
                            \$14439_hd\ := \$ram_value\;
                            eclat_print_string(of_string("bloc "));
                            
                            eclat_print_int(eclat_resize(\$14418\(0 to 30),16));
                            
                            eclat_print_string(of_string(" of size "));
                            
                            eclat_print_int(eclat_add(eclat_resize(eclat_lsr(\$14439_hd\(0 to 30) & "000"& X"000000" & X"2"),16) & X"000" & X"1"));
                            
                            eclat_print_string(of_string(" from "));
                            
                            eclat_print_int(eclat_resize(\$14418\(0 to 30),16));
                            
                            eclat_print_string(of_string(" to "));
                            
                            eclat_print_int(\$14386_loop606_arg\(16 to 31));
                            
                            eclat_print_newline(eclat_unit);
                            
                            \$v5791\ := \$ram_ptr_take\;
                            if \$v5791\(0) = '1' then
                              state_var6677 <= q_wait5790;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(\$14386_loop606_arg\(16 to 31)));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$14439_hd\;
                              state_var6677 <= pause_setI5788;
                            end if;
                          when pause_getII5798 =>
                            \$ram_ptr_take\(0) := '0';
                            \$14434_w\ := \$ram_value\;
                            \$v5796\ := eclat_if(eclat_not(""&\$14434_w\(31)) & 
                                        eclat_if(eclat_le(\$14386_loop606_arg\(48 to 63) & eclat_resize(\$14434_w\(0 to 30),16)) & eclat_lt(eclat_resize(\$14434_w\(0 to 30),16) & eclat_add(\$14386_loop606_arg\(48 to 63) & X"1770")) & eclat_false) & eclat_false);
                            if \$v5796\(0) = '1' then
                              \$14422\ := \$14434_w\ & \$14386_loop606_arg\(16 to 31);
                              \$v5770\ := \$ram_ptr_take\;
                              if \$v5770\(0) = '1' then
                                state_var6677 <= q_wait5769;
                              else
                                \$ram_ptr_take\(0) := '1';
                                \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(\$14386_loop606_arg\(64 to 79) & \$14386_loop606_arg\(0 to 15))));
                                \$ram_write_request\ <= '1';
                                \$ram_write\ <= \$14422\(0 to 31);
                                state_var6677 <= pause_setI5767;
                              end if;
                            else
                              \$v5795\ := \$ram_ptr_take\;
                              if \$v5795\(0) = '1' then
                                state_var6677 <= q_wait5794;
                              else
                                \$ram_ptr_take\(0) := '1';
                                \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$14418\(0 to 30),16)));
                                state_var6677 <= pause_getI5792;
                              end if;
                            end if;
                          when pause_getII5803 =>
                            \$ram_ptr_take\(0) := '0';
                            \$14418\ := \$ram_value\;
                            \$v5801\ := eclat_not(eclat_if(eclat_not(""&\$14418\(31)) & 
                                                  eclat_if(eclat_le(\$14386_loop606_arg\(32 to 47) & eclat_resize(\$14418\(0 to 30),16)) & eclat_lt(eclat_resize(\$14418\(0 to 30),16) & eclat_add(\$14386_loop606_arg\(32 to 47) & X"1770")) & eclat_false) & eclat_false));
                            if \$v5801\(0) = '1' then
                              \$14422\ := \$14418\ & \$14386_loop606_arg\(16 to 31);
                              \$v5770\ := \$ram_ptr_take\;
                              if \$v5770\(0) = '1' then
                                state_var6677 <= q_wait5769;
                              else
                                \$ram_ptr_take\(0) := '1';
                                \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(\$14386_loop606_arg\(64 to 79) & \$14386_loop606_arg\(0 to 15))));
                                \$ram_write_request\ <= '1';
                                \$ram_write\ <= \$14422\(0 to 31);
                                state_var6677 <= pause_setI5767;
                              end if;
                            else
                              \$v5800\ := \$ram_ptr_take\;
                              if \$v5800\(0) = '1' then
                                state_var6677 <= q_wait5799;
                              else
                                \$ram_ptr_take\(0) := '1';
                                \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_resize(\$14418\(0 to 30),16) & X"000" & X"1")));
                                state_var6677 <= pause_getI5797;
                              end if;
                            end if;
                          when pause_getII5808 =>
                            \$ram_ptr_take\(0) := '0';
                            \$14382\ := \$ram_value\;
                            \$14386_loop606_arg\ := X"000" & X"1" & \$14350_aux605_arg\(16 to 31) & \$14350_aux605_arg\(32 to 47) & \$14350_aux605_arg\(48 to 63) & \$14350_aux605_arg\(0 to 15) & eclat_resize(eclat_lsr(eclat_resize(eclat_resize(\$14382\(0 to 30),16),31) & "000"& X"000000" & X"2"),16);
                            state_var6677 <= \$14386_loop606\;
                          when pause_getII5814 =>
                            \$global_end_ptr_take\(0) := '0';
                            \$14345\ := \$global_end_value\;
                            \$14343_copy_root_in_ram604_id\ := "000000000110";
                            \$14343_copy_root_in_ram604_arg\ := X"3e80" & \$14345\ & \$14344_next\ & \$14302\(96 to 111) & \$14302\(112 to 127);
                            state_var6677 <= \$14343_copy_root_in_ram604\;
                          when pause_getII5822 =>
                            \$ram_ptr_take\(0) := '0';
                            \$14710\ := \$ram_value\;
                            \$v5820\ := \$ram_ptr_take\;
                            if \$v5820\(0) = '1' then
                              state_var6677 <= q_wait5819;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(\$14676_loop607_arg\(16 to 31) & \$14676_loop607_arg\(0 to 15))));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$14710\;
                              state_var6677 <= pause_setI5817;
                            end if;
                          when pause_getII5839 =>
                            \$ram_ptr_take\(0) := '0';
                            \$14662_hd\ := \$ram_value\;
                            eclat_print_string(of_string("bloc "));
                            
                            eclat_print_int(eclat_resize(\$14274_wait603_arg\(33 to 63),16));
                            
                            eclat_print_string(of_string(" of size "));
                            
                            eclat_print_int(eclat_add(eclat_resize(eclat_lsr(\$14662_hd\(0 to 30) & "000"& X"000000" & X"2"),16) & X"000" & X"1"));
                            
                            eclat_print_string(of_string(" from "));
                            
                            eclat_print_int(eclat_resize(\$14274_wait603_arg\(33 to 63),16));
                            
                            eclat_print_string(of_string(" to "));
                            
                            eclat_print_int(\$14323\(32 to 47));
                            
                            eclat_print_newline(eclat_unit);
                            
                            \$v5837\ := \$ram_ptr_take\;
                            if \$v5837\(0) = '1' then
                              state_var6677 <= q_wait5836;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(\$14323\(32 to 47)));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$14662_hd\;
                              state_var6677 <= pause_setI5834;
                            end if;
                          when pause_getII5844 =>
                            \$ram_ptr_take\(0) := '0';
                            \$14657_w\ := \$ram_value\;
                            \$v5842\ := eclat_if(eclat_not(""&\$14657_w\(31)) & 
                                        eclat_if(eclat_le(\$14302\(112 to 127) & eclat_resize(\$14657_w\(0 to 30),16)) & eclat_lt(eclat_resize(\$14657_w\(0 to 30),16) & eclat_add(\$14302\(112 to 127) & X"1770")) & eclat_false) & eclat_false);
                            if \$v5842\(0) = '1' then
                              \$14340\ := \$14657_w\ & \$14323\(32 to 47);
                              \$14343_copy_root_in_ram604_id\ := "000000000111";
                              \$14343_copy_root_in_ram604_arg\ := X"0" & X"3e8" & \$14274_wait603_arg\(65 to 80) & \$14340\(32 to 47) & \$14302\(96 to 111) & \$14302\(112 to 127);
                              state_var6677 <= \$14343_copy_root_in_ram604\;
                            else
                              \$v5841\ := \$ram_ptr_take\;
                              if \$v5841\(0) = '1' then
                                state_var6677 <= q_wait5840;
                              else
                                \$ram_ptr_take\(0) := '1';
                                \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$14274_wait603_arg\(33 to 63),16)));
                                state_var6677 <= pause_getI5838;
                              end if;
                            end if;
                          when pause_getII5853 =>
                            \$ram_ptr_take\(0) := '0';
                            \$14806\ := \$ram_value\;
                            \$v5851\ := \$ram_ptr_take\;
                            if \$v5851\(0) = '1' then
                              state_var6677 <= q_wait5850;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(\$14772_loop607_arg\(16 to 31) & \$14772_loop607_arg\(0 to 15))));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$14806\;
                              state_var6677 <= pause_setI5848;
                            end if;
                          when pause_getII5870 =>
                            \$ram_ptr_take\(0) := '0';
                            \$14758_hd\ := \$ram_value\;
                            eclat_print_string(of_string("bloc "));
                            
                            eclat_print_int(eclat_resize(\$14274_wait603_arg\(1 to 31),16));
                            
                            eclat_print_string(of_string(" of size "));
                            
                            eclat_print_int(eclat_add(eclat_resize(eclat_lsr(\$14758_hd\(0 to 30) & "000"& X"000000" & X"2"),16) & X"000" & X"1"));
                            
                            eclat_print_string(of_string(" from "));
                            
                            eclat_print_int(eclat_resize(\$14274_wait603_arg\(1 to 31),16));
                            
                            eclat_print_string(of_string(" to "));
                            
                            eclat_print_int(\$14302\(112 to 127));
                            
                            eclat_print_newline(eclat_unit);
                            
                            \$v5868\ := \$ram_ptr_take\;
                            if \$v5868\(0) = '1' then
                              state_var6677 <= q_wait5867;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(\$14302\(112 to 127)));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$14758_hd\;
                              state_var6677 <= pause_setI5865;
                            end if;
                          when pause_getII5875 =>
                            \$ram_ptr_take\(0) := '0';
                            \$14753_w\ := \$ram_value\;
                            \$v5873\ := eclat_if(eclat_not(""&\$14753_w\(31)) & 
                                        eclat_if(eclat_le(\$14302\(112 to 127) & eclat_resize(\$14753_w\(0 to 30),16)) & eclat_lt(eclat_resize(\$14753_w\(0 to 30),16) & eclat_add(\$14302\(112 to 127) & X"1770")) & eclat_false) & eclat_false);
                            if \$v5873\(0) = '1' then
                              \$14323\ := \$14753_w\ & \$14302\(112 to 127);
                              \$v5847\ := eclat_not(eclat_if(eclat_not(""&\$14274_wait603_arg\(64)) & 
                                                    eclat_if(eclat_le(\$14302\(96 to 111) & eclat_resize(\$14274_wait603_arg\(33 to 63),16)) & eclat_lt(eclat_resize(\$14274_wait603_arg\(33 to 63),16) & eclat_add(\$14302\(96 to 111) & X"1770")) & eclat_false) & eclat_false));
                              if \$v5847\(0) = '1' then
                                \$14340\ := \$14274_wait603_arg\(33 to 64) & \$14323\(32 to 47);
                                \$14343_copy_root_in_ram604_id\ := "000000000111";
                                \$14343_copy_root_in_ram604_arg\ := X"0" & X"3e8" & \$14274_wait603_arg\(65 to 80) & \$14340\(32 to 47) & \$14302\(96 to 111) & \$14302\(112 to 127);
                                state_var6677 <= \$14343_copy_root_in_ram604\;
                              else
                                \$v5846\ := \$ram_ptr_take\;
                                if \$v5846\(0) = '1' then
                                  state_var6677 <= q_wait5845;
                                else
                                  \$ram_ptr_take\(0) := '1';
                                  \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_resize(\$14274_wait603_arg\(33 to 63),16) & X"000" & X"1")));
                                  state_var6677 <= pause_getI5843;
                                end if;
                              end if;
                            else
                              \$v5872\ := \$ram_ptr_take\;
                              if \$v5872\(0) = '1' then
                                state_var6677 <= q_wait5871;
                              else
                                \$ram_ptr_take\(0) := '1';
                                \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$14274_wait603_arg\(1 to 31),16)));
                                state_var6677 <= pause_getI5869;
                              end if;
                            end if;
                          when pause_setI5727 =>
                            \$ram_write_request\ <= '0';
                            state_var6677 <= pause_setII5728;
                          when pause_setI5731 =>
                            \$ram_write_request\ <= '0';
                            state_var6677 <= pause_setII5732;
                          when pause_setI5740 =>
                            \$ram_write_request\ <= '0';
                            state_var6677 <= pause_setII5741;
                          when pause_setI5744 =>
                            \$ram_write_request\ <= '0';
                            state_var6677 <= pause_setII5745;
                          when pause_setI5748 =>
                            \$ram_write_request\ <= '0';
                            state_var6677 <= pause_setII5749;
                          when pause_setI5767 =>
                            \$ram_write_request\ <= '0';
                            state_var6677 <= pause_setII5768;
                          when pause_setI5771 =>
                            \$ram_write_request\ <= '0';
                            state_var6677 <= pause_setII5772;
                          when pause_setI5780 =>
                            \$ram_write_request\ <= '0';
                            state_var6677 <= pause_setII5781;
                          when pause_setI5784 =>
                            \$ram_write_request\ <= '0';
                            state_var6677 <= pause_setII5785;
                          when pause_setI5788 =>
                            \$ram_write_request\ <= '0';
                            state_var6677 <= pause_setII5789;
                          when pause_setI5817 =>
                            \$ram_write_request\ <= '0';
                            state_var6677 <= pause_setII5818;
                          when pause_setI5826 =>
                            \$ram_write_request\ <= '0';
                            state_var6677 <= pause_setII5827;
                          when pause_setI5830 =>
                            \$ram_write_request\ <= '0';
                            state_var6677 <= pause_setII5831;
                          when pause_setI5834 =>
                            \$ram_write_request\ <= '0';
                            state_var6677 <= pause_setII5835;
                          when pause_setI5848 =>
                            \$ram_write_request\ <= '0';
                            state_var6677 <= pause_setII5849;
                          when pause_setI5857 =>
                            \$ram_write_request\ <= '0';
                            state_var6677 <= pause_setII5858;
                          when pause_setI5861 =>
                            \$ram_write_request\ <= '0';
                            state_var6677 <= pause_setII5862;
                          when pause_setI5865 =>
                            \$ram_write_request\ <= '0';
                            state_var6677 <= pause_setII5866;
                          when pause_setII5728 =>
                            \$ram_ptr_take\(0) := '0';
                            eclat_print_string(of_string(" next="));
                            
                            eclat_print_int(\$14547\(32 to 47));
                            
                            eclat_print_newline(eclat_unit);
                            
                            \$14343_copy_root_in_ram604_arg\ := eclat_add(\$14343_copy_root_in_ram604_arg\(0 to 15) & X"000" & X"1") & \$14343_copy_root_in_ram604_arg\(16 to 31) & \$14547\(32 to 47) & \$14343_copy_root_in_ram604_arg\(48 to 63) & \$14343_copy_root_in_ram604_arg\(64 to 79);
                            state_var6677 <= \$14343_copy_root_in_ram604\;
                          when pause_setII5732 =>
                            \$ram_ptr_take\(0) := '0';
                            \$14580_loop607_arg\ := eclat_add(\$14580_loop607_arg\(0 to 15) & X"000" & X"1") & \$14580_loop607_arg\(16 to 31) & \$14580_loop607_arg\(32 to 47) & \$14580_loop607_arg\(48 to 63);
                            state_var6677 <= \$14580_loop607\;
                          when pause_setII5741 =>
                            \$ram_ptr_take\(0) := '0';
                            \$14547\ := eclat_resize(\$14343_copy_root_in_ram604_arg\(32 to 47),31) & eclat_false & eclat_add(\$14343_copy_root_in_ram604_arg\(32 to 47) & eclat_add(eclat_resize(eclat_lsr(\$14566_hd\(0 to 30) & "000"& X"000000" & X"2"),16) & X"000" & X"1"));
                            \$v5730\ := \$ram_ptr_take\;
                            if \$v5730\(0) = '1' then
                              state_var6677 <= q_wait5729;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(\$14343_copy_root_in_ram604_arg\(0 to 15)));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$14547\(0 to 31);
                              state_var6677 <= pause_setI5727;
                            end if;
                          when pause_setII5745 =>
                            \$ram_ptr_take\(0) := '0';
                            \$v5743\ := \$ram_ptr_take\;
                            if \$v5743\(0) = '1' then
                              state_var6677 <= q_wait5742;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_resize(\$14543\(0 to 30),16) & X"000" & X"1")));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= eclat_resize(\$14343_copy_root_in_ram604_arg\(32 to 47),31) & eclat_false;
                              state_var6677 <= pause_setI5740;
                            end if;
                          when pause_setII5749 =>
                            \$ram_ptr_take\(0) := '0';
                            \$14580_loop607_arg\ := X"000" & X"1" & \$14343_copy_root_in_ram604_arg\(32 to 47) & eclat_resize(\$14543\(0 to 30),16) & eclat_resize(eclat_lsr(\$14566_hd\(0 to 30) & "000"& X"000000" & X"2"),16);
                            state_var6677 <= \$14580_loop607\;
                          when pause_setII5768 =>
                            \$ram_ptr_take\(0) := '0';
                            \$14386_loop606_arg\ := eclat_add(\$14386_loop606_arg\(0 to 15) & X"000" & X"1") & \$14422\(32 to 47) & \$14386_loop606_arg\(32 to 47) & \$14386_loop606_arg\(48 to 63) & \$14386_loop606_arg\(64 to 79) & \$14386_loop606_arg\(80 to 95);
                            state_var6677 <= \$14386_loop606\;
                          when pause_setII5772 =>
                            \$ram_ptr_take\(0) := '0';
                            \$14453_loop607_arg\ := eclat_add(\$14453_loop607_arg\(0 to 15) & X"000" & X"1") & \$14453_loop607_arg\(16 to 31) & \$14453_loop607_arg\(32 to 47) & \$14453_loop607_arg\(48 to 63);
                            state_var6677 <= \$14453_loop607\;
                          when pause_setII5781 =>
                            \$ram_ptr_take\(0) := '0';
                            \$14422\ := eclat_resize(\$14386_loop606_arg\(16 to 31),31) & eclat_false & eclat_add(\$14386_loop606_arg\(16 to 31) & eclat_add(eclat_resize(eclat_lsr(\$14439_hd\(0 to 30) & "000"& X"000000" & X"2"),16) & X"000" & X"1"));
                            \$v5770\ := \$ram_ptr_take\;
                            if \$v5770\(0) = '1' then
                              state_var6677 <= q_wait5769;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(\$14386_loop606_arg\(64 to 79) & \$14386_loop606_arg\(0 to 15))));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$14422\(0 to 31);
                              state_var6677 <= pause_setI5767;
                            end if;
                          when pause_setII5785 =>
                            \$ram_ptr_take\(0) := '0';
                            \$v5783\ := \$ram_ptr_take\;
                            if \$v5783\(0) = '1' then
                              state_var6677 <= q_wait5782;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_resize(\$14418\(0 to 30),16) & X"000" & X"1")));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= eclat_resize(\$14386_loop606_arg\(16 to 31),31) & eclat_false;
                              state_var6677 <= pause_setI5780;
                            end if;
                          when pause_setII5789 =>
                            \$ram_ptr_take\(0) := '0';
                            \$14453_loop607_arg\ := X"000" & X"1" & \$14386_loop606_arg\(16 to 31) & eclat_resize(\$14418\(0 to 30),16) & eclat_resize(eclat_lsr(\$14439_hd\(0 to 30) & "000"& X"000000" & X"2"),16);
                            state_var6677 <= \$14453_loop607\;
                          when pause_setII5818 =>
                            \$ram_ptr_take\(0) := '0';
                            \$14676_loop607_arg\ := eclat_add(\$14676_loop607_arg\(0 to 15) & X"000" & X"1") & \$14676_loop607_arg\(16 to 31) & \$14676_loop607_arg\(32 to 47) & \$14676_loop607_arg\(48 to 63);
                            state_var6677 <= \$14676_loop607\;
                          when pause_setII5827 =>
                            \$ram_ptr_take\(0) := '0';
                            \$14340\ := eclat_resize(\$14323\(32 to 47),31) & eclat_false & eclat_add(\$14323\(32 to 47) & eclat_add(eclat_resize(eclat_lsr(\$14662_hd\(0 to 30) & "000"& X"000000" & X"2"),16) & X"000" & X"1"));
                            \$14343_copy_root_in_ram604_id\ := "000000000111";
                            \$14343_copy_root_in_ram604_arg\ := X"0" & X"3e8" & \$14274_wait603_arg\(65 to 80) & \$14340\(32 to 47) & \$14302\(96 to 111) & \$14302\(112 to 127);
                            state_var6677 <= \$14343_copy_root_in_ram604\;
                          when pause_setII5831 =>
                            \$ram_ptr_take\(0) := '0';
                            \$v5829\ := \$ram_ptr_take\;
                            if \$v5829\(0) = '1' then
                              state_var6677 <= q_wait5828;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_resize(\$14274_wait603_arg\(33 to 63),16) & X"000" & X"1")));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= eclat_resize(\$14323\(32 to 47),31) & eclat_false;
                              state_var6677 <= pause_setI5826;
                            end if;
                          when pause_setII5835 =>
                            \$ram_ptr_take\(0) := '0';
                            \$14676_loop607_arg\ := X"000" & X"1" & \$14323\(32 to 47) & eclat_resize(\$14274_wait603_arg\(33 to 63),16) & eclat_resize(eclat_lsr(\$14662_hd\(0 to 30) & "000"& X"000000" & X"2"),16);
                            state_var6677 <= \$14676_loop607\;
                          when pause_setII5849 =>
                            \$ram_ptr_take\(0) := '0';
                            \$14772_loop607_arg\ := eclat_add(\$14772_loop607_arg\(0 to 15) & X"000" & X"1") & \$14772_loop607_arg\(16 to 31) & \$14772_loop607_arg\(32 to 47) & \$14772_loop607_arg\(48 to 63);
                            state_var6677 <= \$14772_loop607\;
                          when pause_setII5858 =>
                            \$ram_ptr_take\(0) := '0';
                            \$14323\ := eclat_resize(\$14302\(112 to 127),31) & eclat_false & eclat_add(\$14302\(112 to 127) & eclat_add(eclat_resize(eclat_lsr(\$14758_hd\(0 to 30) & "000"& X"000000" & X"2"),16) & X"000" & X"1"));
                            \$v5847\ := eclat_not(eclat_if(eclat_not(""&\$14274_wait603_arg\(64)) & 
                                                  eclat_if(eclat_le(\$14302\(96 to 111) & eclat_resize(\$14274_wait603_arg\(33 to 63),16)) & eclat_lt(eclat_resize(\$14274_wait603_arg\(33 to 63),16) & eclat_add(\$14302\(96 to 111) & X"1770")) & eclat_false) & eclat_false));
                            if \$v5847\(0) = '1' then
                              \$14340\ := \$14274_wait603_arg\(33 to 64) & \$14323\(32 to 47);
                              \$14343_copy_root_in_ram604_id\ := "000000000111";
                              \$14343_copy_root_in_ram604_arg\ := X"0" & X"3e8" & \$14274_wait603_arg\(65 to 80) & \$14340\(32 to 47) & \$14302\(96 to 111) & \$14302\(112 to 127);
                              state_var6677 <= \$14343_copy_root_in_ram604\;
                            else
                              \$v5846\ := \$ram_ptr_take\;
                              if \$v5846\(0) = '1' then
                                state_var6677 <= q_wait5845;
                              else
                                \$ram_ptr_take\(0) := '1';
                                \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_resize(\$14274_wait603_arg\(33 to 63),16) & X"000" & X"1")));
                                state_var6677 <= pause_getI5843;
                              end if;
                            end if;
                          when pause_setII5862 =>
                            \$ram_ptr_take\(0) := '0';
                            \$v5860\ := \$ram_ptr_take\;
                            if \$v5860\(0) = '1' then
                              state_var6677 <= q_wait5859;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_resize(\$14274_wait603_arg\(1 to 31),16) & X"000" & X"1")));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= eclat_resize(\$14302\(112 to 127),31) & eclat_false;
                              state_var6677 <= pause_setI5857;
                            end if;
                          when pause_setII5866 =>
                            \$ram_ptr_take\(0) := '0';
                            \$14772_loop607_arg\ := X"000" & X"1" & \$14302\(112 to 127) & eclat_resize(\$14274_wait603_arg\(1 to 31),16) & eclat_resize(eclat_lsr(\$14758_hd\(0 to 30) & "000"& X"000000" & X"2"),16);
                            state_var6677 <= \$14772_loop607\;
                          when q_wait5729 =>
                            \$v5730\ := \$ram_ptr_take\;
                            if \$v5730\(0) = '1' then
                              state_var6677 <= q_wait5729;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(\$14343_copy_root_in_ram604_arg\(0 to 15)));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$14547\(0 to 31);
                              state_var6677 <= pause_setI5727;
                            end if;
                          when q_wait5733 =>
                            \$v5734\ := \$ram_ptr_take\;
                            if \$v5734\(0) = '1' then
                              state_var6677 <= q_wait5733;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(\$14580_loop607_arg\(16 to 31) & \$14580_loop607_arg\(0 to 15))));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$14614\;
                              state_var6677 <= pause_setI5731;
                            end if;
                          when q_wait5737 =>
                            \$v5738\ := \$ram_ptr_take\;
                            if \$v5738\(0) = '1' then
                              state_var6677 <= q_wait5737;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr\ <= to_integer(unsigned(eclat_add(\$14580_loop607_arg\(32 to 47) & \$14580_loop607_arg\(0 to 15))));
                              state_var6677 <= pause_getI5735;
                            end if;
                          when q_wait5742 =>
                            \$v5743\ := \$ram_ptr_take\;
                            if \$v5743\(0) = '1' then
                              state_var6677 <= q_wait5742;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_resize(\$14543\(0 to 30),16) & X"000" & X"1")));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= eclat_resize(\$14343_copy_root_in_ram604_arg\(32 to 47),31) & eclat_false;
                              state_var6677 <= pause_setI5740;
                            end if;
                          when q_wait5746 =>
                            \$v5747\ := \$ram_ptr_take\;
                            if \$v5747\(0) = '1' then
                              state_var6677 <= q_wait5746;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$14543\(0 to 30),16)));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= eclat_resize(\$14343_copy_root_in_ram604_arg\(32 to 47),31) & eclat_false;
                              state_var6677 <= pause_setI5744;
                            end if;
                          when q_wait5750 =>
                            \$v5751\ := \$ram_ptr_take\;
                            if \$v5751\(0) = '1' then
                              state_var6677 <= q_wait5750;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(\$14343_copy_root_in_ram604_arg\(32 to 47)));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$14566_hd\;
                              state_var6677 <= pause_setI5748;
                            end if;
                          when q_wait5754 =>
                            \$v5755\ := \$ram_ptr_take\;
                            if \$v5755\(0) = '1' then
                              state_var6677 <= q_wait5754;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$14543\(0 to 30),16)));
                              state_var6677 <= pause_getI5752;
                            end if;
                          when q_wait5759 =>
                            \$v5760\ := \$ram_ptr_take\;
                            if \$v5760\(0) = '1' then
                              state_var6677 <= q_wait5759;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_resize(\$14543\(0 to 30),16) & X"000" & X"1")));
                              state_var6677 <= pause_getI5757;
                            end if;
                          when q_wait5764 =>
                            \$v5765\ := \$ram_ptr_take\;
                            if \$v5765\(0) = '1' then
                              state_var6677 <= q_wait5764;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr\ <= to_integer(unsigned(\$14343_copy_root_in_ram604_arg\(0 to 15)));
                              state_var6677 <= pause_getI5762;
                            end if;
                          when q_wait5769 =>
                            \$v5770\ := \$ram_ptr_take\;
                            if \$v5770\(0) = '1' then
                              state_var6677 <= q_wait5769;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(\$14386_loop606_arg\(64 to 79) & \$14386_loop606_arg\(0 to 15))));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$14422\(0 to 31);
                              state_var6677 <= pause_setI5767;
                            end if;
                          when q_wait5773 =>
                            \$v5774\ := \$ram_ptr_take\;
                            if \$v5774\(0) = '1' then
                              state_var6677 <= q_wait5773;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(\$14453_loop607_arg\(16 to 31) & \$14453_loop607_arg\(0 to 15))));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$14487\;
                              state_var6677 <= pause_setI5771;
                            end if;
                          when q_wait5777 =>
                            \$v5778\ := \$ram_ptr_take\;
                            if \$v5778\(0) = '1' then
                              state_var6677 <= q_wait5777;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr\ <= to_integer(unsigned(eclat_add(\$14453_loop607_arg\(32 to 47) & \$14453_loop607_arg\(0 to 15))));
                              state_var6677 <= pause_getI5775;
                            end if;
                          when q_wait5782 =>
                            \$v5783\ := \$ram_ptr_take\;
                            if \$v5783\(0) = '1' then
                              state_var6677 <= q_wait5782;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_resize(\$14418\(0 to 30),16) & X"000" & X"1")));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= eclat_resize(\$14386_loop606_arg\(16 to 31),31) & eclat_false;
                              state_var6677 <= pause_setI5780;
                            end if;
                          when q_wait5786 =>
                            \$v5787\ := \$ram_ptr_take\;
                            if \$v5787\(0) = '1' then
                              state_var6677 <= q_wait5786;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$14418\(0 to 30),16)));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= eclat_resize(\$14386_loop606_arg\(16 to 31),31) & eclat_false;
                              state_var6677 <= pause_setI5784;
                            end if;
                          when q_wait5790 =>
                            \$v5791\ := \$ram_ptr_take\;
                            if \$v5791\(0) = '1' then
                              state_var6677 <= q_wait5790;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(\$14386_loop606_arg\(16 to 31)));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$14439_hd\;
                              state_var6677 <= pause_setI5788;
                            end if;
                          when q_wait5794 =>
                            \$v5795\ := \$ram_ptr_take\;
                            if \$v5795\(0) = '1' then
                              state_var6677 <= q_wait5794;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$14418\(0 to 30),16)));
                              state_var6677 <= pause_getI5792;
                            end if;
                          when q_wait5799 =>
                            \$v5800\ := \$ram_ptr_take\;
                            if \$v5800\(0) = '1' then
                              state_var6677 <= q_wait5799;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_resize(\$14418\(0 to 30),16) & X"000" & X"1")));
                              state_var6677 <= pause_getI5797;
                            end if;
                          when q_wait5804 =>
                            \$v5805\ := \$ram_ptr_take\;
                            if \$v5805\(0) = '1' then
                              state_var6677 <= q_wait5804;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr\ <= to_integer(unsigned(eclat_add(\$14386_loop606_arg\(64 to 79) & \$14386_loop606_arg\(0 to 15))));
                              state_var6677 <= pause_getI5802;
                            end if;
                          when q_wait5809 =>
                            \$v5810\ := \$ram_ptr_take\;
                            if \$v5810\(0) = '1' then
                              state_var6677 <= q_wait5809;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr\ <= to_integer(unsigned(\$14350_aux605_arg\(0 to 15)));
                              state_var6677 <= pause_getI5807;
                            end if;
                          when q_wait5815 =>
                            \$v5816\ := \$global_end_ptr_take\;
                            if \$v5816\(0) = '1' then
                              state_var6677 <= q_wait5815;
                            else
                              \$global_end_ptr_take\(0) := '1';
                              \$global_end_ptr\ <= 0;
                              state_var6677 <= pause_getI5813;
                            end if;
                          when q_wait5819 =>
                            \$v5820\ := \$ram_ptr_take\;
                            if \$v5820\(0) = '1' then
                              state_var6677 <= q_wait5819;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(\$14676_loop607_arg\(16 to 31) & \$14676_loop607_arg\(0 to 15))));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$14710\;
                              state_var6677 <= pause_setI5817;
                            end if;
                          when q_wait5823 =>
                            \$v5824\ := \$ram_ptr_take\;
                            if \$v5824\(0) = '1' then
                              state_var6677 <= q_wait5823;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr\ <= to_integer(unsigned(eclat_add(\$14676_loop607_arg\(32 to 47) & \$14676_loop607_arg\(0 to 15))));
                              state_var6677 <= pause_getI5821;
                            end if;
                          when q_wait5828 =>
                            \$v5829\ := \$ram_ptr_take\;
                            if \$v5829\(0) = '1' then
                              state_var6677 <= q_wait5828;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_resize(\$14274_wait603_arg\(33 to 63),16) & X"000" & X"1")));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= eclat_resize(\$14323\(32 to 47),31) & eclat_false;
                              state_var6677 <= pause_setI5826;
                            end if;
                          when q_wait5832 =>
                            \$v5833\ := \$ram_ptr_take\;
                            if \$v5833\(0) = '1' then
                              state_var6677 <= q_wait5832;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$14274_wait603_arg\(33 to 63),16)));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= eclat_resize(\$14323\(32 to 47),31) & eclat_false;
                              state_var6677 <= pause_setI5830;
                            end if;
                          when q_wait5836 =>
                            \$v5837\ := \$ram_ptr_take\;
                            if \$v5837\(0) = '1' then
                              state_var6677 <= q_wait5836;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(\$14323\(32 to 47)));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$14662_hd\;
                              state_var6677 <= pause_setI5834;
                            end if;
                          when q_wait5840 =>
                            \$v5841\ := \$ram_ptr_take\;
                            if \$v5841\(0) = '1' then
                              state_var6677 <= q_wait5840;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$14274_wait603_arg\(33 to 63),16)));
                              state_var6677 <= pause_getI5838;
                            end if;
                          when q_wait5845 =>
                            \$v5846\ := \$ram_ptr_take\;
                            if \$v5846\(0) = '1' then
                              state_var6677 <= q_wait5845;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_resize(\$14274_wait603_arg\(33 to 63),16) & X"000" & X"1")));
                              state_var6677 <= pause_getI5843;
                            end if;
                          when q_wait5850 =>
                            \$v5851\ := \$ram_ptr_take\;
                            if \$v5851\(0) = '1' then
                              state_var6677 <= q_wait5850;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(\$14772_loop607_arg\(16 to 31) & \$14772_loop607_arg\(0 to 15))));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$14806\;
                              state_var6677 <= pause_setI5848;
                            end if;
                          when q_wait5854 =>
                            \$v5855\ := \$ram_ptr_take\;
                            if \$v5855\(0) = '1' then
                              state_var6677 <= q_wait5854;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr\ <= to_integer(unsigned(eclat_add(\$14772_loop607_arg\(32 to 47) & \$14772_loop607_arg\(0 to 15))));
                              state_var6677 <= pause_getI5852;
                            end if;
                          when q_wait5859 =>
                            \$v5860\ := \$ram_ptr_take\;
                            if \$v5860\(0) = '1' then
                              state_var6677 <= q_wait5859;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_resize(\$14274_wait603_arg\(1 to 31),16) & X"000" & X"1")));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= eclat_resize(\$14302\(112 to 127),31) & eclat_false;
                              state_var6677 <= pause_setI5857;
                            end if;
                          when q_wait5863 =>
                            \$v5864\ := \$ram_ptr_take\;
                            if \$v5864\(0) = '1' then
                              state_var6677 <= q_wait5863;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$14274_wait603_arg\(1 to 31),16)));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= eclat_resize(\$14302\(112 to 127),31) & eclat_false;
                              state_var6677 <= pause_setI5861;
                            end if;
                          when q_wait5867 =>
                            \$v5868\ := \$ram_ptr_take\;
                            if \$v5868\(0) = '1' then
                              state_var6677 <= q_wait5867;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(\$14302\(112 to 127)));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$14758_hd\;
                              state_var6677 <= pause_setI5865;
                            end if;
                          when q_wait5871 =>
                            \$v5872\ := \$ram_ptr_take\;
                            if \$v5872\(0) = '1' then
                              state_var6677 <= q_wait5871;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$14274_wait603_arg\(1 to 31),16)));
                              state_var6677 <= pause_getI5869;
                            end if;
                          when q_wait5876 =>
                            \$v5877\ := \$ram_ptr_take\;
                            if \$v5877\(0) = '1' then
                              state_var6677 <= q_wait5876;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_resize(\$14274_wait603_arg\(1 to 31),16) & X"000" & X"1")));
                              state_var6677 <= pause_getI5874;
                            end if;
                          when compute5726 =>
                            rdy5725 := eclat_false;
                            \$v5879\ := eclat_gt(eclat_add(\$14302\(80 to 95) & \$14274_wait603_arg\(81 to 96)) & eclat_add(\$14302\(96 to 111) & X"1770"));
                            if \$v5879\(0) = '1' then
                              eclat_print_newline(eclat_unit);
                              
                              eclat_print_newline(eclat_unit);
                              
                              eclat_print_string(of_string("[================= GC START ======================]"));
                              
                              eclat_print_newline(eclat_unit);
                              
                              eclat_print_newline(eclat_unit);
                              
                              \$v5878\ := eclat_not(eclat_if(eclat_not(""&\$14274_wait603_arg\(32)) & 
                                                    eclat_if(eclat_le(\$14302\(96 to 111) & eclat_resize(\$14274_wait603_arg\(1 to 31),16)) & eclat_lt(eclat_resize(\$14274_wait603_arg\(1 to 31),16) & eclat_add(\$14302\(96 to 111) & X"1770")) & eclat_false) & eclat_false));
                              if \$v5878\(0) = '1' then
                                \$14323\ := \$14274_wait603_arg\(1 to 32) & \$14302\(112 to 127);
                                \$v5847\ := eclat_not(eclat_if(eclat_not(""&\$14274_wait603_arg\(64)) & 
                                                      eclat_if(eclat_le(\$14302\(96 to 111) & eclat_resize(\$14274_wait603_arg\(33 to 63),16)) & eclat_lt(eclat_resize(\$14274_wait603_arg\(33 to 63),16) & eclat_add(\$14302\(96 to 111) & X"1770")) & eclat_false) & eclat_false));
                                if \$v5847\(0) = '1' then
                                  \$14340\ := \$14274_wait603_arg\(33 to 64) & \$14323\(32 to 47);
                                  \$14343_copy_root_in_ram604_id\ := "000000000111";
                                  \$14343_copy_root_in_ram604_arg\ := X"0" & X"3e8" & \$14274_wait603_arg\(65 to 80) & \$14340\(32 to 47) & \$14302\(96 to 111) & \$14302\(112 to 127);
                                  state_var6677 <= \$14343_copy_root_in_ram604\;
                                else
                                  \$v5846\ := \$ram_ptr_take\;
                                  if \$v5846\(0) = '1' then
                                    state_var6677 <= q_wait5845;
                                  else
                                    \$ram_ptr_take\(0) := '1';
                                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_resize(\$14274_wait603_arg\(33 to 63),16) & X"000" & X"1")));
                                    state_var6677 <= pause_getI5843;
                                  end if;
                                end if;
                              else
                                \$v5877\ := \$ram_ptr_take\;
                                if \$v5877\(0) = '1' then
                                  state_var6677 <= q_wait5876;
                                else
                                  \$ram_ptr_take\(0) := '1';
                                  \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_resize(\$14274_wait603_arg\(1 to 31),16) & X"000" & X"1")));
                                  state_var6677 <= pause_getI5874;
                                end if;
                              end if;
                            else
                              result5724 := \$14274_wait603_arg\(1 to 32) & \$14274_wait603_arg\(33 to 64) & \$14302\(80 to 95) & eclat_add(\$14302\(80 to 95) & \$14274_wait603_arg\(81 to 96)) & \$14302\(96 to 111) & \$14302\(112 to 127);
                              rdy5725 := eclat_true;
                              state_var6677 <= compute5726;
                            end if;
                          end case;
                          \$v5881\ := eclat_not(rdy5725);
                          if \$v5881\(0) = '1' then
                            result5724 := \$14302\(0 to 31) & \$14302\(32 to 63) & \$14302\(64 to 79) & \$14302\(80 to 95) & \$14302\(96 to 111) & \$14302\(112 to 127);
                          end if;
                          \$14302\ := result5724 & rdy5725;
                          rdy5722 := eclat_true;
                          state_var6676 <= compute5723;
                        end case;
                        \$14302\ := \$14302\;
                        \$14292\ := \$14302\;
                        \$v5721\ := ""&\$14292\(128);
                        if \$v5721\(0) = '1' then
                          \$14274_wait603_result\ := \$14292\(0 to 31) & \$14292\(32 to 63) & \$14292\(64 to 79);
                          \$14250\ := \$14274_wait603_result\;
                          eclat_print_string(of_string("size:"));
                          
                          eclat_print_int(eclat_if(eclat_eq(\$12199_make_block525_arg\(88 to 103) & X"000" & X"0") & X"000" & X"1" & \$12199_make_block525_arg\(88 to 103)));
                          
                          eclat_print_newline(eclat_unit);
                          
                          \$v5720\ := \$ram_ptr_take\;
                          if \$v5720\(0) = '1' then
                            state_var6675 <= q_wait5719;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$14250\(64 to 79)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= eclat_lor(eclat_lsl(eclat_resize(\$12199_make_block525_arg\(80 to 87),31) & "000"& X"00000" & X"18") & eclat_lsl(eclat_resize(
                            eclat_if(eclat_eq(\$12199_make_block525_arg\(88 to 103) & X"000" & X"0") & X"000" & X"1" & \$12199_make_block525_arg\(88 to 103)),31) & "000"& X"000000" & X"2")) & eclat_true;
                            state_var6675 <= pause_setI5717;
                          end if;
                        else
                          \$14274_wait603_arg\ := eclat_unit & \$14274_wait603_arg\(1 to 32) & \$14274_wait603_arg\(33 to 64) & \$14274_wait603_arg\(65 to 80) & \$14274_wait603_arg\(81 to 96);
                          state_var6675 <= \$14274_wait603\;
                        end if;
                      when pause_getI5884 =>
                        state_var6675 <= pause_getII5885;
                      when pause_getI5916 =>
                        state_var6675 <= pause_getII5917;
                      when pause_getI5921 =>
                        state_var6675 <= pause_getII5922;
                      when pause_getI5926 =>
                        state_var6675 <= pause_getII5927;
                      when pause_getI5937 =>
                        state_var6675 <= pause_getII5938;
                      when pause_getI5942 =>
                        state_var6675 <= pause_getII5943;
                      when pause_getI5950 =>
                        state_var6675 <= pause_getII5951;
                      when pause_getI5959 =>
                        state_var6675 <= pause_getII5960;
                      when pause_getI5969 =>
                        state_var6675 <= pause_getII5970;
                      when pause_getI5974 =>
                        state_var6675 <= pause_getII5975;
                      when pause_getI5978 =>
                        state_var6675 <= pause_getII5979;
                      when pause_getI5982 =>
                        state_var6675 <= pause_getII5983;
                      when pause_getI5986 =>
                        state_var6675 <= pause_getII5987;
                      when pause_getI5990 =>
                        state_var6675 <= pause_getII5991;
                      when pause_getI5994 =>
                        state_var6675 <= pause_getII5995;
                      when pause_getI5998 =>
                        state_var6675 <= pause_getII5999;
                      when pause_getI6002 =>
                        state_var6675 <= pause_getII6003;
                      when pause_getI6014 =>
                        state_var6675 <= pause_getII6015;
                      when pause_getI6022 =>
                        state_var6675 <= pause_getII6023;
                      when pause_getI6030 =>
                        state_var6675 <= pause_getII6031;
                      when pause_getI6038 =>
                        state_var6675 <= pause_getII6039;
                      when pause_getI6046 =>
                        state_var6675 <= pause_getII6047;
                      when pause_getI6054 =>
                        state_var6675 <= pause_getII6055;
                      when pause_getI6062 =>
                        state_var6675 <= pause_getII6063;
                      when pause_getI6070 =>
                        state_var6675 <= pause_getII6071;
                      when pause_getI6074 =>
                        state_var6675 <= pause_getII6075;
                      when pause_getI6078 =>
                        state_var6675 <= pause_getII6079;
                      when pause_getI6082 =>
                        state_var6675 <= pause_getII6083;
                      when pause_getI6086 =>
                        state_var6675 <= pause_getII6087;
                      when pause_getI6094 =>
                        state_var6675 <= pause_getII6095;
                      when pause_getI6102 =>
                        state_var6675 <= pause_getII6103;
                      when pause_getI6110 =>
                        state_var6675 <= pause_getII6111;
                      when pause_getI6122 =>
                        state_var6675 <= pause_getII6123;
                      when pause_getI6127 =>
                        state_var6675 <= pause_getII6128;
                      when pause_getI6131 =>
                        state_var6675 <= pause_getII6132;
                      when pause_getI6151 =>
                        state_var6675 <= pause_getII6152;
                      when pause_getI6155 =>
                        state_var6675 <= pause_getII6156;
                      when pause_getI6159 =>
                        state_var6675 <= pause_getII6160;
                      when pause_getI6163 =>
                        state_var6675 <= pause_getII6164;
                      when pause_getI6171 =>
                        state_var6675 <= pause_getII6172;
                      when pause_getI6179 =>
                        state_var6675 <= pause_getII6180;
                      when pause_getI6187 =>
                        state_var6675 <= pause_getII6188;
                      when pause_getI6195 =>
                        state_var6675 <= pause_getII6196;
                      when pause_getI6199 =>
                        state_var6675 <= pause_getII6200;
                      when pause_getI6203 =>
                        state_var6675 <= pause_getII6204;
                      when pause_getI6207 =>
                        state_var6675 <= pause_getII6208;
                      when pause_getI6215 =>
                        state_var6675 <= pause_getII6216;
                      when pause_getI6219 =>
                        state_var6675 <= pause_getII6220;
                      when pause_getI6223 =>
                        state_var6675 <= pause_getII6224;
                      when pause_getI6227 =>
                        state_var6675 <= pause_getII6228;
                      when pause_getI6235 =>
                        state_var6675 <= pause_getII6236;
                      when pause_getI6239 =>
                        state_var6675 <= pause_getII6240;
                      when pause_getI6243 =>
                        state_var6675 <= pause_getII6244;
                      when pause_getI6247 =>
                        state_var6675 <= pause_getII6248;
                      when pause_getI6251 =>
                        state_var6675 <= pause_getII6252;
                      when pause_getI6255 =>
                        state_var6675 <= pause_getII6256;
                      when pause_getI6259 =>
                        state_var6675 <= pause_getII6260;
                      when pause_getI6279 =>
                        state_var6675 <= pause_getII6280;
                      when pause_getI6283 =>
                        state_var6675 <= pause_getII6284;
                      when pause_getI6295 =>
                        state_var6675 <= pause_getII6296;
                      when pause_getI6299 =>
                        state_var6675 <= pause_getII6300;
                      when pause_getI6319 =>
                        state_var6675 <= pause_getII6320;
                      when pause_getI6323 =>
                        state_var6675 <= pause_getII6324;
                      when pause_getI6327 =>
                        state_var6675 <= pause_getII6328;
                      when pause_getI6331 =>
                        state_var6675 <= pause_getII6332;
                      when pause_getI6335 =>
                        state_var6675 <= pause_getII6336;
                      when pause_getI6344 =>
                        state_var6675 <= pause_getII6345;
                      when pause_getI6349 =>
                        state_var6675 <= pause_getII6350;
                      when pause_getI6353 =>
                        state_var6675 <= pause_getII6354;
                      when pause_getI6357 =>
                        state_var6675 <= pause_getII6358;
                      when pause_getI6374 =>
                        state_var6675 <= pause_getII6375;
                      when pause_getI6378 =>
                        state_var6675 <= pause_getII6379;
                      when pause_getI6394 =>
                        state_var6675 <= pause_getII6395;
                      when pause_getI6402 =>
                        state_var6675 <= pause_getII6403;
                      when pause_getI6406 =>
                        state_var6675 <= pause_getII6407;
                      when pause_getI6410 =>
                        state_var6675 <= pause_getII6411;
                      when pause_getI6431 =>
                        state_var6675 <= pause_getII6432;
                      when pause_getI6440 =>
                        state_var6675 <= pause_getII6441;
                      when pause_getI6449 =>
                        state_var6675 <= pause_getII6450;
                      when pause_getI6453 =>
                        state_var6675 <= pause_getII6454;
                      when pause_getI6462 =>
                        state_var6675 <= pause_getII6463;
                      when pause_getI6466 =>
                        state_var6675 <= pause_getII6467;
                      when pause_getI6470 =>
                        state_var6675 <= pause_getII6471;
                      when pause_getI6479 =>
                        state_var6675 <= pause_getII6480;
                      when pause_getI6483 =>
                        state_var6675 <= pause_getII6484;
                      when pause_getI6487 =>
                        state_var6675 <= pause_getII6488;
                      when pause_getI6491 =>
                        state_var6675 <= pause_getII6492;
                      when pause_getI6500 =>
                        state_var6675 <= pause_getII6501;
                      when pause_getI6504 =>
                        state_var6675 <= pause_getII6505;
                      when pause_getI6508 =>
                        state_var6675 <= pause_getII6509;
                      when pause_getI6512 =>
                        state_var6675 <= pause_getII6513;
                      when pause_getI6524 =>
                        state_var6675 <= pause_getII6525;
                      when pause_getI6532 =>
                        state_var6675 <= pause_getII6533;
                      when pause_getI6537 =>
                        state_var6675 <= pause_getII6538;
                      when pause_getI6545 =>
                        state_var6675 <= pause_getII6546;
                      when pause_getI6559 =>
                        state_var6675 <= pause_getII6560;
                      when pause_getI6563 =>
                        state_var6675 <= pause_getII6564;
                      when pause_getI6567 =>
                        state_var6675 <= pause_getII6568;
                      when pause_getI6571 =>
                        state_var6675 <= pause_getII6572;
                      when pause_getI6583 =>
                        state_var6675 <= pause_getII6584;
                      when pause_getI6596 =>
                        state_var6675 <= pause_getII6597;
                      when pause_getI6605 =>
                        state_var6675 <= pause_getII6606;
                      when pause_getI6632 =>
                        state_var6675 <= pause_getII6633;
                      when pause_getI6637 =>
                        state_var6675 <= pause_getII6638;
                      when pause_getI6642 =>
                        state_var6675 <= pause_getII6643;
                      when pause_getI6647 =>
                        state_var6675 <= pause_getII6648;
                      when pause_getI6652 =>
                        state_var6675 <= pause_getII6653;
                      when pause_getII5885 =>
                        \$ram_ptr_take\(0) := '0';
                        \$14196\ := \$ram_value\;
                        \$12235_apply579_result\ := eclat_resize(\$14196\(0 to 30),16) & \$12235_apply579_arg\(60 to 91) & \$14192_sp\ & \$12235_apply579_arg\(60 to 91) & \$12235_apply579_arg\(3 to 10) & \$12235_apply579_arg\(150 to 165) & \$12235_apply579_arg\(108 to 109);
                        result5714 := \$12235_apply579_result\;
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII5917 =>
                        \$ram_ptr_take\(0) := '0';
                        \$14227_v\ := \$ram_value\;
                        \$14186\ := \$14227_v\ & eclat_sub(\$14183\(32 to 47) & X"000" & X"1");
                        \$v5915\ := ""&\$12235_apply579_arg\(11);
                        if \$v5915\(0) = '1' then
                          \$14189_sp\ := eclat_add(eclat_sub(\$14186\(32 to 47) & \$12235_apply579_arg\(12 to 27)) & \$12235_apply579_arg\(28 to 43));
                          \$v5902\ := ""&\$12235_apply579_arg\(2);
                          if \$v5902\(0) = '1' then
                            \$v5901\ := \$ram_ptr_take\;
                            if \$v5901\(0) = '1' then
                              state_var6675 <= q_wait5900;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(\$14189_sp\));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$14186\(0 to 31);
                              state_var6675 <= pause_setI5898;
                            end if;
                          else
                            \$14190_sp\ := \$14189_sp\;
                            \$v5897\ := ""&\$12235_apply579_arg\(1);
                            if \$v5897\(0) = '1' then
                              \$v5896\ := \$ram_ptr_take\;
                              if \$v5896\(0) = '1' then
                                state_var6675 <= q_wait5895;
                              else
                                \$ram_ptr_take\(0) := '1';
                                \$ram_ptr_write\ <= to_integer(unsigned(\$14190_sp\));
                                \$ram_write_request\ <= '1';
                                \$ram_write\ <= \$14183\(0 to 31);
                                state_var6675 <= pause_setI5893;
                              end if;
                            else
                              \$14191_sp\ := \$14190_sp\;
                              \$v5892\ := ""&\$12235_apply579_arg\(0);
                              if \$v5892\(0) = '1' then
                                \$v5891\ := \$ram_ptr_take\;
                                if \$v5891\(0) = '1' then
                                  state_var6675 <= q_wait5890;
                                else
                                  \$ram_ptr_take\(0) := '1';
                                  \$ram_ptr_write\ <= to_integer(unsigned(\$14191_sp\));
                                  \$ram_write_request\ <= '1';
                                  \$ram_write\ <= \$14180\(0 to 31);
                                  state_var6675 <= pause_setI5888;
                                end if;
                              else
                                \$14192_sp\ := \$14191_sp\;
                                \$v5887\ := \$ram_ptr_take\;
                                if \$v5887\(0) = '1' then
                                  state_var6675 <= q_wait5886;
                                else
                                  \$ram_ptr_take\(0) := '1';
                                  \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12235_apply579_arg\(60 to 90),16) & X"000" & X"0") & X"000" & X"1")));
                                  state_var6675 <= pause_getI5884;
                                end if;
                              end if;
                            end if;
                          end if;
                        else
                          \$v5914\ := \$ram_ptr_take\;
                          if \$v5914\(0) = '1' then
                            state_var6675 <= q_wait5913;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$14186\(32 to 47)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= eclat_resize(\$12235_apply579_arg\(142 to 149),31) & eclat_true;
                            state_var6675 <= pause_setI5911;
                          end if;
                        end if;
                      when pause_getII5922 =>
                        \$ram_ptr_take\(0) := '0';
                        \$14230_v\ := \$ram_value\;
                        \$14183\ := \$14230_v\ & eclat_sub(\$14180\(32 to 47) & X"000" & X"1");
                        \$v5920\ := ""&\$12235_apply579_arg\(2);
                        if \$v5920\(0) = '1' then
                          \$v5919\ := \$ram_ptr_take\;
                          if \$v5919\(0) = '1' then
                            state_var6675 <= q_wait5918;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$14183\(32 to 47) & X"000" & X"1")));
                            state_var6675 <= pause_getI5916;
                          end if;
                        else
                          \$14186\ := "000"& X"000000" & X"1" & eclat_true & \$14183\(32 to 47);
                          \$v5915\ := ""&\$12235_apply579_arg\(11);
                          if \$v5915\(0) = '1' then
                            \$14189_sp\ := eclat_add(eclat_sub(\$14186\(32 to 47) & \$12235_apply579_arg\(12 to 27)) & \$12235_apply579_arg\(28 to 43));
                            \$v5902\ := ""&\$12235_apply579_arg\(2);
                            if \$v5902\(0) = '1' then
                              \$v5901\ := \$ram_ptr_take\;
                              if \$v5901\(0) = '1' then
                                state_var6675 <= q_wait5900;
                              else
                                \$ram_ptr_take\(0) := '1';
                                \$ram_ptr_write\ <= to_integer(unsigned(\$14189_sp\));
                                \$ram_write_request\ <= '1';
                                \$ram_write\ <= \$14186\(0 to 31);
                                state_var6675 <= pause_setI5898;
                              end if;
                            else
                              \$14190_sp\ := \$14189_sp\;
                              \$v5897\ := ""&\$12235_apply579_arg\(1);
                              if \$v5897\(0) = '1' then
                                \$v5896\ := \$ram_ptr_take\;
                                if \$v5896\(0) = '1' then
                                  state_var6675 <= q_wait5895;
                                else
                                  \$ram_ptr_take\(0) := '1';
                                  \$ram_ptr_write\ <= to_integer(unsigned(\$14190_sp\));
                                  \$ram_write_request\ <= '1';
                                  \$ram_write\ <= \$14183\(0 to 31);
                                  state_var6675 <= pause_setI5893;
                                end if;
                              else
                                \$14191_sp\ := \$14190_sp\;
                                \$v5892\ := ""&\$12235_apply579_arg\(0);
                                if \$v5892\(0) = '1' then
                                  \$v5891\ := \$ram_ptr_take\;
                                  if \$v5891\(0) = '1' then
                                    state_var6675 <= q_wait5890;
                                  else
                                    \$ram_ptr_take\(0) := '1';
                                    \$ram_ptr_write\ <= to_integer(unsigned(\$14191_sp\));
                                    \$ram_write_request\ <= '1';
                                    \$ram_write\ <= \$14180\(0 to 31);
                                    state_var6675 <= pause_setI5888;
                                  end if;
                                else
                                  \$14192_sp\ := \$14191_sp\;
                                  \$v5887\ := \$ram_ptr_take\;
                                  if \$v5887\(0) = '1' then
                                    state_var6675 <= q_wait5886;
                                  else
                                    \$ram_ptr_take\(0) := '1';
                                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12235_apply579_arg\(60 to 90),16) & X"000" & X"0") & X"000" & X"1")));
                                    state_var6675 <= pause_getI5884;
                                  end if;
                                end if;
                              end if;
                            end if;
                          else
                            \$v5914\ := \$ram_ptr_take\;
                            if \$v5914\(0) = '1' then
                              state_var6675 <= q_wait5913;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(\$14186\(32 to 47)));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= eclat_resize(\$12235_apply579_arg\(142 to 149),31) & eclat_true;
                              state_var6675 <= pause_setI5911;
                            end if;
                          end if;
                        end if;
                      when pause_getII5927 =>
                        \$ram_ptr_take\(0) := '0';
                        \$14233_v\ := \$ram_value\;
                        \$14180\ := \$14233_v\ & eclat_sub(\$12235_apply579_arg\(92 to 107) & X"000" & X"1");
                        \$v5925\ := ""&\$12235_apply579_arg\(1);
                        if \$v5925\(0) = '1' then
                          \$v5924\ := \$ram_ptr_take\;
                          if \$v5924\(0) = '1' then
                            state_var6675 <= q_wait5923;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$14180\(32 to 47) & X"000" & X"1")));
                            state_var6675 <= pause_getI5921;
                          end if;
                        else
                          \$14183\ := "000"& X"000000" & X"1" & eclat_true & \$14180\(32 to 47);
                          \$v5920\ := ""&\$12235_apply579_arg\(2);
                          if \$v5920\(0) = '1' then
                            \$v5919\ := \$ram_ptr_take\;
                            if \$v5919\(0) = '1' then
                              state_var6675 <= q_wait5918;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$14183\(32 to 47) & X"000" & X"1")));
                              state_var6675 <= pause_getI5916;
                            end if;
                          else
                            \$14186\ := "000"& X"000000" & X"1" & eclat_true & \$14183\(32 to 47);
                            \$v5915\ := ""&\$12235_apply579_arg\(11);
                            if \$v5915\(0) = '1' then
                              \$14189_sp\ := eclat_add(eclat_sub(\$14186\(32 to 47) & \$12235_apply579_arg\(12 to 27)) & \$12235_apply579_arg\(28 to 43));
                              \$v5902\ := ""&\$12235_apply579_arg\(2);
                              if \$v5902\(0) = '1' then
                                \$v5901\ := \$ram_ptr_take\;
                                if \$v5901\(0) = '1' then
                                  state_var6675 <= q_wait5900;
                                else
                                  \$ram_ptr_take\(0) := '1';
                                  \$ram_ptr_write\ <= to_integer(unsigned(\$14189_sp\));
                                  \$ram_write_request\ <= '1';
                                  \$ram_write\ <= \$14186\(0 to 31);
                                  state_var6675 <= pause_setI5898;
                                end if;
                              else
                                \$14190_sp\ := \$14189_sp\;
                                \$v5897\ := ""&\$12235_apply579_arg\(1);
                                if \$v5897\(0) = '1' then
                                  \$v5896\ := \$ram_ptr_take\;
                                  if \$v5896\(0) = '1' then
                                    state_var6675 <= q_wait5895;
                                  else
                                    \$ram_ptr_take\(0) := '1';
                                    \$ram_ptr_write\ <= to_integer(unsigned(\$14190_sp\));
                                    \$ram_write_request\ <= '1';
                                    \$ram_write\ <= \$14183\(0 to 31);
                                    state_var6675 <= pause_setI5893;
                                  end if;
                                else
                                  \$14191_sp\ := \$14190_sp\;
                                  \$v5892\ := ""&\$12235_apply579_arg\(0);
                                  if \$v5892\(0) = '1' then
                                    \$v5891\ := \$ram_ptr_take\;
                                    if \$v5891\(0) = '1' then
                                      state_var6675 <= q_wait5890;
                                    else
                                      \$ram_ptr_take\(0) := '1';
                                      \$ram_ptr_write\ <= to_integer(unsigned(\$14191_sp\));
                                      \$ram_write_request\ <= '1';
                                      \$ram_write\ <= \$14180\(0 to 31);
                                      state_var6675 <= pause_setI5888;
                                    end if;
                                  else
                                    \$14192_sp\ := \$14191_sp\;
                                    \$v5887\ := \$ram_ptr_take\;
                                    if \$v5887\(0) = '1' then
                                      state_var6675 <= q_wait5886;
                                    else
                                      \$ram_ptr_take\(0) := '1';
                                      \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12235_apply579_arg\(60 to 90),16) & X"000" & X"0") & X"000" & X"1")));
                                      state_var6675 <= pause_getI5884;
                                    end if;
                                  end if;
                                end if;
                              end if;
                            else
                              \$v5914\ := \$ram_ptr_take\;
                              if \$v5914\(0) = '1' then
                                state_var6675 <= q_wait5913;
                              else
                                \$ram_ptr_take\(0) := '1';
                                \$ram_ptr_write\ <= to_integer(unsigned(\$14186\(32 to 47)));
                                \$ram_write_request\ <= '1';
                                \$ram_write\ <= eclat_resize(\$12235_apply579_arg\(142 to 149),31) & eclat_true;
                                state_var6675 <= pause_setI5911;
                              end if;
                            end if;
                          end if;
                        end if;
                      when pause_getII5938 =>
                        \$ram_ptr_take\(0) := '0';
                        \$14082_v\ := \$ram_value\;
                        \$v5936\ := \$12237_binop_int584_arg\(0 to 31);
                        case \$v5936\ is
                        when X"0000000" & X"0" =>
                          \$14086_res\ := eclat_add(\$12237_binop_int584_arg\(48 to 78) & \$14082_v\(0 to 30));
                          \$12237_binop_int584_result\ := eclat_add(\$12237_binop_int584_arg\(32 to 47) & X"000" & X"1") & \$14086_res\ & eclat_true & eclat_sub(\$12237_binop_int584_arg\(80 to 95) & X"000" & X"1") & \$12237_binop_int584_arg\(96 to 151) & \$12237_binop_int584_arg\(152 to 153);
                          result5714 := \$12237_binop_int584_result\;
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        when X"0000000" & X"1" =>
                          \$14086_res\ := eclat_sub(\$12237_binop_int584_arg\(48 to 78) & \$14082_v\(0 to 30));
                          \$12237_binop_int584_result\ := eclat_add(\$12237_binop_int584_arg\(32 to 47) & X"000" & X"1") & \$14086_res\ & eclat_true & eclat_sub(\$12237_binop_int584_arg\(80 to 95) & X"000" & X"1") & \$12237_binop_int584_arg\(96 to 151) & \$12237_binop_int584_arg\(152 to 153);
                          result5714 := \$12237_binop_int584_result\;
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        when X"0000000" & X"2" =>
                          \$14086_res\ := eclat_mult(\$12237_binop_int584_arg\(48 to 78) & \$14082_v\(0 to 30));
                          \$12237_binop_int584_result\ := eclat_add(\$12237_binop_int584_arg\(32 to 47) & X"000" & X"1") & \$14086_res\ & eclat_true & eclat_sub(\$12237_binop_int584_arg\(80 to 95) & X"000" & X"1") & \$12237_binop_int584_arg\(96 to 151) & \$12237_binop_int584_arg\(152 to 153);
                          result5714 := \$12237_binop_int584_result\;
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        when X"0000000" & X"3" =>
                          \$v5933\ := eclat_eq(\$14082_v\(0 to 30) & "000"& X"000000" & X"0");
                          if \$v5933\(0) = '1' then
                            \$14086_res\ := "000"& X"000000" & X"0";
                            \$12237_binop_int584_result\ := eclat_add(\$12237_binop_int584_arg\(32 to 47) & X"000" & X"1") & \$14086_res\ & eclat_true & eclat_sub(\$12237_binop_int584_arg\(80 to 95) & X"000" & X"1") & \$12237_binop_int584_arg\(96 to 151) & \$12237_binop_int584_arg\(152 to 153);
                            result5714 := \$12237_binop_int584_result\;
                            rdy5715 := eclat_true;
                            state_var6675 <= compute5716;
                          else
                            \$14090_modulo609_arg\ := eclat_abs(\$12237_binop_int584_arg\(48 to 78)) & eclat_abs(\$14082_v\(0 to 30));
                            state_var6675 <= \$14090_modulo609\;
                          end if;
                        when X"0000000" & X"4" =>
                          \$v5935\ := eclat_eq(\$14082_v\(0 to 30) & "000"& X"000000" & X"0");
                          if \$v5935\(0) = '1' then
                            \$14086_res\ := "000"& X"000000" & X"0";
                            \$12237_binop_int584_result\ := eclat_add(\$12237_binop_int584_arg\(32 to 47) & X"000" & X"1") & \$14086_res\ & eclat_true & eclat_sub(\$12237_binop_int584_arg\(80 to 95) & X"000" & X"1") & \$12237_binop_int584_arg\(96 to 151) & \$12237_binop_int584_arg\(152 to 153);
                            result5714 := \$12237_binop_int584_result\;
                            rdy5715 := eclat_true;
                            state_var6675 <= compute5716;
                          else
                            \$14105_modulo609_arg\ := eclat_abs(\$12237_binop_int584_arg\(48 to 78)) & eclat_abs(\$14082_v\(0 to 30));
                            state_var6675 <= \$14105_modulo609\;
                          end if;
                        when X"0000000" & X"5" =>
                          \$14086_res\ := eclat_land(\$12237_binop_int584_arg\(48 to 78) & \$14082_v\(0 to 30));
                          \$12237_binop_int584_result\ := eclat_add(\$12237_binop_int584_arg\(32 to 47) & X"000" & X"1") & \$14086_res\ & eclat_true & eclat_sub(\$12237_binop_int584_arg\(80 to 95) & X"000" & X"1") & \$12237_binop_int584_arg\(96 to 151) & \$12237_binop_int584_arg\(152 to 153);
                          result5714 := \$12237_binop_int584_result\;
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        when X"0000000" & X"6" =>
                          \$14086_res\ := eclat_lor(\$12237_binop_int584_arg\(48 to 78) & \$14082_v\(0 to 30));
                          \$12237_binop_int584_result\ := eclat_add(\$12237_binop_int584_arg\(32 to 47) & X"000" & X"1") & \$14086_res\ & eclat_true & eclat_sub(\$12237_binop_int584_arg\(80 to 95) & X"000" & X"1") & \$12237_binop_int584_arg\(96 to 151) & \$12237_binop_int584_arg\(152 to 153);
                          result5714 := \$12237_binop_int584_result\;
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        when X"0000000" & X"7" =>
                          \$14086_res\ := eclat_lxor(\$12237_binop_int584_arg\(48 to 78) & \$14082_v\(0 to 30));
                          \$12237_binop_int584_result\ := eclat_add(\$12237_binop_int584_arg\(32 to 47) & X"000" & X"1") & \$14086_res\ & eclat_true & eclat_sub(\$12237_binop_int584_arg\(80 to 95) & X"000" & X"1") & \$12237_binop_int584_arg\(96 to 151) & \$12237_binop_int584_arg\(152 to 153);
                          result5714 := \$12237_binop_int584_result\;
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        when X"0000000" & X"8" =>
                          \$14086_res\ := eclat_lsl(\$12237_binop_int584_arg\(48 to 78) & \$14082_v\(0 to 30));
                          \$12237_binop_int584_result\ := eclat_add(\$12237_binop_int584_arg\(32 to 47) & X"000" & X"1") & \$14086_res\ & eclat_true & eclat_sub(\$12237_binop_int584_arg\(80 to 95) & X"000" & X"1") & \$12237_binop_int584_arg\(96 to 151) & \$12237_binop_int584_arg\(152 to 153);
                          result5714 := \$12237_binop_int584_result\;
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        when X"0000000" & X"9" =>
                          \$14086_res\ := eclat_lsr(\$12237_binop_int584_arg\(48 to 78) & \$14082_v\(0 to 30));
                          \$12237_binop_int584_result\ := eclat_add(\$12237_binop_int584_arg\(32 to 47) & X"000" & X"1") & \$14086_res\ & eclat_true & eclat_sub(\$12237_binop_int584_arg\(80 to 95) & X"000" & X"1") & \$12237_binop_int584_arg\(96 to 151) & \$12237_binop_int584_arg\(152 to 153);
                          result5714 := \$12237_binop_int584_result\;
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        when X"0000000" & X"a" =>
                          \$14086_res\ := eclat_asr(\$12237_binop_int584_arg\(48 to 78) & \$14082_v\(0 to 30));
                          \$12237_binop_int584_result\ := eclat_add(\$12237_binop_int584_arg\(32 to 47) & X"000" & X"1") & \$14086_res\ & eclat_true & eclat_sub(\$12237_binop_int584_arg\(80 to 95) & X"000" & X"1") & \$12237_binop_int584_arg\(96 to 151) & \$12237_binop_int584_arg\(152 to 153);
                          result5714 := \$12237_binop_int584_result\;
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        when X"0000000" & X"b" =>
                          \$14086_res\ := eclat_if(eclat_lt(\$12237_binop_int584_arg\(48 to 78) & "000"& X"000000" & X"0") & 
                                          eclat_if(eclat_lt(\$14082_v\(0 to 30) & "000"& X"000000" & X"0") & 
                                          eclat_if(eclat_gt(\$12237_binop_int584_arg\(48 to 78) & \$14082_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"0") & 
                                          eclat_if(eclat_lt(\$14082_v\(0 to 30) & "000"& X"000000" & X"0") & "000"& X"000000" & X"0" & 
                                          eclat_if(eclat_lt(\$12237_binop_int584_arg\(48 to 78) & \$14082_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                          \$12237_binop_int584_result\ := eclat_add(\$12237_binop_int584_arg\(32 to 47) & X"000" & X"1") & \$14086_res\ & eclat_true & eclat_sub(\$12237_binop_int584_arg\(80 to 95) & X"000" & X"1") & \$12237_binop_int584_arg\(96 to 151) & \$12237_binop_int584_arg\(152 to 153);
                          result5714 := \$12237_binop_int584_result\;
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        when X"0000000" & X"c" =>
                          \$14086_res\ := eclat_if(eclat_lt(\$12237_binop_int584_arg\(48 to 78) & "000"& X"000000" & X"0") & 
                                          eclat_if(eclat_lt(\$14082_v\(0 to 30) & "000"& X"000000" & X"0") & 
                                          eclat_if(eclat_le(\$12237_binop_int584_arg\(48 to 78) & \$14082_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & "000"& X"000000" & X"1") & 
                                          eclat_if(eclat_lt(\$14082_v\(0 to 30) & "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & 
                                          eclat_if(eclat_ge(\$12237_binop_int584_arg\(48 to 78) & \$14082_v\(0 to 30)) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0")));
                          \$12237_binop_int584_result\ := eclat_add(\$12237_binop_int584_arg\(32 to 47) & X"000" & X"1") & \$14086_res\ & eclat_true & eclat_sub(\$12237_binop_int584_arg\(80 to 95) & X"000" & X"1") & \$12237_binop_int584_arg\(96 to 151) & \$12237_binop_int584_arg\(152 to 153);
                          result5714 := \$12237_binop_int584_result\;
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        when others =>
                          \$14086_res\ := "000"& X"000000" & X"0";
                          \$12237_binop_int584_result\ := eclat_add(\$12237_binop_int584_arg\(32 to 47) & X"000" & X"1") & \$14086_res\ & eclat_true & eclat_sub(\$12237_binop_int584_arg\(80 to 95) & X"000" & X"1") & \$12237_binop_int584_arg\(96 to 151) & \$12237_binop_int584_arg\(152 to 153);
                          result5714 := \$12237_binop_int584_result\;
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        end case;
                      when pause_getII5943 =>
                        \$ram_ptr_take\(0) := '0';
                        \$14048_v\ := \$ram_value\;
                        \$12238_compare585_id\ := "000000001101";
                        \$12238_compare585_arg\ := \$12239_binop_compare586_arg\(0 to 31) & \$12239_binop_compare586_arg\(48 to 78) & \$14048_v\(0 to 30);
                        state_var6675 <= \$12238_compare585\;
                      when pause_getII5951 =>
                        \$ram_ptr_take\(0) := '0';
                        \$14003_v\ := \$ram_value\;
                        \$v5949\ := \$ram_ptr_take\;
                        if \$v5949\(0) = '1' then
                          state_var6675 <= q_wait5948;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$13996\(64 to 94),16) & X"000" & X"2") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$14003_v\;
                          state_var6675 <= pause_setI5946;
                        end if;
                      when pause_getII5960 =>
                        \$ram_ptr_take\(0) := '0';
                        \$14014_v\ := \$ram_value\;
                        \$v5958\ := \$ram_ptr_take\;
                        if \$v5958\(0) = '1' then
                          state_var6675 <= q_wait5957;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$13996\(64 to 94),16) & X"000" & X"1") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$14014_v\;
                          state_var6675 <= pause_setI5955;
                        end if;
                      when pause_getII5970 =>
                        \$code_ptr_take\(0) := '0';
                        \$13972_arg\ := \$code_value\;
                        \$12241_branch_if589_result\ := eclat_add(eclat_add(\$12241_branch_if589_arg\(1 to 16) & X"000" & X"1") & eclat_resize(\$13972_arg\,16)) & \$12241_branch_if589_arg\(17 to 48) & \$12241_branch_if589_arg\(49 to 64) & \$12241_branch_if589_arg\(65 to 120) & \$12241_branch_if589_arg\(121 to 122);
                        result5714 := \$12241_branch_if589_result\;
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII5975 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13328_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$13328_v\ & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII5979 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13333_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$13333_v\ & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII5983 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13338_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$13338_v\ & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII5987 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13343_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$13343_v\ & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII5991 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13348_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$13348_v\ & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII5995 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13353_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$13353_v\ & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII5999 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13358_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$13358_v\ & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6003 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13363_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$13363_v\ & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6015 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13377_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$13377_v\ & eclat_add(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6023 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13386_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$13386_v\ & eclat_add(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6031 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13395_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$13395_v\ & eclat_add(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6039 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13404_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$13404_v\ & eclat_add(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6047 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13413_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$13413_v\ & eclat_add(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6055 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13422_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$13422_v\ & eclat_add(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6063 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13431_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$13431_v\ & eclat_add(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6071 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13442\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$13442\ & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6075 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13453\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$13453\ & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6079 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13464\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$13464\ & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6083 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13475\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$13475\ & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6087 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13487\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$13487\ & eclat_add(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6095 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13500\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$13500\ & eclat_add(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6103 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13513\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$13513\ & eclat_add(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6111 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13526\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$13526\ & eclat_add(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6123 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13589\ := \$ram_value\;
                        \$v6121\ := \$ram_ptr_take\;
                        if \$v6121\(0) = '1' then
                          state_var6675 <= q_wait6120;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$13539_loop_push598_arg\(0 to 15)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$13589\;
                          state_var6675 <= pause_setI6118;
                        end if;
                      when pause_getII6128 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13547_next_env\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$12190\(16 to 47) & \$13543_sp\ & \$13547_next_env\ & eclat_add(\$12190\(96 to 103) & eclat_sub(eclat_resize(eclat_resize(eclat_lsr(eclat_resize(eclat_resize(\$13538_hd\(0 to 30),16),31) & "000"& X"000000" & X"2"),16),8) & "00000010")) & \$12190\(104 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6132 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13538_hd\ := \$ram_value\;
                        \$13539_loop_push598_arg\ := \$12190\(48 to 63) & "00000000" & \$12190\(64 to 95) & eclat_resize(eclat_resize(eclat_lsr(eclat_resize(eclat_resize(\$13538_hd\(0 to 30),16),31) & "000"& X"000000" & X"2"),16),8);
                        state_var6675 <= \$13539_loop_push598\;
                      when pause_getII6152 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13646_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$13646_v\ & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6156 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13661_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$13661_v\ & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6160 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13676_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$13676_v\ & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6164 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13691_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$13691_v\ & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6172 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13699_v\ := \$ram_value\;
                        \$v6170\ := \$ram_ptr_take\;
                        if \$v6170\(0) = '1' then
                          state_var6675 <= q_wait6169;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & X"000" & X"0") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$13699_v\;
                          state_var6675 <= pause_setI6167;
                        end if;
                      when pause_getII6180 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13712_v\ := \$ram_value\;
                        \$v6178\ := \$ram_ptr_take\;
                        if \$v6178\(0) = '1' then
                          state_var6675 <= q_wait6177;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & X"000" & X"1") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$13712_v\;
                          state_var6675 <= pause_setI6175;
                        end if;
                      when pause_getII6188 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13725_v\ := \$ram_value\;
                        \$v6186\ := \$ram_ptr_take\;
                        if \$v6186\(0) = '1' then
                          state_var6675 <= q_wait6185;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & X"000" & X"2") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$13725_v\;
                          state_var6675 <= pause_setI6183;
                        end if;
                      when pause_getII6196 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13738_v\ := \$ram_value\;
                        \$v6194\ := \$ram_ptr_take\;
                        if \$v6194\(0) = '1' then
                          state_var6675 <= q_wait6193;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & X"000" & X"3") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$13738_v\;
                          state_var6675 <= pause_setI6191;
                        end if;
                      when pause_getII6200 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13754_hd\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & eclat_resize(eclat_resize(eclat_lsr(eclat_resize(eclat_resize(\$13754_hd\(0 to 30),16),31) & "000"& X"000000" & X"2"),16),31) & eclat_true & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6204 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13774_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$13774_v\ & eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6208 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13767_v\ := \$ram_value\;
                        \$v6206\ := \$ram_ptr_take\;
                        if \$v6206\(0) = '1' then
                          state_var6675 <= q_wait6205;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & eclat_resize(\$13767_v\(0 to 30),16)) & X"000" & X"1")));
                          state_var6675 <= pause_getI6203;
                        end if;
                      when pause_getII6216 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13785_v\ := \$ram_value\;
                        \$v6214\ := \$ram_ptr_take\;
                        if \$v6214\(0) = '1' then
                          state_var6675 <= q_wait6213;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & eclat_resize(\$13784_v\(0 to 30),16)) & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$13785_v\;
                          state_var6675 <= pause_setI6211;
                        end if;
                      when pause_getII6220 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13784_v\ := \$ram_value\;
                        \$v6218\ := \$ram_ptr_take\;
                        if \$v6218\(0) = '1' then
                          state_var6675 <= q_wait6217;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6215;
                        end if;
                      when pause_getII6224 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13814_next_acc\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$13814_next_acc\ & eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6228 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13807_v\ := \$ram_value\;
                        \$v6226\ := \$ram_ptr_take\;
                        if \$v6226\(0) = '1' then
                          state_var6675 <= q_wait6225;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & eclat_resize(\$13807_v\(0 to 30),16)) & X"000" & X"1")));
                          state_var6675 <= pause_getI6223;
                        end if;
                      when pause_getII6236 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13825_v\ := \$ram_value\;
                        \$v6234\ := \$ram_ptr_take\;
                        if \$v6234\(0) = '1' then
                          state_var6675 <= q_wait6233;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & eclat_resize(\$13824_v\(0 to 30),16)) & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$13825_v\;
                          state_var6675 <= pause_setI6231;
                        end if;
                      when pause_getII6240 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13824_v\ := \$ram_value\;
                        \$v6238\ := \$ram_ptr_take\;
                        if \$v6238\(0) = '1' then
                          state_var6675 <= q_wait6237;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6235;
                        end if;
                      when pause_getII6244 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13854_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$12190\(16 to 47) & eclat_sub(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1") & X"000" & X"2") & \$12190\(64 to 95) & \$12190\(96 to 103) & eclat_resize(\$13854_v\(0 to 30),16) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6248 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13878_v\ := \$ram_value\;
                        result5714 := eclat_resize(\$13869_v\(0 to 30),16) & \$12190\(16 to 47) & eclat_sub(eclat_sub(eclat_sub(eclat_sub(\$12190\(104 to 119) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1") & X"000" & X"1") & \$13877_v\ & eclat_resize(\$13878_v\(0 to 30),8) & eclat_resize(\$13873_v\(0 to 30),16) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6252 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13877_v\ := \$ram_value\;
                        \$v6250\ := \$ram_ptr_take\;
                        if \$v6250\(0) = '1' then
                          state_var6675 <= q_wait6249;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_sub(eclat_sub(\$12190\(104 to 119) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6247;
                        end if;
                      when pause_getII6256 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13873_v\ := \$ram_value\;
                        \$v6254\ := \$ram_ptr_take\;
                        if \$v6254\(0) = '1' then
                          state_var6675 <= q_wait6253;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_sub(\$12190\(104 to 119) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6251;
                        end if;
                      when pause_getII6260 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13869_v\ := \$ram_value\;
                        \$v6258\ := \$ram_ptr_take\;
                        if \$v6258\(0) = '1' then
                          state_var6675 <= q_wait6257;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(104 to 119) & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6255;
                        end if;
                      when pause_getII6280 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12604_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$12604_v\ & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6284 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12612_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"2") & \$12612_v\ & eclat_add(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6296 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12634\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"2") & \$12634\ & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6300 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12648\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"2") & \$12648\ & eclat_add(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6320 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12683\ := \$ram_value\;
                        result5714 := eclat_resize(\$12683\(0 to 30),16) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(16 to 47) & eclat_sub(eclat_resize(\$12246_argument1\,8) & "00000001") & \$12190\(104 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6324 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12754\ := \$ram_value\;
                        result5714 := eclat_resize(\$12754\(0 to 30),16) & \$12190\(16 to 47) & eclat_sub(\$12190\(48 to 63) & eclat_resize(\$12246_argument1\,16)) & \$12190\(16 to 47) & eclat_sub(\$12190\(96 to 103) & "00000001") & \$12190\(104 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6328 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12714_v\ := \$ram_value\;
                        result5714 := eclat_resize(\$12709_v\(0 to 30),16) & \$12190\(16 to 47) & eclat_sub(eclat_sub(eclat_sub(eclat_sub(\$12190\(48 to 63) & eclat_resize(\$12246_argument1\,16)) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1") & \$12713_v\ & eclat_resize(\$12714_v\(0 to 30),8) & \$12190\(104 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6332 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12713_v\ := \$ram_value\;
                        \$v6330\ := \$ram_ptr_take\;
                        if \$v6330\(0) = '1' then
                          state_var6675 <= q_wait6329;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_sub(eclat_sub(\$12190\(48 to 63) & eclat_resize(\$12246_argument1\,16)) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6327;
                        end if;
                      when pause_getII6336 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12709_v\ := \$ram_value\;
                        \$v6334\ := \$ram_ptr_take\;
                        if \$v6334\(0) = '1' then
                          state_var6675 <= q_wait6333;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_sub(\$12190\(48 to 63) & eclat_resize(\$12246_argument1\,16)) & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6331;
                        end if;
                      when pause_getII6345 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12820_v\ := \$ram_value\;
                        \$v6343\ := \$ram_ptr_take\;
                        if \$v6343\(0) = '1' then
                          state_var6675 <= q_wait6342;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12782_w597_arg\(32 to 62),16) & eclat_resize(eclat_add(\$12782_w597_arg\(0 to 7) & "00000010"),16)) & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12820_v\;
                          state_var6675 <= pause_setI6340;
                        end if;
                      when pause_getII6350 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12789_v\ := \$ram_value\;
                        result5714 := eclat_resize(\$12784_v\(0 to 30),16) & \$12770\(64 to 95) & eclat_sub(eclat_sub(eclat_sub(\$12783_sp\ & X"000" & X"1") & X"000" & X"1") & X"000" & X"1") & \$12788_v\ & eclat_resize(\$12789_v\(0 to 30),8) & \$12190\(104 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6354 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12788_v\ := \$ram_value\;
                        \$v6352\ := \$ram_ptr_take\;
                        if \$v6352\(0) = '1' then
                          state_var6675 <= q_wait6351;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_sub(\$12783_sp\ & X"000" & X"1") & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6349;
                        end if;
                      when pause_getII6358 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12784_v\ := \$ram_value\;
                        \$v6356\ := \$ram_ptr_take\;
                        if \$v6356\(0) = '1' then
                          state_var6675 <= q_wait6355;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12783_sp\ & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6353;
                        end if;
                      when pause_getII6375 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12872_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"2") & \$12872_v\ & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6379 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12878_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"2") & \$12878_v\ & eclat_add(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6395 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12920_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"2") & \$12920_v\ & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6403 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12929_v\ := \$ram_value\;
                        \$v6401\ := \$ram_ptr_take\;
                        if \$v6401\(0) = '1' then
                          state_var6675 <= q_wait6400;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & eclat_resize(\$12246_argument1\,16)) & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12929_v\;
                          state_var6675 <= pause_setI6398;
                        end if;
                      when pause_getII6407 =>
                        \$code_ptr_take\(0) := '0';
                        \$12954\ := \$code_value\;
                        result5714 := eclat_add(eclat_add(\$12190\(0 to 15) & X"000" & X"2") & eclat_resize(\$12954\,16)) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6411 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12965_hd\ := \$ram_value\;
                        \$12953_ofs\ := eclat_add(eclat_resize(\$12246_argument1\,16) & eclat_lsr(eclat_resize(\$12965_hd\(0 to 30),16) & X"00" & X"18"));
                        \$v6409\ := \$code_ptr_take\;
                        if \$v6409\(0) = '1' then
                          state_var6675 <= q_wait6408;
                        else
                          \$code_ptr_take\(0) := '1';
                          \$code_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(\$12190\(0 to 15) & X"000" & X"2") & \$12953_ofs\)));
                          state_var6675 <= pause_getI6406;
                        end if;
                      when pause_getII6432 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13035_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"2") & \$13023\(0 to 31) & eclat_sub(\$13023\(80 to 95) & X"000" & X"1") & \$13035_v\ & \$13023\(128 to 135) & \$13023\(136 to 151) & \$13023\(152 to 153);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6441 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13064_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"2") & \$13052\(0 to 31) & eclat_sub(\$13052\(80 to 95) & X"000" & X"1") & \$13064_v\ & \$13052\(128 to 135) & \$13052\(136 to 151) & \$13052\(152 to 153);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6450 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6448\ := \$ram_ptr_take\;
                        if \$v6448\(0) = '1' then
                          state_var6675 <= q_wait6447;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_sub(\$12190\(48 to 63) & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(64 to 95);
                          state_var6675 <= pause_setI6445;
                        end if;
                      when pause_getII6454 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13100_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"2") & \$13088\(0 to 31) & eclat_sub(\$13088\(80 to 95) & X"000" & X"1") & \$13100_v\ & \$13088\(128 to 135) & \$13088\(136 to 151) & \$13088\(152 to 153);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6463 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6461\ := \$ram_ptr_take\;
                        if \$v6461\(0) = '1' then
                          state_var6675 <= q_wait6460;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(64 to 95);
                          state_var6675 <= pause_setI6458;
                        end if;
                      when pause_getII6467 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6465\ := \$ram_ptr_take\;
                        if \$v6465\(0) = '1' then
                          state_var6675 <= q_wait6464;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6462;
                        end if;
                      when pause_getII6471 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13146_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"2") & \$13134\(0 to 31) & eclat_sub(\$13134\(80 to 95) & X"000" & X"1") & \$13146_v\ & \$13134\(128 to 135) & \$13134\(136 to 151) & \$13134\(152 to 153);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6480 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6478\ := \$ram_ptr_take\;
                        if \$v6478\(0) = '1' then
                          state_var6675 <= q_wait6477;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(64 to 95);
                          state_var6675 <= pause_setI6475;
                        end if;
                      when pause_getII6484 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6482\ := \$ram_ptr_take\;
                        if \$v6482\(0) = '1' then
                          state_var6675 <= q_wait6481;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6479;
                        end if;
                      when pause_getII6488 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6486\ := \$ram_ptr_take\;
                        if \$v6486\(0) = '1' then
                          state_var6675 <= q_wait6485;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6483;
                        end if;
                      when pause_getII6492 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13204_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"2") & \$13192\(0 to 31) & eclat_sub(\$13192\(80 to 95) & X"000" & X"1") & \$13204_v\ & \$13192\(128 to 135) & \$13192\(136 to 151) & \$13192\(152 to 153);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6501 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6499\ := \$ram_ptr_take\;
                        if \$v6499\(0) = '1' then
                          state_var6675 <= q_wait6498;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(64 to 95);
                          state_var6675 <= pause_setI6496;
                        end if;
                      when pause_getII6505 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6503\ := \$ram_ptr_take\;
                        if \$v6503\(0) = '1' then
                          state_var6675 <= q_wait6502;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6500;
                        end if;
                      when pause_getII6509 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6507\ := \$ram_ptr_take\;
                        if \$v6507\(0) = '1' then
                          state_var6675 <= q_wait6506;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6504;
                        end if;
                      when pause_getII6513 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6511\ := \$ram_ptr_take\;
                        if \$v6511\(0) = '1' then
                          state_var6675 <= q_wait6510;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6508;
                        end if;
                      when pause_getII6525 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13278_f0\ := \$ram_value\;
                        \$v6523\ := \$ram_ptr_take\;
                        if \$v6523\(0) = '1' then
                          state_var6675 <= q_wait6522;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & X"000" & X"0") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= eclat_add(\$13278_f0\(0 to 30) & \$12246_argument1\) & eclat_true;
                          state_var6675 <= pause_setI6520;
                        end if;
                      when pause_getII6533 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12455\ := \$ram_value\;
                        \$v6531\ := \$ram_ptr_take\;
                        if \$v6531\(0) = '1' then
                          state_var6675 <= q_wait6530;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_sub(\$12421_w594_arg\(16 to 31) & \$12421_w594_arg\(32 to 47)) & \$12421_w594_arg\(48 to 63)) & \$12421_w594_arg\(0 to 15))));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12455\;
                          state_var6675 <= pause_setI6528;
                        end if;
                      when pause_getII6538 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12426\ := \$ram_value\;
                        result5714 := eclat_resize(\$12426\(0 to 30),16) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(16 to 47) & eclat_sub(eclat_add(\$12190\(96 to 103) & eclat_resize(\$12246_argument1\,8)) & "00000001") & \$12190\(104 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6546 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12490_v\ := \$ram_value\;
                        \$v6544\ := \$ram_ptr_take\;
                        if \$v6544\(0) = '1' then
                          state_var6675 <= q_wait6543;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12474_fill595_arg\(48 to 78),16) & \$12474_fill595_arg\(0 to 15)) & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12490_v\;
                          state_var6675 <= pause_setI6541;
                        end if;
                      when pause_getII6560 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12528_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"3") & \$12528_v\ & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6564 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12524\ := \$ram_value\;
                        \$v6562\ := \$ram_ptr_take\;
                        if \$v6562\(0) = '1' then
                          state_var6675 <= q_wait6561;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12524\(0 to 30),16) & eclat_resize(\$12248_argument2\,16)) & X"000" & X"1")));
                          state_var6675 <= pause_getI6559;
                        end if;
                      when pause_getII6568 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12544_v\ := \$ram_value\;
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"3") & \$12544_v\ & eclat_add(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6572 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12540\ := \$ram_value\;
                        \$v6570\ := \$ram_ptr_take\;
                        if \$v6570\(0) = '1' then
                          state_var6675 <= q_wait6569;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12540\(0 to 30),16) & eclat_resize(\$12248_argument2\,16)) & X"000" & X"1")));
                          state_var6675 <= pause_getI6567;
                        end if;
                      when pause_getII6584 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12580_v\ := \$ram_value\;
                        \$v6582\ := \$ram_ptr_take\;
                        if \$v6582\(0) = '1' then
                          state_var6675 <= q_wait6581;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12564_fill596_arg\(48 to 78),16) & \$12564_fill596_arg\(0 to 15)) & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12580_v\;
                          state_var6675 <= pause_setI6579;
                        end if;
                      when pause_getII6597 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12376_v\ := \$ram_value\;
                        \$v6595\ := \$ram_ptr_take\;
                        if \$v6595\(0) = '1' then
                          state_var6675 <= q_wait6594;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12265_w0591_arg\(64 to 94),16) & eclat_sub(eclat_add(\$12265_w0591_arg\(0 to 15) & eclat_mult(X"000" & X"2" & \$12265_w0591_arg\(32 to 47))) & X"000" & X"1")) & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12376_v\;
                          state_var6675 <= pause_setI6592;
                        end if;
                      when pause_getII6606 =>
                        \$code_ptr_take\(0) := '0';
                        \$12321\ := \$code_value\;
                        \$v6604\ := \$ram_ptr_take\;
                        if \$v6604\(0) = '1' then
                          state_var6675 <= q_wait6603;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12267_w1592_arg\(48 to 78),16) & eclat_mult(X"000" & X"2" & \$12267_w1592_arg\(0 to 15))) & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= eclat_resize(eclat_add(eclat_add(\$12267_w1592_arg\(16 to 31) & X"000" & X"2") & eclat_resize(\$12321\,16)),31) & eclat_true;
                          state_var6675 <= pause_setI6601;
                        end if;
                      when pause_getII6633 =>
                        \$code_ptr_take\(0) := '0';
                        \$12253\ := \$code_value\;
                        eclat_print_int(\$12253\);
                        
                        eclat_print_newline(eclat_unit);
                        
                        result5714 := \$12190\(0 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_getII6638 =>
                        \$code_ptr_take\(0) := '0';
                        \$12250_argument3\ := \$code_value\;
                        \$v6636\ := eclat_resize(\$12243\,8);
                        case \$v6636\ is
                        when "00101100" =>
                          \$v6631\ := eclat_gt(eclat_resize(\$12248_argument2\,16) & X"000" & X"0");
                          if \$v6631\(0) = '1' then
                            \$v6630\ := \$ram_ptr_take\;
                            if \$v6630\(0) = '1' then
                              state_var6675 <= q_wait6629;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$12190\(16 to 47);
                              state_var6675 <= pause_setI6627;
                            end if;
                          else
                            \$12256_sp\ := \$12190\(48 to 63);
                            \$12199_make_block525_id\ := "000001010011";
                            \$12199_make_block525_arg\ := \$12256_sp\ & \$12190\(16 to 47) & \$12190\(64 to 95) & "11110111" & eclat_add(eclat_sub(eclat_mult(X"000" & X"2" & eclat_resize(\$12246_argument1\,16)) & X"000" & X"1") & eclat_resize(\$12248_argument2\,16));
                            state_var6675 <= \$12199_make_block525\;
                          end if;
                        when others =>
                          eclat_print_string(of_string("unknown opcode : "));
                          
                          \$v6635\ := \$code_ptr_take\;
                          if \$v6635\(0) = '1' then
                            state_var6675 <= q_wait6634;
                          else
                            \$code_ptr_take\(0) := '1';
                            \$code_ptr\ <= to_integer(unsigned(\$12190\(0 to 15)));
                            state_var6675 <= pause_getI6632;
                          end if;
                        end case;
                      when pause_getII6643 =>
                        \$code_ptr_take\(0) := '0';
                        \$12248_argument2\ := \$code_value\;
                        \$v6641\ := eclat_resize(\$12243\,8);
                        case \$v6641\ is
                        when "00100100" =>
                          \$12421_w594_arg\ := X"000" & X"1" & \$12190\(48 to 63) & eclat_resize(\$12246_argument1\,16) & eclat_resize(\$12248_argument2\,16);
                          state_var6675 <= \$12421_w594\;
                        when "00101011" =>
                          \$v6558\ := eclat_gt(eclat_resize(\$12246_argument1\,16) & X"000" & X"0");
                          if \$v6558\(0) = '1' then
                            \$v6557\ := \$ram_ptr_take\;
                            if \$v6557\(0) = '1' then
                              state_var6675 <= q_wait6556;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$12190\(16 to 47);
                              state_var6675 <= pause_setI6554;
                            end if;
                          else
                            \$12465_sp\ := \$12190\(48 to 63);
                            \$12199_make_block525_id\ := "000001000111";
                            \$12199_make_block525_arg\ := \$12465_sp\ & \$12190\(16 to 47) & \$12190\(64 to 95) & "11110111" & eclat_add(eclat_resize(\$12246_argument1\,16) & X"000" & X"1");
                            state_var6675 <= \$12199_make_block525\;
                          end if;
                        when "00110111" =>
                          \$v6566\ := \$ram_ptr_take\;
                          if \$v6566\(0) = '1' then
                            state_var6675 <= q_wait6565;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_add(X"3e80" & eclat_resize(\$12246_argument1\,16))));
                            state_var6675 <= pause_getI6563;
                          end if;
                        when "00111000" =>
                          \$v6578\ := \$ram_ptr_take\;
                          if \$v6578\(0) = '1' then
                            state_var6675 <= q_wait6577;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(16 to 47);
                            state_var6675 <= pause_setI6575;
                          end if;
                        when "00111110" =>
                          \$12199_make_block525_id\ := "000001001001";
                          \$12199_make_block525_arg\ := \$12190\(48 to 63) & \$12190\(16 to 47) & \$12190\(64 to 95) & eclat_resize(\$12248_argument2\,8) & eclat_resize(\$12246_argument1\,16);
                          state_var6675 <= \$12199_make_block525\;
                        when "10000011" =>
                          \$12245_compbranch590_arg\ := X"0000000" & X"0" & \$12246_argument1\ & \$12248_argument2\ & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          state_var6675 <= \$12245_compbranch590\;
                        when "10000100" =>
                          \$12245_compbranch590_arg\ := X"0000000" & X"1" & \$12246_argument1\ & \$12248_argument2\ & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          state_var6675 <= \$12245_compbranch590\;
                        when "10000101" =>
                          \$12245_compbranch590_arg\ := X"0000000" & X"2" & \$12246_argument1\ & \$12248_argument2\ & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          state_var6675 <= \$12245_compbranch590\;
                        when "10000110" =>
                          \$12245_compbranch590_arg\ := X"0000000" & X"3" & \$12246_argument1\ & \$12248_argument2\ & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          state_var6675 <= \$12245_compbranch590\;
                        when "10000111" =>
                          \$12245_compbranch590_arg\ := X"0000000" & X"4" & \$12246_argument1\ & \$12248_argument2\ & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          state_var6675 <= \$12245_compbranch590\;
                        when "10001000" =>
                          \$12245_compbranch590_arg\ := X"0000000" & X"5" & \$12246_argument1\ & \$12248_argument2\ & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          state_var6675 <= \$12245_compbranch590\;
                        when others =>
                          \$v6640\ := \$code_ptr_take\;
                          if \$v6640\(0) = '1' then
                            state_var6675 <= q_wait6639;
                          else
                            \$code_ptr_take\(0) := '1';
                            \$code_ptr\ <= to_integer(unsigned(eclat_add(\$12190\(0 to 15) & X"000" & X"3")));
                            state_var6675 <= pause_getI6637;
                          end if;
                        end case;
                      when pause_getII6648 =>
                        \$code_ptr_take\(0) := '0';
                        \$12246_argument1\ := \$code_value\;
                        \$v6646\ := eclat_resize(\$12243\,8);
                        case \$v6646\ is
                        when "00001000" =>
                          \$v6282\ := \$ram_ptr_take\;
                          if \$v6282\(0) = '1' then
                            state_var6675 <= q_wait6281;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & eclat_resize(\$12246_argument1\,16)) & X"000" & X"1")));
                            state_var6675 <= pause_getI6279;
                          end if;
                        when "00010010" =>
                          \$v6290\ := \$ram_ptr_take\;
                          if \$v6290\(0) = '1' then
                            state_var6675 <= q_wait6289;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(16 to 47);
                            state_var6675 <= pause_setI6287;
                          end if;
                        when "00010011" =>
                          result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"2") & \$12190\(16 to 47) & eclat_sub(\$12190\(48 to 63) & eclat_resize(\$12246_argument1\,16)) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        when "00010100" =>
                          \$v6294\ := \$ram_ptr_take\;
                          if \$v6294\(0) = '1' then
                            state_var6675 <= q_wait6293;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & eclat_resize(\$12246_argument1\,16))));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(16 to 47);
                            state_var6675 <= pause_setI6291;
                          end if;
                        when "00011001" =>
                          \$v6298\ := \$ram_ptr_take\;
                          if \$v6298\(0) = '1' then
                            state_var6675 <= q_wait6297;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(64 to 94),16) & eclat_sub(eclat_resize(\$12246_argument1\,16) & X"000" & X"1")) & X"000" & X"1")));
                            state_var6675 <= pause_getI6295;
                          end if;
                        when "00011110" =>
                          \$v6306\ := \$ram_ptr_take\;
                          if \$v6306\(0) = '1' then
                            state_var6675 <= q_wait6305;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(16 to 47);
                            state_var6675 <= pause_setI6303;
                          end if;
                        when "00011111" =>
                          \$v6318\ := \$ram_ptr_take\;
                          if \$v6318\(0) = '1' then
                            state_var6675 <= q_wait6317;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= eclat_resize(\$12190\(96 to 103),31) & eclat_true;
                            state_var6675 <= pause_setI6315;
                          end if;
                        when "00100000" =>
                          \$v6322\ := \$ram_ptr_take\;
                          if \$v6322\(0) = '1' then
                            state_var6675 <= q_wait6321;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & X"000" & X"0") & X"000" & X"1")));
                            state_var6675 <= pause_getI6319;
                          end if;
                        when "00100101" =>
                          \$12235_apply579_arg\ := eclat_true & eclat_false & eclat_false & \$12190\(96 to 103) & eclat_true & eclat_resize(\$12246_argument1\,16) & X"000" & X"1" & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(120 to 121) & \$12190\(64 to 95) & \$12190\(96 to 103) & \$12190\(104 to 119);
                          state_var6675 <= \$12235_apply579\;
                        when "00100110" =>
                          \$12235_apply579_arg\ := eclat_true & eclat_true & eclat_false & eclat_add(\$12190\(96 to 103) & "00000001") & eclat_true & eclat_resize(\$12246_argument1\,16) & X"000" & X"2" & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(120 to 121) & \$12190\(64 to 95) & \$12190\(96 to 103) & \$12190\(104 to 119);
                          state_var6675 <= \$12235_apply579\;
                        when "00100111" =>
                          \$12235_apply579_arg\ := eclat_true & eclat_true & eclat_true & eclat_add(\$12190\(96 to 103) & "00000010") & eclat_true & eclat_resize(\$12246_argument1\,16) & X"000" & X"3" & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(120 to 121) & \$12190\(64 to 95) & \$12190\(96 to 103) & \$12190\(104 to 119);
                          state_var6675 <= \$12235_apply579\;
                        when "00101000" =>
                          \$v6339\ := eclat_gt(\$12190\(96 to 103) & "00000000");
                          if \$v6339\(0) = '1' then
                            \$v6326\ := \$ram_ptr_take\;
                            if \$v6326\(0) = '1' then
                              state_var6675 <= q_wait6325;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & X"000" & X"0") & X"000" & X"1")));
                              state_var6675 <= pause_getI6323;
                            end if;
                          else
                            \$v6338\ := \$ram_ptr_take\;
                            if \$v6338\(0) = '1' then
                              state_var6675 <= q_wait6337;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & eclat_resize(\$12246_argument1\,16)) & X"000" & X"1")));
                              state_var6675 <= pause_getI6335;
                            end if;
                          end if;
                        when "00101010" =>
                          \$v6369\ := eclat_ge(\$12190\(96 to 103) & eclat_resize(\$12246_argument1\,8));
                          if \$v6369\(0) = '1' then
                            result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"2") & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 95) & eclat_sub(\$12190\(96 to 103) & eclat_resize(\$12246_argument1\,8)) & \$12190\(104 to 119) & \$12190\(120 to 121);
                            rdy5715 := eclat_true;
                            state_var6675 <= compute5716;
                          else
                            \$12199_make_block525_id\ := "000000111000";
                            \$12199_make_block525_arg\ := \$12190\(48 to 63) & \$12190\(16 to 47) & \$12190\(64 to 95) & "11110111" & eclat_resize(eclat_add(\$12190\(96 to 103) & "00000011"),16);
                            state_var6675 <= \$12199_make_block525\;
                          end if;
                        when "00110000" =>
                          \$12236_offsetclosure_n580_arg\ := eclat_add(\$12190\(0 to 15) & X"000" & X"2") & \$12190\(48 to 63) & eclat_resize(\$12246_argument1\,16) & \$12190\(64 to 119) & \$12190\(120 to 121) & \$12190\(64 to 95);
                          state_var6675 <= \$12236_offsetclosure_n580\;
                        when "00110100" =>
                          \$v6373\ := \$ram_ptr_take\;
                          if \$v6373\(0) = '1' then
                            state_var6675 <= q_wait6372;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(16 to 47);
                            state_var6675 <= pause_setI6370;
                          end if;
                        when "00110101" =>
                          \$v6377\ := \$ram_ptr_take\;
                          if \$v6377\(0) = '1' then
                            state_var6675 <= q_wait6376;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_add(X"3e80" & eclat_resize(\$12246_argument1\,16))));
                            state_var6675 <= pause_getI6374;
                          end if;
                        when "00110110" =>
                          \$v6385\ := \$ram_ptr_take\;
                          if \$v6385\(0) = '1' then
                            state_var6675 <= q_wait6384;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(16 to 47);
                            state_var6675 <= pause_setI6382;
                          end if;
                        when "00111001" =>
                          \$v6389\ := \$ram_ptr_take\;
                          if \$v6389\(0) = '1' then
                            state_var6675 <= q_wait6388;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(X"3e80" & eclat_resize(\$12246_argument1\,16))));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(16 to 47);
                            state_var6675 <= pause_setI6386;
                          end if;
                        when "00111011" =>
                          \$12240_make_block_n587_arg\ := eclat_add(\$12190\(0 to 15) & X"000" & X"2") & \$12190\(48 to 63) & eclat_false & eclat_false & eclat_false & \$12246_argument1\ & X"000" & X"0" & \$12190\(16 to 47) & \$12190\(120 to 121) & \$12190\(64 to 95) & \$12190\(96 to 103) & \$12190\(104 to 119);
                          state_var6675 <= \$12240_make_block_n587\;
                        when "00111101" =>
                          \$v6393\ := \$ram_ptr_take\;
                          if \$v6393\(0) = '1' then
                            state_var6675 <= q_wait6392;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(16 to 47);
                            state_var6675 <= pause_setI6390;
                          end if;
                        when "00111111" =>
                          \$12240_make_block_n587_arg\ := eclat_add(\$12190\(0 to 15) & X"000" & X"2") & \$12190\(48 to 63) & eclat_true & eclat_false & eclat_false & \$12246_argument1\ & X"000" & X"1" & \$12190\(16 to 47) & \$12190\(120 to 121) & \$12190\(64 to 95) & \$12190\(96 to 103) & \$12190\(104 to 119);
                          state_var6675 <= \$12240_make_block_n587\;
                        when "01000000" =>
                          \$12240_make_block_n587_arg\ := eclat_add(\$12190\(0 to 15) & X"000" & X"2") & \$12190\(48 to 63) & eclat_true & eclat_true & eclat_false & \$12246_argument1\ & X"000" & X"2" & \$12190\(16 to 47) & \$12190\(120 to 121) & \$12190\(64 to 95) & \$12190\(96 to 103) & \$12190\(104 to 119);
                          state_var6675 <= \$12240_make_block_n587\;
                        when "01000001" =>
                          \$12240_make_block_n587_arg\ := eclat_add(\$12190\(0 to 15) & X"000" & X"2") & \$12190\(48 to 63) & eclat_true & eclat_true & eclat_true & \$12246_argument1\ & X"000" & X"3" & \$12190\(16 to 47) & \$12190\(120 to 121) & \$12190\(64 to 95) & \$12190\(96 to 103) & \$12190\(104 to 119);
                          state_var6675 <= \$12240_make_block_n587\;
                        when "01000010" =>
                          eclat_print_string(of_string("fatal error: "));
                          
                          eclat_print_string(of_string("unsupported instruction SETFLOATFIELD"));
                          
                          eclat_print_newline(eclat_unit);
                          
                          state_var6675 <= \$12909_forever611\;
                        when "01000111" =>
                          assert eclat_not(""&\$12190\(47)) = eclat_true report "assertion failed" severity error;
                          
                          \$v6397\ := \$ram_ptr_take\;
                          if \$v6397\(0) = '1' then
                            state_var6675 <= q_wait6396;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & eclat_resize(\$12246_argument1\,16)) & X"000" & X"1")));
                            state_var6675 <= pause_getI6394;
                          end if;
                        when "01001101" =>
                          \$v6405\ := \$ram_ptr_take\;
                          if \$v6405\(0) = '1' then
                            state_var6675 <= q_wait6404;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12190\(48 to 63) & X"000" & X"1")));
                            state_var6675 <= pause_getI6402;
                          end if;
                        when "01001110" =>
                          eclat_print_string(of_string("fatal error: "));
                          
                          eclat_print_string(of_string("unsupported instruction SETFLOATFIELD"));
                          
                          eclat_print_newline(eclat_unit);
                          
                          state_var6675 <= \$12946_forever611\;
                        when "01010111" =>
                          \$v6414\ := ""&\$12190\(47);
                          if \$v6414\(0) = '1' then
                            \$12953_ofs\ := eclat_resize(\$12190\(16 to 46),16);
                            \$v6409\ := \$code_ptr_take\;
                            if \$v6409\(0) = '1' then
                              state_var6675 <= q_wait6408;
                            else
                              \$code_ptr_take\(0) := '1';
                              \$code_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(\$12190\(0 to 15) & X"000" & X"2") & \$12953_ofs\)));
                              state_var6675 <= pause_getI6406;
                            end if;
                          else
                            \$v6413\ := \$ram_ptr_take\;
                            if \$v6413\(0) = '1' then
                              state_var6675 <= q_wait6412;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$12190\(16 to 46),16)));
                              state_var6675 <= pause_getI6410;
                            end if;
                          end if;
                        when "01010100" =>
                          result5714 := eclat_add(eclat_add(\$12190\(0 to 15) & X"000" & X"1") & eclat_resize(\$12246_argument1\,16)) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        when "01011001" =>
                          \$v6430\ := \$ram_ptr_take\;
                          if \$v6430\(0) = '1' then
                            state_var6675 <= q_wait6429;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= eclat_resize(\$12190\(96 to 103),31) & eclat_true;
                            state_var6675 <= pause_setI6427;
                          end if;
                        when "01011100" =>
                          result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 95) & \$12190\(96 to 103) & \$12190\(104 to 119) & \$12190\(120 to 121);
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        when "01011101" =>
                          \$v6439\ := \$ram_ptr_take\;
                          if \$v6439\(0) = '1' then
                            state_var6675 <= q_wait6438;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(64 to 95);
                            state_var6675 <= pause_setI6436;
                          end if;
                        when "01011110" =>
                          \$v6452\ := \$ram_ptr_take\;
                          if \$v6452\(0) = '1' then
                            state_var6675 <= q_wait6451;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12190\(48 to 63) & X"000" & X"1")));
                            state_var6675 <= pause_getI6449;
                          end if;
                        when "01011111" =>
                          \$v6469\ := \$ram_ptr_take\;
                          if \$v6469\(0) = '1' then
                            state_var6675 <= q_wait6468;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12190\(48 to 63) & X"000" & X"1")));
                            state_var6675 <= pause_getI6466;
                          end if;
                        when "01100000" =>
                          \$v6490\ := \$ram_ptr_take\;
                          if \$v6490\(0) = '1' then
                            state_var6675 <= q_wait6489;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12190\(48 to 63) & X"000" & X"1")));
                            state_var6675 <= pause_getI6487;
                          end if;
                        when "01100001" =>
                          \$v6515\ := \$ram_ptr_take\;
                          if \$v6515\(0) = '1' then
                            state_var6675 <= q_wait6514;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12190\(48 to 63) & X"000" & X"1")));
                            state_var6675 <= pause_getI6512;
                          end if;
                        when "01100010" =>
                          eclat_print_string(of_string("fatal error: "));
                          
                          eclat_print_string(of_string("unsupported instruction CALLN"));
                          
                          eclat_print_newline(eclat_unit);
                          
                          state_var6675 <= \$13261_forever611\;
                        when "01100111" =>
                          result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"2") & \$12246_argument1\ & eclat_true & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        when "01101100" =>
                          \$v6519\ := \$ram_ptr_take\;
                          if \$v6519\(0) = '1' then
                            state_var6675 <= q_wait6518;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(16 to 47);
                            state_var6675 <= pause_setI6516;
                          end if;
                        when "01111111" =>
                          result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"2") & eclat_add(\$12190\(16 to 46) & \$12246_argument1\) & eclat_true & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        when "10000000" =>
                          \$v6527\ := \$ram_ptr_take\;
                          if \$v6527\(0) = '1' then
                            state_var6675 <= q_wait6526;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & X"000" & X"0") & X"000" & X"1")));
                            state_var6675 <= pause_getI6524;
                          end if;
                        when "10001011" =>
                          \$12245_compbranch590_arg\ := X"0000000" & X"2" & \$12246_argument1\ & \$12190\(16 to 46) & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          state_var6675 <= \$12245_compbranch590\;
                        when "10001100" =>
                          \$12245_compbranch590_arg\ := X"0000000" & X"5" & \$12246_argument1\ & \$12190\(16 to 46) & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          state_var6675 <= \$12245_compbranch590\;
                        when others =>
                          \$v6645\ := \$code_ptr_take\;
                          if \$v6645\(0) = '1' then
                            state_var6675 <= q_wait6644;
                          else
                            \$code_ptr_take\(0) := '1';
                            \$code_ptr\ <= to_integer(unsigned(eclat_add(\$12190\(0 to 15) & X"000" & X"2")));
                            state_var6675 <= pause_getI6642;
                          end if;
                        end case;
                      when pause_getII6653 =>
                        \$code_ptr_take\(0) := '0';
                        \$12243\ := \$code_value\;
                        \$v6651\ := eclat_resize(\$12243\,8);
                        case \$v6651\ is
                        when "00000000" =>
                          \$v5977\ := \$ram_ptr_take\;
                          if \$v5977\(0) = '1' then
                            state_var6675 <= q_wait5976;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"0") & X"000" & X"1")));
                            state_var6675 <= pause_getI5974;
                          end if;
                        when "00000001" =>
                          \$v5981\ := \$ram_ptr_take\;
                          if \$v5981\(0) = '1' then
                            state_var6675 <= q_wait5980;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1")));
                            state_var6675 <= pause_getI5978;
                          end if;
                        when "00000010" =>
                          \$v5985\ := \$ram_ptr_take\;
                          if \$v5985\(0) = '1' then
                            state_var6675 <= q_wait5984;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"2") & X"000" & X"1")));
                            state_var6675 <= pause_getI5982;
                          end if;
                        when "00000011" =>
                          \$v5989\ := \$ram_ptr_take\;
                          if \$v5989\(0) = '1' then
                            state_var6675 <= q_wait5988;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"3") & X"000" & X"1")));
                            state_var6675 <= pause_getI5986;
                          end if;
                        when "00000100" =>
                          \$v5993\ := \$ram_ptr_take\;
                          if \$v5993\(0) = '1' then
                            state_var6675 <= q_wait5992;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"4") & X"000" & X"1")));
                            state_var6675 <= pause_getI5990;
                          end if;
                        when "00000101" =>
                          \$v5997\ := \$ram_ptr_take\;
                          if \$v5997\(0) = '1' then
                            state_var6675 <= q_wait5996;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"5") & X"000" & X"1")));
                            state_var6675 <= pause_getI5994;
                          end if;
                        when "00000110" =>
                          \$v6001\ := \$ram_ptr_take\;
                          if \$v6001\(0) = '1' then
                            state_var6675 <= q_wait6000;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"6") & X"000" & X"1")));
                            state_var6675 <= pause_getI5998;
                          end if;
                        when "00000111" =>
                          \$v6005\ := \$ram_ptr_take\;
                          if \$v6005\(0) = '1' then
                            state_var6675 <= q_wait6004;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"7") & X"000" & X"1")));
                            state_var6675 <= pause_getI6002;
                          end if;
                        when "00001001" =>
                          \$v6009\ := \$ram_ptr_take\;
                          if \$v6009\(0) = '1' then
                            state_var6675 <= q_wait6008;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(16 to 47);
                            state_var6675 <= pause_setI6006;
                          end if;
                        when "00001010" =>
                          \$v6013\ := \$ram_ptr_take\;
                          if \$v6013\(0) = '1' then
                            state_var6675 <= q_wait6012;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(16 to 47);
                            state_var6675 <= pause_setI6010;
                          end if;
                        when "00001011" =>
                          \$v6021\ := \$ram_ptr_take\;
                          if \$v6021\(0) = '1' then
                            state_var6675 <= q_wait6020;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(16 to 47);
                            state_var6675 <= pause_setI6018;
                          end if;
                        when "00001100" =>
                          \$v6029\ := \$ram_ptr_take\;
                          if \$v6029\(0) = '1' then
                            state_var6675 <= q_wait6028;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(16 to 47);
                            state_var6675 <= pause_setI6026;
                          end if;
                        when "00001101" =>
                          \$v6037\ := \$ram_ptr_take\;
                          if \$v6037\(0) = '1' then
                            state_var6675 <= q_wait6036;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(16 to 47);
                            state_var6675 <= pause_setI6034;
                          end if;
                        when "00001110" =>
                          \$v6045\ := \$ram_ptr_take\;
                          if \$v6045\(0) = '1' then
                            state_var6675 <= q_wait6044;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(16 to 47);
                            state_var6675 <= pause_setI6042;
                          end if;
                        when "00001111" =>
                          \$v6053\ := \$ram_ptr_take\;
                          if \$v6053\(0) = '1' then
                            state_var6675 <= q_wait6052;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(16 to 47);
                            state_var6675 <= pause_setI6050;
                          end if;
                        when "00010000" =>
                          \$v6061\ := \$ram_ptr_take\;
                          if \$v6061\(0) = '1' then
                            state_var6675 <= q_wait6060;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(16 to 47);
                            state_var6675 <= pause_setI6058;
                          end if;
                        when "00010001" =>
                          \$v6069\ := \$ram_ptr_take\;
                          if \$v6069\(0) = '1' then
                            state_var6675 <= q_wait6068;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(16 to 47);
                            state_var6675 <= pause_setI6066;
                          end if;
                        when "00010101" =>
                          \$v6073\ := \$ram_ptr_take\;
                          if \$v6073\(0) = '1' then
                            state_var6675 <= q_wait6072;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(64 to 94),16) & eclat_sub(X"000" & X"1" & X"000" & X"1")) & X"000" & X"1")));
                            state_var6675 <= pause_getI6070;
                          end if;
                        when "00010110" =>
                          \$v6077\ := \$ram_ptr_take\;
                          if \$v6077\(0) = '1' then
                            state_var6675 <= q_wait6076;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(64 to 94),16) & eclat_sub(X"000" & X"2" & X"000" & X"1")) & X"000" & X"1")));
                            state_var6675 <= pause_getI6074;
                          end if;
                        when "00010111" =>
                          \$v6081\ := \$ram_ptr_take\;
                          if \$v6081\(0) = '1' then
                            state_var6675 <= q_wait6080;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(64 to 94),16) & eclat_sub(X"000" & X"3" & X"000" & X"1")) & X"000" & X"1")));
                            state_var6675 <= pause_getI6078;
                          end if;
                        when "00011000" =>
                          \$v6085\ := \$ram_ptr_take\;
                          if \$v6085\(0) = '1' then
                            state_var6675 <= q_wait6084;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(64 to 94),16) & eclat_sub(X"000" & X"4" & X"000" & X"1")) & X"000" & X"1")));
                            state_var6675 <= pause_getI6082;
                          end if;
                        when "00011010" =>
                          \$v6093\ := \$ram_ptr_take\;
                          if \$v6093\(0) = '1' then
                            state_var6675 <= q_wait6092;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(16 to 47);
                            state_var6675 <= pause_setI6090;
                          end if;
                        when "00011011" =>
                          \$v6101\ := \$ram_ptr_take\;
                          if \$v6101\(0) = '1' then
                            state_var6675 <= q_wait6100;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(16 to 47);
                            state_var6675 <= pause_setI6098;
                          end if;
                        when "00011100" =>
                          \$v6109\ := \$ram_ptr_take\;
                          if \$v6109\(0) = '1' then
                            state_var6675 <= q_wait6108;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(16 to 47);
                            state_var6675 <= pause_setI6106;
                          end if;
                        when "00011101" =>
                          \$v6117\ := \$ram_ptr_take\;
                          if \$v6117\(0) = '1' then
                            state_var6675 <= q_wait6116;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(16 to 47);
                            state_var6675 <= pause_setI6114;
                          end if;
                        when "00100001" =>
                          \$12235_apply579_arg\ := eclat_true & eclat_false & eclat_false & "00000000" & eclat_false & X"000" & X"0" & X"000" & X"0" & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(120 to 121) & \$12190\(64 to 95) & \$12190\(96 to 103) & \$12190\(104 to 119);
                          state_var6675 <= \$12235_apply579\;
                        when "00100010" =>
                          \$12235_apply579_arg\ := eclat_true & eclat_true & eclat_false & "00000001" & eclat_false & X"000" & X"0" & X"000" & X"0" & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(120 to 121) & \$12190\(64 to 95) & \$12190\(96 to 103) & \$12190\(104 to 119);
                          state_var6675 <= \$12235_apply579\;
                        when "00100011" =>
                          \$12235_apply579_arg\ := eclat_true & eclat_true & eclat_true & "00000010" & eclat_false & X"000" & X"0" & X"000" & X"0" & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(120 to 121) & \$12190\(64 to 95) & \$12190\(96 to 103) & \$12190\(104 to 119);
                          state_var6675 <= \$12235_apply579\;
                        when "00101001" =>
                          \$v6134\ := \$ram_ptr_take\;
                          if \$v6134\(0) = '1' then
                            state_var6675 <= q_wait6133;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$12190\(64 to 94),16)));
                            state_var6675 <= pause_getI6131;
                          end if;
                        when "00101101" =>
                          \$12236_offsetclosure_n580_arg\ := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$12190\(48 to 63) & eclat_sub(X"000" & X"0" & X"000" & X"2") & \$12190\(64 to 119) & \$12190\(120 to 121) & \$12190\(64 to 95);
                          state_var6675 <= \$12236_offsetclosure_n580\;
                        when "00101110" =>
                          \$12236_offsetclosure_n580_arg\ := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$12190\(48 to 63) & X"000" & X"0" & \$12190\(64 to 119) & \$12190\(120 to 121) & \$12190\(64 to 95);
                          state_var6675 <= \$12236_offsetclosure_n580\;
                        when "00101111" =>
                          \$12236_offsetclosure_n580_arg\ := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$12190\(48 to 63) & X"000" & X"2" & \$12190\(64 to 119) & \$12190\(120 to 121) & \$12190\(64 to 95);
                          state_var6675 <= \$12236_offsetclosure_n580\;
                        when "00110001" =>
                          \$v6138\ := \$ram_ptr_take\;
                          if \$v6138\(0) = '1' then
                            state_var6675 <= q_wait6137;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(16 to 47);
                            state_var6675 <= pause_setI6135;
                          end if;
                        when "00110010" =>
                          \$v6142\ := \$ram_ptr_take\;
                          if \$v6142\(0) = '1' then
                            state_var6675 <= q_wait6141;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(16 to 47);
                            state_var6675 <= pause_setI6139;
                          end if;
                        when "00110011" =>
                          \$v6146\ := \$ram_ptr_take\;
                          if \$v6146\(0) = '1' then
                            state_var6675 <= q_wait6145;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(16 to 47);
                            state_var6675 <= pause_setI6143;
                          end if;
                        when "00111010" =>
                          \$12240_make_block_n587_arg\ := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$12190\(48 to 63) & eclat_false & eclat_false & eclat_false & "000"& X"000000" & X"0" & X"000" & X"0" & \$12190\(16 to 47) & \$12190\(120 to 121) & \$12190\(64 to 95) & \$12190\(96 to 103) & \$12190\(104 to 119);
                          state_var6675 <= \$12240_make_block_n587\;
                        when "00111100" =>
                          \$v6150\ := \$ram_ptr_take\;
                          if \$v6150\(0) = '1' then
                            state_var6675 <= q_wait6149;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(16 to 47);
                            state_var6675 <= pause_setI6147;
                          end if;
                        when "01000011" =>
                          assert eclat_not(""&\$12190\(47)) = eclat_true report "assertion failed" severity error;
                          
                          \$v6154\ := \$ram_ptr_take\;
                          if \$v6154\(0) = '1' then
                            state_var6675 <= q_wait6153;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & X"000" & X"0") & X"000" & X"1")));
                            state_var6675 <= pause_getI6151;
                          end if;
                        when "01000100" =>
                          assert eclat_not(""&\$12190\(47)) = eclat_true report "assertion failed" severity error;
                          
                          \$v6158\ := \$ram_ptr_take\;
                          if \$v6158\(0) = '1' then
                            state_var6675 <= q_wait6157;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & X"000" & X"1") & X"000" & X"1")));
                            state_var6675 <= pause_getI6155;
                          end if;
                        when "01000101" =>
                          assert eclat_not(""&\$12190\(47)) = eclat_true report "assertion failed" severity error;
                          
                          \$v6162\ := \$ram_ptr_take\;
                          if \$v6162\(0) = '1' then
                            state_var6675 <= q_wait6161;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & X"000" & X"2") & X"000" & X"1")));
                            state_var6675 <= pause_getI6159;
                          end if;
                        when "01000110" =>
                          assert eclat_not(""&\$12190\(47)) = eclat_true report "assertion failed" severity error;
                          
                          \$v6166\ := \$ram_ptr_take\;
                          if \$v6166\(0) = '1' then
                            state_var6675 <= q_wait6165;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & X"000" & X"3") & X"000" & X"1")));
                            state_var6675 <= pause_getI6163;
                          end if;
                        when "01001001" =>
                          \$v6174\ := \$ram_ptr_take\;
                          if \$v6174\(0) = '1' then
                            state_var6675 <= q_wait6173;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12190\(48 to 63) & X"000" & X"1")));
                            state_var6675 <= pause_getI6171;
                          end if;
                        when "01001010" =>
                          \$v6182\ := \$ram_ptr_take\;
                          if \$v6182\(0) = '1' then
                            state_var6675 <= q_wait6181;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12190\(48 to 63) & X"000" & X"1")));
                            state_var6675 <= pause_getI6179;
                          end if;
                        when "01001011" =>
                          \$v6190\ := \$ram_ptr_take\;
                          if \$v6190\(0) = '1' then
                            state_var6675 <= q_wait6189;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12190\(48 to 63) & X"000" & X"1")));
                            state_var6675 <= pause_getI6187;
                          end if;
                        when "01001100" =>
                          \$v6198\ := \$ram_ptr_take\;
                          if \$v6198\(0) = '1' then
                            state_var6675 <= q_wait6197;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12190\(48 to 63) & X"000" & X"1")));
                            state_var6675 <= pause_getI6195;
                          end if;
                        when "01001111" =>
                          \$v6202\ := \$ram_ptr_take\;
                          if \$v6202\(0) = '1' then
                            state_var6675 <= q_wait6201;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$12190\(16 to 46),16)));
                            state_var6675 <= pause_getI6199;
                          end if;
                        when "01010000" =>
                          \$v6210\ := \$ram_ptr_take\;
                          if \$v6210\(0) = '1' then
                            state_var6675 <= q_wait6209;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12190\(48 to 63) & X"000" & X"1")));
                            state_var6675 <= pause_getI6207;
                          end if;
                        when "01010001" =>
                          \$v6222\ := \$ram_ptr_take\;
                          if \$v6222\(0) = '1' then
                            state_var6675 <= q_wait6221;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12190\(48 to 63) & X"000" & X"1")));
                            state_var6675 <= pause_getI6219;
                          end if;
                        when "01010010" =>
                          \$v6230\ := \$ram_ptr_take\;
                          if \$v6230\(0) = '1' then
                            state_var6675 <= q_wait6229;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12190\(48 to 63) & X"000" & X"1")));
                            state_var6675 <= pause_getI6227;
                          end if;
                        when "01010011" =>
                          \$v6242\ := \$ram_ptr_take\;
                          if \$v6242\(0) = '1' then
                            state_var6675 <= q_wait6241;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12190\(48 to 63) & X"000" & X"1")));
                            state_var6675 <= pause_getI6239;
                          end if;
                        when "01010101" =>
                          \$12241_branch_if589_arg\ := eclat_false & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          state_var6675 <= \$12241_branch_if589\;
                        when "01010110" =>
                          \$12241_branch_if589_arg\ := eclat_true & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          state_var6675 <= \$12241_branch_if589\;
                        when "01011000" =>
                          result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & 
                          eclat_if(eclat_eq(\$12190\(16 to 46) & "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        when "01011010" =>
                          \$v6246\ := \$ram_ptr_take\;
                          if \$v6246\(0) = '1' then
                            state_var6675 <= q_wait6245;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1")));
                            state_var6675 <= pause_getI6243;
                          end if;
                        when "01011011" =>
                          \$v6262\ := \$ram_ptr_take\;
                          if \$v6262\(0) = '1' then
                            state_var6675 <= q_wait6261;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12190\(104 to 119) & X"000" & X"1")));
                            state_var6675 <= pause_getI6259;
                          end if;
                        when "01100011" =>
                          result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"0" & eclat_true & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        when "01100100" =>
                          result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        when "01100101" =>
                          result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"2" & eclat_true & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        when "01100110" =>
                          result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"3" & eclat_true & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        when "01101000" =>
                          \$v6266\ := \$ram_ptr_take\;
                          if \$v6266\(0) = '1' then
                            state_var6675 <= q_wait6265;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(16 to 47);
                            state_var6675 <= pause_setI6263;
                          end if;
                        when "01101001" =>
                          \$v6270\ := \$ram_ptr_take\;
                          if \$v6270\(0) = '1' then
                            state_var6675 <= q_wait6269;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(16 to 47);
                            state_var6675 <= pause_setI6267;
                          end if;
                        when "01101010" =>
                          \$v6274\ := \$ram_ptr_take\;
                          if \$v6274\(0) = '1' then
                            state_var6675 <= q_wait6273;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(16 to 47);
                            state_var6675 <= pause_setI6271;
                          end if;
                        when "01101011" =>
                          \$v6278\ := \$ram_ptr_take\;
                          if \$v6278\(0) = '1' then
                            state_var6675 <= q_wait6277;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12190\(16 to 47);
                            state_var6675 <= pause_setI6275;
                          end if;
                        when "01101110" =>
                          \$12237_binop_int584_arg\ := X"0000000" & X"0" & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          state_var6675 <= \$12237_binop_int584\;
                        when "01101111" =>
                          \$12237_binop_int584_arg\ := X"0000000" & X"1" & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          state_var6675 <= \$12237_binop_int584\;
                        when "01110000" =>
                          \$12237_binop_int584_arg\ := X"0000000" & X"2" & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          state_var6675 <= \$12237_binop_int584\;
                        when "01110001" =>
                          \$12237_binop_int584_arg\ := X"0000000" & X"3" & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          state_var6675 <= \$12237_binop_int584\;
                        when "01110010" =>
                          \$12237_binop_int584_arg\ := X"0000000" & X"4" & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          state_var6675 <= \$12237_binop_int584\;
                        when "01110011" =>
                          \$12237_binop_int584_arg\ := X"0000000" & X"5" & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          state_var6675 <= \$12237_binop_int584\;
                        when "01110100" =>
                          \$12237_binop_int584_arg\ := X"0000000" & X"6" & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          state_var6675 <= \$12237_binop_int584\;
                        when "01110101" =>
                          \$12237_binop_int584_arg\ := X"0000000" & X"7" & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          state_var6675 <= \$12237_binop_int584\;
                        when "01110110" =>
                          \$12237_binop_int584_arg\ := X"0000000" & X"8" & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          state_var6675 <= \$12237_binop_int584\;
                        when "01110111" =>
                          \$12237_binop_int584_arg\ := X"0000000" & X"9" & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          state_var6675 <= \$12237_binop_int584\;
                        when "01111000" =>
                          \$12237_binop_int584_arg\ := X"0000000" & X"a" & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          state_var6675 <= \$12237_binop_int584\;
                        when "10000010" =>
                          eclat_print_string(of_string("fatal error: "));
                          
                          eclat_print_string(of_string("unsupported instruction GETMETHOD"));
                          
                          eclat_print_newline(eclat_unit);
                          
                          state_var6675 <= \$13928_forever611\;
                        when "10001001" =>
                          \$12237_binop_int584_arg\ := X"0000000" & X"b" & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          state_var6675 <= \$12237_binop_int584\;
                        when "10001010" =>
                          \$12237_binop_int584_arg\ := X"0000000" & X"c" & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          state_var6675 <= \$12237_binop_int584\;
                        when "10001101" =>
                          eclat_print_string(of_string("fatal error: "));
                          
                          eclat_print_string(of_string("unsupported instruction GETPUBMET"));
                          
                          eclat_print_newline(eclat_unit);
                          
                          state_var6675 <= \$13935_forever611\;
                        when "10001110" =>
                          eclat_print_string(of_string("fatal error: "));
                          
                          eclat_print_string(of_string("unsupported instruction GETDYNMET"));
                          
                          eclat_print_newline(eclat_unit);
                          
                          state_var6675 <= \$13942_forever611\;
                        when "01111001" =>
                          \$12239_binop_compare586_arg\ := X"0000000" & X"0" & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          state_var6675 <= \$12239_binop_compare586\;
                        when "01111010" =>
                          \$12239_binop_compare586_arg\ := X"0000000" & X"1" & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          state_var6675 <= \$12239_binop_compare586\;
                        when "01111011" =>
                          \$12239_binop_compare586_arg\ := X"0000000" & X"2" & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          state_var6675 <= \$12239_binop_compare586\;
                        when "01111100" =>
                          \$12239_binop_compare586_arg\ := X"0000000" & X"3" & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          state_var6675 <= \$12239_binop_compare586\;
                        when "01111101" =>
                          \$12239_binop_compare586_arg\ := X"0000000" & X"4" & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          state_var6675 <= \$12239_binop_compare586\;
                        when "01111110" =>
                          \$12239_binop_compare586_arg\ := X"0000000" & X"5" & \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          state_var6675 <= \$12239_binop_compare586\;
                        when "10000001" =>
                          result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & 
                          eclat_if(""&\$12190\(47) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        when "10001111" =>
                          eclat_print_string(of_string("STOP : "));
                          
                          result5714 := \$12190\(0 to 15) & \$12190\(16 to 47) & \$12190\(48 to 63) & \$12190\(64 to 119) & eclat_true & ""&\$12190\(121);
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        when others =>
                          \$v6650\ := \$code_ptr_take\;
                          if \$v6650\(0) = '1' then
                            state_var6675 <= q_wait6649;
                          else
                            \$code_ptr_take\(0) := '1';
                            \$code_ptr\ <= to_integer(unsigned(eclat_add(\$12190\(0 to 15) & X"000" & X"1")));
                            state_var6675 <= pause_getI6647;
                          end if;
                        end case;
                      when pause_setI5717 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII5718;
                      when pause_setI5888 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII5889;
                      when pause_setI5893 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII5894;
                      when pause_setI5898 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII5899;
                      when pause_setI5903 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII5904;
                      when pause_setI5907 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII5908;
                      when pause_setI5911 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII5912;
                      when pause_setI5946 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII5947;
                      when pause_setI5955 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII5956;
                      when pause_setI5964 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII5965;
                      when pause_setI6006 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6007;
                      when pause_setI6010 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6011;
                      when pause_setI6018 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6019;
                      when pause_setI6026 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6027;
                      when pause_setI6034 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6035;
                      when pause_setI6042 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6043;
                      when pause_setI6050 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6051;
                      when pause_setI6058 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6059;
                      when pause_setI6066 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6067;
                      when pause_setI6090 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6091;
                      when pause_setI6098 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6099;
                      when pause_setI6106 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6107;
                      when pause_setI6114 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6115;
                      when pause_setI6118 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6119;
                      when pause_setI6135 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6136;
                      when pause_setI6139 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6140;
                      when pause_setI6143 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6144;
                      when pause_setI6147 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6148;
                      when pause_setI6167 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6168;
                      when pause_setI6175 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6176;
                      when pause_setI6183 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6184;
                      when pause_setI6191 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6192;
                      when pause_setI6211 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6212;
                      when pause_setI6231 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6232;
                      when pause_setI6263 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6264;
                      when pause_setI6267 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6268;
                      when pause_setI6271 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6272;
                      when pause_setI6275 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6276;
                      when pause_setI6287 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6288;
                      when pause_setI6291 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6292;
                      when pause_setI6303 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6304;
                      when pause_setI6307 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6308;
                      when pause_setI6311 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6312;
                      when pause_setI6315 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6316;
                      when pause_setI6340 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6341;
                      when pause_setI6361 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6362;
                      when pause_setI6365 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6366;
                      when pause_setI6370 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6371;
                      when pause_setI6382 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6383;
                      when pause_setI6386 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6387;
                      when pause_setI6390 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6391;
                      when pause_setI6398 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6399;
                      when pause_setI6415 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6416;
                      when pause_setI6419 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6420;
                      when pause_setI6423 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6424;
                      when pause_setI6427 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6428;
                      when pause_setI6436 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6437;
                      when pause_setI6445 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6446;
                      when pause_setI6458 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6459;
                      when pause_setI6475 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6476;
                      when pause_setI6496 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6497;
                      when pause_setI6516 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6517;
                      when pause_setI6520 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6521;
                      when pause_setI6528 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6529;
                      when pause_setI6541 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6542;
                      when pause_setI6550 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6551;
                      when pause_setI6554 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6555;
                      when pause_setI6575 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6576;
                      when pause_setI6579 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6580;
                      when pause_setI6588 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6589;
                      when pause_setI6592 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6593;
                      when pause_setI6601 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6602;
                      when pause_setI6609 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6610;
                      when pause_setI6614 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6615;
                      when pause_setI6619 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6620;
                      when pause_setI6623 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6624;
                      when pause_setI6627 =>
                        \$ram_write_request\ <= '0';
                        state_var6675 <= pause_setII6628;
                      when pause_setII5718 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12199_make_block525_result\ := \$14250\(0 to 31) & \$14250\(32 to 63) & eclat_resize(\$14250\(64 to 79),31) & eclat_false;
                        case \$12199_make_block525_id\ is
                        when "000000001110" =>
                          \$13996\ := \$12199_make_block525_result\;
                          \$v5968\ := ""&\$12240_make_block_n587_arg\(32);
                          if \$v5968\(0) = '1' then
                            \$v5967\ := \$ram_ptr_take\;
                            if \$v5967\(0) = '1' then
                              state_var6675 <= q_wait5966;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$13996\(64 to 94),16) & X"000" & X"0") & X"000" & X"1")));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$13996\(0 to 31);
                              state_var6675 <= pause_setI5964;
                            end if;
                          else
                            \$v5963\ := ""&\$12240_make_block_n587_arg\(33);
                            if \$v5963\(0) = '1' then
                              \$v5962\ := \$ram_ptr_take\;
                              if \$v5962\(0) = '1' then
                                state_var6675 <= q_wait5961;
                              else
                                \$ram_ptr_take\(0) := '1';
                                \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12240_make_block_n587_arg\(16 to 31) & X"000" & X"1")));
                                state_var6675 <= pause_getI5959;
                              end if;
                            else
                              \$14001_sp\ := \$12240_make_block_n587_arg\(16 to 31);
                              \$v5954\ := ""&\$12240_make_block_n587_arg\(34);
                              if \$v5954\(0) = '1' then
                                \$v5953\ := \$ram_ptr_take\;
                                if \$v5953\(0) = '1' then
                                  state_var6675 <= q_wait5952;
                                else
                                  \$ram_ptr_take\(0) := '1';
                                  \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$14001_sp\ & X"000" & X"1")));
                                  state_var6675 <= pause_getI5950;
                                end if;
                              else
                                \$14002_sp\ := \$14001_sp\;
                                \$12240_make_block_n587_result\ := \$12240_make_block_n587_arg\(0 to 15) & \$13996\(64 to 95) & \$14002_sp\ & \$13996\(32 to 63) & \$12240_make_block_n587_arg\(148 to 155) & \$12240_make_block_n587_arg\(156 to 171) & \$12240_make_block_n587_arg\(114 to 115);
                                result5714 := \$12240_make_block_n587_result\;
                                rdy5715 := eclat_true;
                                state_var6675 <= compute5716;
                              end if;
                            end if;
                          end if;
                        when "000000111000" =>
                          \$12770\ := \$12199_make_block525_result\;
                          \$v6368\ := \$ram_ptr_take\;
                          if \$v6368\(0) = '1' then
                            state_var6675 <= q_wait6367;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12770\(64 to 94),16) & X"000" & X"0") & X"000" & X"1")));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= eclat_resize(eclat_sub(eclat_add(\$12190\(0 to 15) & X"000" & X"2") & X"000" & X"3"),31) & eclat_true;
                            state_var6675 <= pause_setI6365;
                          end if;
                        when "000001000111" =>
                          \$12466\ := \$12199_make_block525_result\;
                          \$v6553\ := \$ram_ptr_take\;
                          if \$v6553\(0) = '1' then
                            state_var6675 <= q_wait6552;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12466\(64 to 94),16) & X"000" & X"0") & X"000" & X"1")));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= eclat_resize(eclat_add(eclat_add(\$12190\(0 to 15) & X"000" & X"2") & eclat_resize(\$12248_argument2\,16)),31) & eclat_true;
                            state_var6675 <= pause_setI6550;
                          end if;
                        when "000001001001" =>
                          \$12556\ := \$12199_make_block525_result\;
                          \$v6591\ := \$ram_ptr_take\;
                          if \$v6591\(0) = '1' then
                            state_var6675 <= q_wait6590;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12556\(64 to 94),16) & X"000" & X"0") & X"000" & X"1")));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$12556\(0 to 31);
                            state_var6675 <= pause_setI6588;
                          end if;
                        when "000001010011" =>
                          \$12257\ := \$12199_make_block525_result\;
                          \$v6626\ := \$ram_ptr_take\;
                          if \$v6626\(0) = '1' then
                            state_var6675 <= q_wait6625;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12257\(64 to 94),16) & X"000" & X"0") & X"000" & X"1")));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= eclat_resize(eclat_add(eclat_add(\$12190\(0 to 15) & X"000" & X"3") & eclat_resize(\$12250_argument3\,16)),31) & eclat_true;
                            state_var6675 <= pause_setI6623;
                          end if;
                        when others =>
                          
                        end case;
                      when pause_setII5889 =>
                        \$ram_ptr_take\(0) := '0';
                        \$14192_sp\ := eclat_add(\$14191_sp\ & X"000" & X"1");
                        \$v5887\ := \$ram_ptr_take\;
                        if \$v5887\(0) = '1' then
                          state_var6675 <= q_wait5886;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12235_apply579_arg\(60 to 90),16) & X"000" & X"0") & X"000" & X"1")));
                          state_var6675 <= pause_getI5884;
                        end if;
                      when pause_setII5894 =>
                        \$ram_ptr_take\(0) := '0';
                        \$14191_sp\ := eclat_add(\$14190_sp\ & X"000" & X"1");
                        \$v5892\ := ""&\$12235_apply579_arg\(0);
                        if \$v5892\(0) = '1' then
                          \$v5891\ := \$ram_ptr_take\;
                          if \$v5891\(0) = '1' then
                            state_var6675 <= q_wait5890;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$14191_sp\));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$14180\(0 to 31);
                            state_var6675 <= pause_setI5888;
                          end if;
                        else
                          \$14192_sp\ := \$14191_sp\;
                          \$v5887\ := \$ram_ptr_take\;
                          if \$v5887\(0) = '1' then
                            state_var6675 <= q_wait5886;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12235_apply579_arg\(60 to 90),16) & X"000" & X"0") & X"000" & X"1")));
                            state_var6675 <= pause_getI5884;
                          end if;
                        end if;
                      when pause_setII5899 =>
                        \$ram_ptr_take\(0) := '0';
                        \$14190_sp\ := eclat_add(\$14189_sp\ & X"000" & X"1");
                        \$v5897\ := ""&\$12235_apply579_arg\(1);
                        if \$v5897\(0) = '1' then
                          \$v5896\ := \$ram_ptr_take\;
                          if \$v5896\(0) = '1' then
                            state_var6675 <= q_wait5895;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$14190_sp\));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$14183\(0 to 31);
                            state_var6675 <= pause_setI5893;
                          end if;
                        else
                          \$14191_sp\ := \$14190_sp\;
                          \$v5892\ := ""&\$12235_apply579_arg\(0);
                          if \$v5892\(0) = '1' then
                            \$v5891\ := \$ram_ptr_take\;
                            if \$v5891\(0) = '1' then
                              state_var6675 <= q_wait5890;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(\$14191_sp\));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$14180\(0 to 31);
                              state_var6675 <= pause_setI5888;
                            end if;
                          else
                            \$14192_sp\ := \$14191_sp\;
                            \$v5887\ := \$ram_ptr_take\;
                            if \$v5887\(0) = '1' then
                              state_var6675 <= q_wait5886;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12235_apply579_arg\(60 to 90),16) & X"000" & X"0") & X"000" & X"1")));
                              state_var6675 <= pause_getI5884;
                            end if;
                          end if;
                        end if;
                      when pause_setII5904 =>
                        \$ram_ptr_take\(0) := '0';
                        \$14189_sp\ := eclat_add(eclat_add(eclat_add(\$14186\(32 to 47) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1");
                        \$v5902\ := ""&\$12235_apply579_arg\(2);
                        if \$v5902\(0) = '1' then
                          \$v5901\ := \$ram_ptr_take\;
                          if \$v5901\(0) = '1' then
                            state_var6675 <= q_wait5900;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr_write\ <= to_integer(unsigned(\$14189_sp\));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$14186\(0 to 31);
                            state_var6675 <= pause_setI5898;
                          end if;
                        else
                          \$14190_sp\ := \$14189_sp\;
                          \$v5897\ := ""&\$12235_apply579_arg\(1);
                          if \$v5897\(0) = '1' then
                            \$v5896\ := \$ram_ptr_take\;
                            if \$v5896\(0) = '1' then
                              state_var6675 <= q_wait5895;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr_write\ <= to_integer(unsigned(\$14190_sp\));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$14183\(0 to 31);
                              state_var6675 <= pause_setI5893;
                            end if;
                          else
                            \$14191_sp\ := \$14190_sp\;
                            \$v5892\ := ""&\$12235_apply579_arg\(0);
                            if \$v5892\(0) = '1' then
                              \$v5891\ := \$ram_ptr_take\;
                              if \$v5891\(0) = '1' then
                                state_var6675 <= q_wait5890;
                              else
                                \$ram_ptr_take\(0) := '1';
                                \$ram_ptr_write\ <= to_integer(unsigned(\$14191_sp\));
                                \$ram_write_request\ <= '1';
                                \$ram_write\ <= \$14180\(0 to 31);
                                state_var6675 <= pause_setI5888;
                              end if;
                            else
                              \$14192_sp\ := \$14191_sp\;
                              \$v5887\ := \$ram_ptr_take\;
                              if \$v5887\(0) = '1' then
                                state_var6675 <= q_wait5886;
                              else
                                \$ram_ptr_take\(0) := '1';
                                \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12235_apply579_arg\(60 to 90),16) & X"000" & X"0") & X"000" & X"1")));
                                state_var6675 <= pause_getI5884;
                              end if;
                            end if;
                          end if;
                        end if;
                      when pause_setII5908 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v5906\ := \$ram_ptr_take\;
                        if \$v5906\(0) = '1' then
                          state_var6675 <= q_wait5905;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(\$14186\(32 to 47) & X"000" & X"1") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= eclat_resize(eclat_add(\$12235_apply579_arg\(44 to 59) & X"000" & X"1"),31) & eclat_true;
                          state_var6675 <= pause_setI5903;
                        end if;
                      when pause_setII5912 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v5910\ := \$ram_ptr_take\;
                        if \$v5910\(0) = '1' then
                          state_var6675 <= q_wait5909;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(\$14186\(32 to 47) & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12235_apply579_arg\(110 to 141);
                          state_var6675 <= pause_setI5907;
                        end if;
                      when pause_setII5947 =>
                        \$ram_ptr_take\(0) := '0';
                        \$14002_sp\ := eclat_sub(\$14001_sp\ & X"000" & X"1");
                        \$12240_make_block_n587_result\ := \$12240_make_block_n587_arg\(0 to 15) & \$13996\(64 to 95) & \$14002_sp\ & \$13996\(32 to 63) & \$12240_make_block_n587_arg\(148 to 155) & \$12240_make_block_n587_arg\(156 to 171) & \$12240_make_block_n587_arg\(114 to 115);
                        result5714 := \$12240_make_block_n587_result\;
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_setII5956 =>
                        \$ram_ptr_take\(0) := '0';
                        \$14001_sp\ := eclat_sub(\$12240_make_block_n587_arg\(16 to 31) & X"000" & X"1");
                        \$v5954\ := ""&\$12240_make_block_n587_arg\(34);
                        if \$v5954\(0) = '1' then
                          \$v5953\ := \$ram_ptr_take\;
                          if \$v5953\(0) = '1' then
                            state_var6675 <= q_wait5952;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$14001_sp\ & X"000" & X"1")));
                            state_var6675 <= pause_getI5950;
                          end if;
                        else
                          \$14002_sp\ := \$14001_sp\;
                          \$12240_make_block_n587_result\ := \$12240_make_block_n587_arg\(0 to 15) & \$13996\(64 to 95) & \$14002_sp\ & \$13996\(32 to 63) & \$12240_make_block_n587_arg\(148 to 155) & \$12240_make_block_n587_arg\(156 to 171) & \$12240_make_block_n587_arg\(114 to 115);
                          result5714 := \$12240_make_block_n587_result\;
                          rdy5715 := eclat_true;
                          state_var6675 <= compute5716;
                        end if;
                      when pause_setII5965 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v5963\ := ""&\$12240_make_block_n587_arg\(33);
                        if \$v5963\(0) = '1' then
                          \$v5962\ := \$ram_ptr_take\;
                          if \$v5962\(0) = '1' then
                            state_var6675 <= q_wait5961;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12240_make_block_n587_arg\(16 to 31) & X"000" & X"1")));
                            state_var6675 <= pause_getI5959;
                          end if;
                        else
                          \$14001_sp\ := \$12240_make_block_n587_arg\(16 to 31);
                          \$v5954\ := ""&\$12240_make_block_n587_arg\(34);
                          if \$v5954\(0) = '1' then
                            \$v5953\ := \$ram_ptr_take\;
                            if \$v5953\(0) = '1' then
                              state_var6675 <= q_wait5952;
                            else
                              \$ram_ptr_take\(0) := '1';
                              \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$14001_sp\ & X"000" & X"1")));
                              state_var6675 <= pause_getI5950;
                            end if;
                          else
                            \$14002_sp\ := \$14001_sp\;
                            \$12240_make_block_n587_result\ := \$12240_make_block_n587_arg\(0 to 15) & \$13996\(64 to 95) & \$14002_sp\ & \$13996\(32 to 63) & \$12240_make_block_n587_arg\(148 to 155) & \$12240_make_block_n587_arg\(156 to 171) & \$12240_make_block_n587_arg\(114 to 115);
                            result5714 := \$12240_make_block_n587_result\;
                            rdy5715 := eclat_true;
                            state_var6675 <= compute5716;
                          end if;
                        end if;
                      when pause_setII6007 =>
                        \$ram_ptr_take\(0) := '0';
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$12190\(16 to 47) & eclat_add(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_setII6011 =>
                        \$ram_ptr_take\(0) := '0';
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & \$12190\(16 to 47) & eclat_add(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_setII6019 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6017\ := \$ram_ptr_take\;
                        if \$v6017\(0) = '1' then
                          state_var6675 <= q_wait6016;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_add(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6014;
                        end if;
                      when pause_setII6027 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6025\ := \$ram_ptr_take\;
                        if \$v6025\(0) = '1' then
                          state_var6675 <= q_wait6024;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_add(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"2") & X"000" & X"1")));
                          state_var6675 <= pause_getI6022;
                        end if;
                      when pause_setII6035 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6033\ := \$ram_ptr_take\;
                        if \$v6033\(0) = '1' then
                          state_var6675 <= q_wait6032;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_add(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"3") & X"000" & X"1")));
                          state_var6675 <= pause_getI6030;
                        end if;
                      when pause_setII6043 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6041\ := \$ram_ptr_take\;
                        if \$v6041\(0) = '1' then
                          state_var6675 <= q_wait6040;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_add(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"4") & X"000" & X"1")));
                          state_var6675 <= pause_getI6038;
                        end if;
                      when pause_setII6051 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6049\ := \$ram_ptr_take\;
                        if \$v6049\(0) = '1' then
                          state_var6675 <= q_wait6048;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_add(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"5") & X"000" & X"1")));
                          state_var6675 <= pause_getI6046;
                        end if;
                      when pause_setII6059 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6057\ := \$ram_ptr_take\;
                        if \$v6057\(0) = '1' then
                          state_var6675 <= q_wait6056;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_add(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"6") & X"000" & X"1")));
                          state_var6675 <= pause_getI6054;
                        end if;
                      when pause_setII6067 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6065\ := \$ram_ptr_take\;
                        if \$v6065\(0) = '1' then
                          state_var6675 <= q_wait6064;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_add(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"7") & X"000" & X"1")));
                          state_var6675 <= pause_getI6062;
                        end if;
                      when pause_setII6091 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6089\ := \$ram_ptr_take\;
                        if \$v6089\(0) = '1' then
                          state_var6675 <= q_wait6088;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(64 to 94),16) & eclat_sub(X"000" & X"1" & X"000" & X"1")) & X"000" & X"1")));
                          state_var6675 <= pause_getI6086;
                        end if;
                      when pause_setII6099 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6097\ := \$ram_ptr_take\;
                        if \$v6097\(0) = '1' then
                          state_var6675 <= q_wait6096;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(64 to 94),16) & eclat_sub(X"000" & X"2" & X"000" & X"1")) & X"000" & X"1")));
                          state_var6675 <= pause_getI6094;
                        end if;
                      when pause_setII6107 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6105\ := \$ram_ptr_take\;
                        if \$v6105\(0) = '1' then
                          state_var6675 <= q_wait6104;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(64 to 94),16) & eclat_sub(X"000" & X"3" & X"000" & X"1")) & X"000" & X"1")));
                          state_var6675 <= pause_getI6102;
                        end if;
                      when pause_setII6115 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6113\ := \$ram_ptr_take\;
                        if \$v6113\(0) = '1' then
                          state_var6675 <= q_wait6112;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(64 to 94),16) & eclat_sub(X"000" & X"4" & X"000" & X"1")) & X"000" & X"1")));
                          state_var6675 <= pause_getI6110;
                        end if;
                      when pause_setII6119 =>
                        \$ram_ptr_take\(0) := '0';
                        \$13539_loop_push598_arg\ := eclat_add(\$13539_loop_push598_arg\(0 to 15) & X"000" & X"1") & eclat_add(\$13539_loop_push598_arg\(16 to 23) & "00000001") & \$13539_loop_push598_arg\(24 to 55) & \$13539_loop_push598_arg\(56 to 63);
                        state_var6675 <= \$13539_loop_push598\;
                      when pause_setII6136 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12236_offsetclosure_n580_arg\ := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & eclat_add(\$12190\(48 to 63) & X"000" & X"1") & eclat_sub(X"000" & X"0" & X"000" & X"2") & \$12190\(64 to 119) & \$12190\(120 to 121) & \$12190\(64 to 95);
                        state_var6675 <= \$12236_offsetclosure_n580\;
                      when pause_setII6140 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12236_offsetclosure_n580_arg\ := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & eclat_add(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"0" & \$12190\(64 to 119) & \$12190\(120 to 121) & \$12190\(64 to 95);
                        state_var6675 <= \$12236_offsetclosure_n580\;
                      when pause_setII6144 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12236_offsetclosure_n580_arg\ := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & eclat_add(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"2" & \$12190\(64 to 119) & \$12190\(120 to 121) & \$12190\(64 to 95);
                        state_var6675 <= \$12236_offsetclosure_n580\;
                      when pause_setII6148 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12240_make_block_n587_arg\ := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & eclat_add(\$12190\(48 to 63) & X"000" & X"1") & eclat_false & eclat_false & eclat_false & "000"& X"000000" & X"0" & X"000" & X"0" & \$12190\(16 to 47) & \$12190\(120 to 121) & \$12190\(64 to 95) & \$12190\(96 to 103) & \$12190\(104 to 119);
                        state_var6675 <= \$12240_make_block_n587\;
                      when pause_setII6168 =>
                        \$ram_ptr_take\(0) := '0';
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_setII6176 =>
                        \$ram_ptr_take\(0) := '0';
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_setII6184 =>
                        \$ram_ptr_take\(0) := '0';
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_setII6192 =>
                        \$ram_ptr_take\(0) := '0';
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_setII6212 =>
                        \$ram_ptr_take\(0) := '0';
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_setII6232 =>
                        \$ram_ptr_take\(0) := '0';
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_setII6264 =>
                        \$ram_ptr_take\(0) := '0';
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"0" & eclat_true & eclat_add(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_setII6268 =>
                        \$ram_ptr_take\(0) := '0';
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & eclat_add(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_setII6272 =>
                        \$ram_ptr_take\(0) := '0';
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"2" & eclat_true & eclat_add(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_setII6276 =>
                        \$ram_ptr_take\(0) := '0';
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"3" & eclat_true & eclat_add(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_setII6288 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6286\ := \$ram_ptr_take\;
                        if \$v6286\(0) = '1' then
                          state_var6675 <= q_wait6285;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_add(\$12190\(48 to 63) & X"000" & X"1") & eclat_resize(\$12246_argument1\,16)) & X"000" & X"1")));
                          state_var6675 <= pause_getI6283;
                        end if;
                      when pause_setII6292 =>
                        \$ram_ptr_take\(0) := '0';
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"2") & "000"& X"000000" & X"1" & eclat_true & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_setII6304 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6302\ := \$ram_ptr_take\;
                        if \$v6302\(0) = '1' then
                          state_var6675 <= q_wait6301;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(64 to 94),16) & eclat_sub(eclat_resize(\$12246_argument1\,16) & X"000" & X"1")) & X"000" & X"1")));
                          state_var6675 <= pause_getI6299;
                        end if;
                      when pause_setII6308 =>
                        \$ram_ptr_take\(0) := '0';
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"2") & \$12190\(16 to 47) & eclat_add(eclat_add(eclat_add(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_setII6312 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6310\ := \$ram_ptr_take\;
                        if \$v6310\(0) = '1' then
                          state_var6675 <= q_wait6309;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= eclat_resize(eclat_add(eclat_add(\$12190\(0 to 15) & X"000" & X"1") & eclat_resize(\$12246_argument1\,16)),31) & eclat_true;
                          state_var6675 <= pause_setI6307;
                        end if;
                      when pause_setII6316 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6314\ := \$ram_ptr_take\;
                        if \$v6314\(0) = '1' then
                          state_var6675 <= q_wait6313;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(\$12190\(48 to 63) & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(64 to 95);
                          state_var6675 <= pause_setI6311;
                        end if;
                      when pause_setII6341 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12782_w597_arg\ := eclat_add(\$12782_w597_arg\(0 to 7) & "00000001") & eclat_sub(\$12782_w597_arg\(8 to 23) & X"000" & X"1") & \$12782_w597_arg\(24 to 31) & \$12782_w597_arg\(32 to 63);
                        state_var6675 <= \$12782_w597\;
                      when pause_setII6362 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12782_w597_arg\ := "00000000" & \$12190\(48 to 63) & \$12190\(96 to 103) & \$12770\(64 to 95);
                        state_var6675 <= \$12782_w597\;
                      when pause_setII6366 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6364\ := \$ram_ptr_take\;
                        if \$v6364\(0) = '1' then
                          state_var6675 <= q_wait6363;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12770\(64 to 94),16) & X"000" & X"1") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12770\(32 to 63);
                          state_var6675 <= pause_setI6361;
                        end if;
                      when pause_setII6371 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12236_offsetclosure_n580_arg\ := eclat_add(\$12190\(0 to 15) & X"000" & X"2") & eclat_add(\$12190\(48 to 63) & X"000" & X"1") & eclat_resize(\$12246_argument1\,16) & \$12190\(64 to 119) & \$12190\(120 to 121) & \$12190\(64 to 95);
                        state_var6675 <= \$12236_offsetclosure_n580\;
                      when pause_setII6383 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6381\ := \$ram_ptr_take\;
                        if \$v6381\(0) = '1' then
                          state_var6675 <= q_wait6380;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(X"3e80" & eclat_resize(\$12246_argument1\,16))));
                          state_var6675 <= pause_getI6378;
                        end if;
                      when pause_setII6387 =>
                        \$ram_ptr_take\(0) := '0';
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"2") & "000"& X"000000" & X"1" & eclat_true & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_setII6391 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12240_make_block_n587_arg\ := eclat_add(\$12190\(0 to 15) & X"000" & X"2") & eclat_add(\$12190\(48 to 63) & X"000" & X"1") & eclat_false & eclat_false & eclat_false & \$12246_argument1\ & X"000" & X"0" & \$12190\(16 to 47) & \$12190\(120 to 121) & \$12190\(64 to 95) & \$12190\(96 to 103) & \$12190\(104 to 119);
                        state_var6675 <= \$12240_make_block_n587\;
                      when pause_setII6399 =>
                        \$ram_ptr_take\(0) := '0';
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"2") & "000"& X"000000" & X"1" & eclat_true & eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_setII6416 =>
                        \$ram_ptr_take\(0) := '0';
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"2") & \$12190\(16 to 47) & eclat_add(eclat_add(eclat_add(eclat_add(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1") & X"000" & X"1") & \$12190\(64 to 95) & \$12190\(96 to 103) & eclat_add(eclat_add(eclat_add(eclat_add(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1") & X"000" & X"1") & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_setII6420 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6418\ := \$ram_ptr_take\;
                        if \$v6418\(0) = '1' then
                          state_var6675 <= q_wait6417;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_add(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= eclat_resize(eclat_add(eclat_add(\$12190\(0 to 15) & X"000" & X"1") & eclat_resize(\$12246_argument1\,16)),31) & eclat_true;
                          state_var6675 <= pause_setI6415;
                        end if;
                      when pause_setII6424 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6422\ := \$ram_ptr_take\;
                        if \$v6422\(0) = '1' then
                          state_var6675 <= q_wait6421;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= eclat_resize(\$12190\(104 to 119),31) & eclat_true;
                          state_var6675 <= pause_setI6419;
                        end if;
                      when pause_setII6428 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6426\ := \$ram_ptr_take\;
                        if \$v6426\(0) = '1' then
                          state_var6675 <= q_wait6425;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(\$12190\(48 to 63) & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(64 to 95);
                          state_var6675 <= pause_setI6423;
                        end if;
                      when pause_setII6437 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6435\ := \$12246_argument1\;
                        case \$v6435\ is
                        when "000"& X"000000" & X"0" =>
                          eclat_print_string(of_string("======> "));
                          
                          eclat_print_int(\$12190\(16 to 46));
                          
                          eclat_print_newline(eclat_unit);
                          
                          \$13023\ := "000"& X"000000" & X"1" & eclat_true & \$12190\(0 to 15) & \$12190\(16 to 47) & eclat_add(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 95) & \$12190\(96 to 103) & \$12190\(104 to 119) & \$12190\(120 to 121);
                          \$v6434\ := \$ram_ptr_take\;
                          if \$v6434\(0) = '1' then
                            state_var6675 <= q_wait6433;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$13023\(80 to 95) & X"000" & X"1")));
                            state_var6675 <= pause_getI6431;
                          end if;
                        when others =>
                          eclat_print_string(of_string("unknown primitive"));
                          
                          \$13023\ := "000"& X"000000" & X"1" & eclat_true & \$12190\(0 to 15) & \$12190\(16 to 47) & eclat_add(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 95) & \$12190\(96 to 103) & \$12190\(104 to 119) & \$12190\(120 to 121);
                          \$v6434\ := \$ram_ptr_take\;
                          if \$v6434\(0) = '1' then
                            state_var6675 <= q_wait6433;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$13023\(80 to 95) & X"000" & X"1")));
                            state_var6675 <= pause_getI6431;
                          end if;
                        end case;
                      when pause_setII6446 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6444\ := \$12246_argument1\;
                        case \$v6444\ is
                        when "000"& X"000000" & X"0" =>
                          eclat_print_string(of_string("======> "));
                          
                          eclat_print_int(\$12190\(16 to 46));
                          
                          eclat_print_newline(eclat_unit);
                          
                          \$13052\ := "000"& X"000000" & X"1" & eclat_true & \$12190\(0 to 15) & \$12190\(16 to 47) & eclat_add(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1") & \$12190\(64 to 95) & \$12190\(96 to 103) & \$12190\(104 to 119) & \$12190\(120 to 121);
                          \$v6443\ := \$ram_ptr_take\;
                          if \$v6443\(0) = '1' then
                            state_var6675 <= q_wait6442;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$13052\(80 to 95) & X"000" & X"1")));
                            state_var6675 <= pause_getI6440;
                          end if;
                        when others =>
                          eclat_print_string(of_string("unknown primitive"));
                          
                          \$13052\ := "000"& X"000000" & X"1" & eclat_true & \$12190\(0 to 15) & \$12190\(16 to 47) & eclat_add(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1") & \$12190\(64 to 95) & \$12190\(96 to 103) & \$12190\(104 to 119) & \$12190\(120 to 121);
                          \$v6443\ := \$ram_ptr_take\;
                          if \$v6443\(0) = '1' then
                            state_var6675 <= q_wait6442;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$13052\(80 to 95) & X"000" & X"1")));
                            state_var6675 <= pause_getI6440;
                          end if;
                        end case;
                      when pause_setII6459 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6457\ := \$12246_argument1\;
                        case \$v6457\ is
                        when "000"& X"000000" & X"0" =>
                          eclat_print_string(of_string("======> "));
                          
                          eclat_print_int(\$12190\(16 to 46));
                          
                          eclat_print_newline(eclat_unit);
                          
                          \$13088\ := "000"& X"000000" & X"1" & eclat_true & \$12190\(0 to 15) & \$12190\(16 to 47) & eclat_add(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1") & \$12190\(64 to 95) & \$12190\(96 to 103) & \$12190\(104 to 119) & \$12190\(120 to 121);
                          \$v6456\ := \$ram_ptr_take\;
                          if \$v6456\(0) = '1' then
                            state_var6675 <= q_wait6455;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$13088\(80 to 95) & X"000" & X"1")));
                            state_var6675 <= pause_getI6453;
                          end if;
                        when others =>
                          eclat_print_string(of_string("unknown primitive"));
                          
                          \$13088\ := "000"& X"000000" & X"1" & eclat_true & \$12190\(0 to 15) & \$12190\(16 to 47) & eclat_add(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1") & \$12190\(64 to 95) & \$12190\(96 to 103) & \$12190\(104 to 119) & \$12190\(120 to 121);
                          \$v6456\ := \$ram_ptr_take\;
                          if \$v6456\(0) = '1' then
                            state_var6675 <= q_wait6455;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$13088\(80 to 95) & X"000" & X"1")));
                            state_var6675 <= pause_getI6453;
                          end if;
                        end case;
                      when pause_setII6476 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6474\ := \$12246_argument1\;
                        case \$v6474\ is
                        when "000"& X"000000" & X"0" =>
                          eclat_print_string(of_string("======> "));
                          
                          eclat_print_int(\$12190\(16 to 46));
                          
                          eclat_print_newline(eclat_unit);
                          
                          \$13134\ := "000"& X"000000" & X"1" & eclat_true & \$12190\(0 to 15) & \$12190\(16 to 47) & eclat_add(eclat_sub(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1") & X"000" & X"1") & \$12190\(64 to 95) & \$12190\(96 to 103) & \$12190\(104 to 119) & \$12190\(120 to 121);
                          \$v6473\ := \$ram_ptr_take\;
                          if \$v6473\(0) = '1' then
                            state_var6675 <= q_wait6472;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$13134\(80 to 95) & X"000" & X"1")));
                            state_var6675 <= pause_getI6470;
                          end if;
                        when others =>
                          eclat_print_string(of_string("unknown primitive"));
                          
                          \$13134\ := "000"& X"000000" & X"1" & eclat_true & \$12190\(0 to 15) & \$12190\(16 to 47) & eclat_add(eclat_sub(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1") & X"000" & X"1") & \$12190\(64 to 95) & \$12190\(96 to 103) & \$12190\(104 to 119) & \$12190\(120 to 121);
                          \$v6473\ := \$ram_ptr_take\;
                          if \$v6473\(0) = '1' then
                            state_var6675 <= q_wait6472;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$13134\(80 to 95) & X"000" & X"1")));
                            state_var6675 <= pause_getI6470;
                          end if;
                        end case;
                      when pause_setII6497 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6495\ := \$12246_argument1\;
                        case \$v6495\ is
                        when "000"& X"000000" & X"0" =>
                          eclat_print_string(of_string("======> "));
                          
                          eclat_print_int(\$12190\(16 to 46));
                          
                          eclat_print_newline(eclat_unit);
                          
                          \$13192\ := "000"& X"000000" & X"1" & eclat_true & \$12190\(0 to 15) & \$12190\(16 to 47) & eclat_add(eclat_sub(eclat_sub(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1") & X"000" & X"1") & X"000" & X"1") & \$12190\(64 to 95) & \$12190\(96 to 103) & \$12190\(104 to 119) & \$12190\(120 to 121);
                          \$v6494\ := \$ram_ptr_take\;
                          if \$v6494\(0) = '1' then
                            state_var6675 <= q_wait6493;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$13192\(80 to 95) & X"000" & X"1")));
                            state_var6675 <= pause_getI6491;
                          end if;
                        when others =>
                          eclat_print_string(of_string("unknown primitive"));
                          
                          \$13192\ := "000"& X"000000" & X"1" & eclat_true & \$12190\(0 to 15) & \$12190\(16 to 47) & eclat_add(eclat_sub(eclat_sub(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1") & X"000" & X"1") & X"000" & X"1") & \$12190\(64 to 95) & \$12190\(96 to 103) & \$12190\(104 to 119) & \$12190\(120 to 121);
                          \$v6494\ := \$ram_ptr_take\;
                          if \$v6494\(0) = '1' then
                            state_var6675 <= q_wait6493;
                          else
                            \$ram_ptr_take\(0) := '1';
                            \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$13192\(80 to 95) & X"000" & X"1")));
                            state_var6675 <= pause_getI6491;
                          end if;
                        end case;
                      when pause_setII6517 =>
                        \$ram_ptr_take\(0) := '0';
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"2") & \$12246_argument1\ & eclat_true & eclat_add(\$12190\(48 to 63) & X"000" & X"1") & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_setII6521 =>
                        \$ram_ptr_take\(0) := '0';
                        result5714 := eclat_add(\$12190\(0 to 15) & X"000" & X"2") & "000"& X"000000" & X"1" & eclat_true & \$12190\(48 to 63) & \$12190\(64 to 119) & \$12190\(120 to 121);
                        rdy5715 := eclat_true;
                        state_var6675 <= compute5716;
                      when pause_setII6529 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12421_w594_arg\ := eclat_add(\$12421_w594_arg\(0 to 15) & X"000" & X"1") & \$12421_w594_arg\(16 to 31) & \$12421_w594_arg\(32 to 47) & \$12421_w594_arg\(48 to 63);
                        state_var6675 <= \$12421_w594\;
                      when pause_setII6542 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12474_fill595_arg\ := eclat_add(\$12474_fill595_arg\(0 to 15) & X"000" & X"1") & eclat_sub(\$12474_fill595_arg\(16 to 31) & X"000" & X"1") & \$12474_fill595_arg\(32 to 47) & \$12474_fill595_arg\(48 to 79);
                        state_var6675 <= \$12474_fill595\;
                      when pause_setII6551 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12474_fill595_arg\ := X"000" & X"1" & \$12465_sp\ & eclat_resize(\$12246_argument1\,16) & \$12466\(64 to 95);
                        state_var6675 <= \$12474_fill595\;
                      when pause_setII6555 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12465_sp\ := eclat_add(\$12190\(48 to 63) & X"000" & X"1");
                        \$12199_make_block525_id\ := "000001000111";
                        \$12199_make_block525_arg\ := \$12465_sp\ & \$12190\(16 to 47) & \$12190\(64 to 95) & "11110111" & eclat_add(eclat_resize(\$12246_argument1\,16) & X"000" & X"1");
                        state_var6675 <= \$12199_make_block525\;
                      when pause_setII6576 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6574\ := \$ram_ptr_take\;
                        if \$v6574\(0) = '1' then
                          state_var6675 <= q_wait6573;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(X"3e80" & eclat_resize(\$12246_argument1\,16))));
                          state_var6675 <= pause_getI6571;
                        end if;
                      when pause_setII6580 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12564_fill596_arg\ := eclat_add(\$12564_fill596_arg\(0 to 15) & X"000" & X"1") & eclat_sub(\$12564_fill596_arg\(16 to 31) & X"000" & X"1") & \$12564_fill596_arg\(32 to 47) & \$12564_fill596_arg\(48 to 79);
                        state_var6675 <= \$12564_fill596\;
                      when pause_setII6589 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12564_fill596_arg\ := X"000" & X"1" & \$12190\(48 to 63) & eclat_resize(\$12246_argument1\,16) & \$12556\(64 to 95);
                        state_var6675 <= \$12564_fill596\;
                      when pause_setII6593 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12265_w0591_arg\ := eclat_add(\$12265_w0591_arg\(0 to 15) & X"000" & X"1") & eclat_sub(\$12265_w0591_arg\(16 to 31) & X"000" & X"1") & \$12265_w0591_arg\(32 to 47) & \$12265_w0591_arg\(48 to 63) & \$12265_w0591_arg\(64 to 95);
                        state_var6675 <= \$12265_w0591\;
                      when pause_setII6602 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12267_w1592_arg\ := eclat_add(\$12267_w1592_arg\(0 to 15) & X"000" & X"1") & \$12267_w1592_arg\(16 to 31) & \$12267_w1592_arg\(32 to 47) & \$12267_w1592_arg\(48 to 79);
                        state_var6675 <= \$12267_w1592\;
                      when pause_setII6610 =>
                        \$ram_ptr_take\(0) := '0';
                        \$v6608\ := \$code_ptr_take\;
                        if \$v6608\(0) = '1' then
                          state_var6675 <= q_wait6607;
                        else
                          \$code_ptr_take\(0) := '1';
                          \$code_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(\$12267_w1592_arg\(16 to 31) & X"000" & X"3") & \$12267_w1592_arg\(0 to 15))));
                          state_var6675 <= pause_getI6605;
                        end if;
                      when pause_setII6615 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12270_w3593_arg\ := eclat_add(\$12270_w3593_arg\(0 to 15) & X"000" & X"1") & eclat_add(\$12270_w3593_arg\(16 to 31) & X"000" & X"1") & \$12270_w3593_arg\(32 to 47) & \$12270_w3593_arg\(48 to 79);
                        state_var6675 <= \$12270_w3593\;
                      when pause_setII6620 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12270_w3593_arg\ := X"000" & X"1" & eclat_add(\$12266_sp\ & X"000" & X"1") & eclat_resize(\$12246_argument1\,16) & \$12257\(64 to 95);
                        state_var6675 <= \$12270_w3593\;
                      when pause_setII6624 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12265_w0591_arg\ := X"000" & X"0" & \$12256_sp\ & eclat_resize(\$12246_argument1\,16) & eclat_resize(\$12248_argument2\,16) & \$12257\(64 to 95);
                        state_var6675 <= \$12265_w0591\;
                      when pause_setII6628 =>
                        \$ram_ptr_take\(0) := '0';
                        \$12256_sp\ := eclat_add(\$12190\(48 to 63) & X"000" & X"1");
                        \$12199_make_block525_id\ := "000001010011";
                        \$12199_make_block525_arg\ := \$12256_sp\ & \$12190\(16 to 47) & \$12190\(64 to 95) & "11110111" & eclat_add(eclat_sub(eclat_mult(X"000" & X"2" & eclat_resize(\$12246_argument1\,16)) & X"000" & X"1") & eclat_resize(\$12248_argument2\,16));
                        state_var6675 <= \$12199_make_block525\;
                      when q_wait5719 =>
                        \$v5720\ := \$ram_ptr_take\;
                        if \$v5720\(0) = '1' then
                          state_var6675 <= q_wait5719;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$14250\(64 to 79)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= eclat_lor(eclat_lsl(eclat_resize(\$12199_make_block525_arg\(80 to 87),31) & "000"& X"00000" & X"18") & eclat_lsl(eclat_resize(
                          eclat_if(eclat_eq(\$12199_make_block525_arg\(88 to 103) & X"000" & X"0") & X"000" & X"1" & \$12199_make_block525_arg\(88 to 103)),31) & "000"& X"000000" & X"2")) & eclat_true;
                          state_var6675 <= pause_setI5717;
                        end if;
                      when q_wait5886 =>
                        \$v5887\ := \$ram_ptr_take\;
                        if \$v5887\(0) = '1' then
                          state_var6675 <= q_wait5886;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12235_apply579_arg\(60 to 90),16) & X"000" & X"0") & X"000" & X"1")));
                          state_var6675 <= pause_getI5884;
                        end if;
                      when q_wait5890 =>
                        \$v5891\ := \$ram_ptr_take\;
                        if \$v5891\(0) = '1' then
                          state_var6675 <= q_wait5890;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$14191_sp\));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$14180\(0 to 31);
                          state_var6675 <= pause_setI5888;
                        end if;
                      when q_wait5895 =>
                        \$v5896\ := \$ram_ptr_take\;
                        if \$v5896\(0) = '1' then
                          state_var6675 <= q_wait5895;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$14190_sp\));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$14183\(0 to 31);
                          state_var6675 <= pause_setI5893;
                        end if;
                      when q_wait5900 =>
                        \$v5901\ := \$ram_ptr_take\;
                        if \$v5901\(0) = '1' then
                          state_var6675 <= q_wait5900;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$14189_sp\));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$14186\(0 to 31);
                          state_var6675 <= pause_setI5898;
                        end if;
                      when q_wait5905 =>
                        \$v5906\ := \$ram_ptr_take\;
                        if \$v5906\(0) = '1' then
                          state_var6675 <= q_wait5905;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(\$14186\(32 to 47) & X"000" & X"1") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= eclat_resize(eclat_add(\$12235_apply579_arg\(44 to 59) & X"000" & X"1"),31) & eclat_true;
                          state_var6675 <= pause_setI5903;
                        end if;
                      when q_wait5909 =>
                        \$v5910\ := \$ram_ptr_take\;
                        if \$v5910\(0) = '1' then
                          state_var6675 <= q_wait5909;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(\$14186\(32 to 47) & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12235_apply579_arg\(110 to 141);
                          state_var6675 <= pause_setI5907;
                        end if;
                      when q_wait5913 =>
                        \$v5914\ := \$ram_ptr_take\;
                        if \$v5914\(0) = '1' then
                          state_var6675 <= q_wait5913;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$14186\(32 to 47)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= eclat_resize(\$12235_apply579_arg\(142 to 149),31) & eclat_true;
                          state_var6675 <= pause_setI5911;
                        end if;
                      when q_wait5918 =>
                        \$v5919\ := \$ram_ptr_take\;
                        if \$v5919\(0) = '1' then
                          state_var6675 <= q_wait5918;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$14183\(32 to 47) & X"000" & X"1")));
                          state_var6675 <= pause_getI5916;
                        end if;
                      when q_wait5923 =>
                        \$v5924\ := \$ram_ptr_take\;
                        if \$v5924\(0) = '1' then
                          state_var6675 <= q_wait5923;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$14180\(32 to 47) & X"000" & X"1")));
                          state_var6675 <= pause_getI5921;
                        end if;
                      when q_wait5928 =>
                        \$v5929\ := \$ram_ptr_take\;
                        if \$v5929\(0) = '1' then
                          state_var6675 <= q_wait5928;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12235_apply579_arg\(92 to 107) & X"000" & X"1")));
                          state_var6675 <= pause_getI5926;
                        end if;
                      when q_wait5939 =>
                        \$v5940\ := \$ram_ptr_take\;
                        if \$v5940\(0) = '1' then
                          state_var6675 <= q_wait5939;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12237_binop_int584_arg\(80 to 95) & X"000" & X"1")));
                          state_var6675 <= pause_getI5937;
                        end if;
                      when q_wait5944 =>
                        \$v5945\ := \$ram_ptr_take\;
                        if \$v5945\(0) = '1' then
                          state_var6675 <= q_wait5944;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12239_binop_compare586_arg\(80 to 95) & X"000" & X"1")));
                          state_var6675 <= pause_getI5942;
                        end if;
                      when q_wait5948 =>
                        \$v5949\ := \$ram_ptr_take\;
                        if \$v5949\(0) = '1' then
                          state_var6675 <= q_wait5948;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$13996\(64 to 94),16) & X"000" & X"2") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$14003_v\;
                          state_var6675 <= pause_setI5946;
                        end if;
                      when q_wait5952 =>
                        \$v5953\ := \$ram_ptr_take\;
                        if \$v5953\(0) = '1' then
                          state_var6675 <= q_wait5952;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$14001_sp\ & X"000" & X"1")));
                          state_var6675 <= pause_getI5950;
                        end if;
                      when q_wait5957 =>
                        \$v5958\ := \$ram_ptr_take\;
                        if \$v5958\(0) = '1' then
                          state_var6675 <= q_wait5957;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$13996\(64 to 94),16) & X"000" & X"1") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$14014_v\;
                          state_var6675 <= pause_setI5955;
                        end if;
                      when q_wait5961 =>
                        \$v5962\ := \$ram_ptr_take\;
                        if \$v5962\(0) = '1' then
                          state_var6675 <= q_wait5961;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12240_make_block_n587_arg\(16 to 31) & X"000" & X"1")));
                          state_var6675 <= pause_getI5959;
                        end if;
                      when q_wait5966 =>
                        \$v5967\ := \$ram_ptr_take\;
                        if \$v5967\(0) = '1' then
                          state_var6675 <= q_wait5966;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$13996\(64 to 94),16) & X"000" & X"0") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$13996\(0 to 31);
                          state_var6675 <= pause_setI5964;
                        end if;
                      when q_wait5971 =>
                        \$v5972\ := \$code_ptr_take\;
                        if \$v5972\(0) = '1' then
                          state_var6675 <= q_wait5971;
                        else
                          \$code_ptr_take\(0) := '1';
                          \$code_ptr\ <= to_integer(unsigned(eclat_add(\$12241_branch_if589_arg\(1 to 16) & X"000" & X"1")));
                          state_var6675 <= pause_getI5969;
                        end if;
                      when q_wait5976 =>
                        \$v5977\ := \$ram_ptr_take\;
                        if \$v5977\(0) = '1' then
                          state_var6675 <= q_wait5976;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"0") & X"000" & X"1")));
                          state_var6675 <= pause_getI5974;
                        end if;
                      when q_wait5980 =>
                        \$v5981\ := \$ram_ptr_take\;
                        if \$v5981\(0) = '1' then
                          state_var6675 <= q_wait5980;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI5978;
                        end if;
                      when q_wait5984 =>
                        \$v5985\ := \$ram_ptr_take\;
                        if \$v5985\(0) = '1' then
                          state_var6675 <= q_wait5984;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"2") & X"000" & X"1")));
                          state_var6675 <= pause_getI5982;
                        end if;
                      when q_wait5988 =>
                        \$v5989\ := \$ram_ptr_take\;
                        if \$v5989\(0) = '1' then
                          state_var6675 <= q_wait5988;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"3") & X"000" & X"1")));
                          state_var6675 <= pause_getI5986;
                        end if;
                      when q_wait5992 =>
                        \$v5993\ := \$ram_ptr_take\;
                        if \$v5993\(0) = '1' then
                          state_var6675 <= q_wait5992;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"4") & X"000" & X"1")));
                          state_var6675 <= pause_getI5990;
                        end if;
                      when q_wait5996 =>
                        \$v5997\ := \$ram_ptr_take\;
                        if \$v5997\(0) = '1' then
                          state_var6675 <= q_wait5996;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"5") & X"000" & X"1")));
                          state_var6675 <= pause_getI5994;
                        end if;
                      when q_wait6000 =>
                        \$v6001\ := \$ram_ptr_take\;
                        if \$v6001\(0) = '1' then
                          state_var6675 <= q_wait6000;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"6") & X"000" & X"1")));
                          state_var6675 <= pause_getI5998;
                        end if;
                      when q_wait6004 =>
                        \$v6005\ := \$ram_ptr_take\;
                        if \$v6005\(0) = '1' then
                          state_var6675 <= q_wait6004;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"7") & X"000" & X"1")));
                          state_var6675 <= pause_getI6002;
                        end if;
                      when q_wait6008 =>
                        \$v6009\ := \$ram_ptr_take\;
                        if \$v6009\(0) = '1' then
                          state_var6675 <= q_wait6008;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6006;
                        end if;
                      when q_wait6012 =>
                        \$v6013\ := \$ram_ptr_take\;
                        if \$v6013\(0) = '1' then
                          state_var6675 <= q_wait6012;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6010;
                        end if;
                      when q_wait6016 =>
                        \$v6017\ := \$ram_ptr_take\;
                        if \$v6017\(0) = '1' then
                          state_var6675 <= q_wait6016;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_add(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6014;
                        end if;
                      when q_wait6020 =>
                        \$v6021\ := \$ram_ptr_take\;
                        if \$v6021\(0) = '1' then
                          state_var6675 <= q_wait6020;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6018;
                        end if;
                      when q_wait6024 =>
                        \$v6025\ := \$ram_ptr_take\;
                        if \$v6025\(0) = '1' then
                          state_var6675 <= q_wait6024;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_add(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"2") & X"000" & X"1")));
                          state_var6675 <= pause_getI6022;
                        end if;
                      when q_wait6028 =>
                        \$v6029\ := \$ram_ptr_take\;
                        if \$v6029\(0) = '1' then
                          state_var6675 <= q_wait6028;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6026;
                        end if;
                      when q_wait6032 =>
                        \$v6033\ := \$ram_ptr_take\;
                        if \$v6033\(0) = '1' then
                          state_var6675 <= q_wait6032;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_add(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"3") & X"000" & X"1")));
                          state_var6675 <= pause_getI6030;
                        end if;
                      when q_wait6036 =>
                        \$v6037\ := \$ram_ptr_take\;
                        if \$v6037\(0) = '1' then
                          state_var6675 <= q_wait6036;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6034;
                        end if;
                      when q_wait6040 =>
                        \$v6041\ := \$ram_ptr_take\;
                        if \$v6041\(0) = '1' then
                          state_var6675 <= q_wait6040;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_add(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"4") & X"000" & X"1")));
                          state_var6675 <= pause_getI6038;
                        end if;
                      when q_wait6044 =>
                        \$v6045\ := \$ram_ptr_take\;
                        if \$v6045\(0) = '1' then
                          state_var6675 <= q_wait6044;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6042;
                        end if;
                      when q_wait6048 =>
                        \$v6049\ := \$ram_ptr_take\;
                        if \$v6049\(0) = '1' then
                          state_var6675 <= q_wait6048;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_add(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"5") & X"000" & X"1")));
                          state_var6675 <= pause_getI6046;
                        end if;
                      when q_wait6052 =>
                        \$v6053\ := \$ram_ptr_take\;
                        if \$v6053\(0) = '1' then
                          state_var6675 <= q_wait6052;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6050;
                        end if;
                      when q_wait6056 =>
                        \$v6057\ := \$ram_ptr_take\;
                        if \$v6057\(0) = '1' then
                          state_var6675 <= q_wait6056;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_add(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"6") & X"000" & X"1")));
                          state_var6675 <= pause_getI6054;
                        end if;
                      when q_wait6060 =>
                        \$v6061\ := \$ram_ptr_take\;
                        if \$v6061\(0) = '1' then
                          state_var6675 <= q_wait6060;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6058;
                        end if;
                      when q_wait6064 =>
                        \$v6065\ := \$ram_ptr_take\;
                        if \$v6065\(0) = '1' then
                          state_var6675 <= q_wait6064;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_add(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"7") & X"000" & X"1")));
                          state_var6675 <= pause_getI6062;
                        end if;
                      when q_wait6068 =>
                        \$v6069\ := \$ram_ptr_take\;
                        if \$v6069\(0) = '1' then
                          state_var6675 <= q_wait6068;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6066;
                        end if;
                      when q_wait6072 =>
                        \$v6073\ := \$ram_ptr_take\;
                        if \$v6073\(0) = '1' then
                          state_var6675 <= q_wait6072;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(64 to 94),16) & eclat_sub(X"000" & X"1" & X"000" & X"1")) & X"000" & X"1")));
                          state_var6675 <= pause_getI6070;
                        end if;
                      when q_wait6076 =>
                        \$v6077\ := \$ram_ptr_take\;
                        if \$v6077\(0) = '1' then
                          state_var6675 <= q_wait6076;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(64 to 94),16) & eclat_sub(X"000" & X"2" & X"000" & X"1")) & X"000" & X"1")));
                          state_var6675 <= pause_getI6074;
                        end if;
                      when q_wait6080 =>
                        \$v6081\ := \$ram_ptr_take\;
                        if \$v6081\(0) = '1' then
                          state_var6675 <= q_wait6080;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(64 to 94),16) & eclat_sub(X"000" & X"3" & X"000" & X"1")) & X"000" & X"1")));
                          state_var6675 <= pause_getI6078;
                        end if;
                      when q_wait6084 =>
                        \$v6085\ := \$ram_ptr_take\;
                        if \$v6085\(0) = '1' then
                          state_var6675 <= q_wait6084;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(64 to 94),16) & eclat_sub(X"000" & X"4" & X"000" & X"1")) & X"000" & X"1")));
                          state_var6675 <= pause_getI6082;
                        end if;
                      when q_wait6088 =>
                        \$v6089\ := \$ram_ptr_take\;
                        if \$v6089\(0) = '1' then
                          state_var6675 <= q_wait6088;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(64 to 94),16) & eclat_sub(X"000" & X"1" & X"000" & X"1")) & X"000" & X"1")));
                          state_var6675 <= pause_getI6086;
                        end if;
                      when q_wait6092 =>
                        \$v6093\ := \$ram_ptr_take\;
                        if \$v6093\(0) = '1' then
                          state_var6675 <= q_wait6092;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6090;
                        end if;
                      when q_wait6096 =>
                        \$v6097\ := \$ram_ptr_take\;
                        if \$v6097\(0) = '1' then
                          state_var6675 <= q_wait6096;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(64 to 94),16) & eclat_sub(X"000" & X"2" & X"000" & X"1")) & X"000" & X"1")));
                          state_var6675 <= pause_getI6094;
                        end if;
                      when q_wait6100 =>
                        \$v6101\ := \$ram_ptr_take\;
                        if \$v6101\(0) = '1' then
                          state_var6675 <= q_wait6100;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6098;
                        end if;
                      when q_wait6104 =>
                        \$v6105\ := \$ram_ptr_take\;
                        if \$v6105\(0) = '1' then
                          state_var6675 <= q_wait6104;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(64 to 94),16) & eclat_sub(X"000" & X"3" & X"000" & X"1")) & X"000" & X"1")));
                          state_var6675 <= pause_getI6102;
                        end if;
                      when q_wait6108 =>
                        \$v6109\ := \$ram_ptr_take\;
                        if \$v6109\(0) = '1' then
                          state_var6675 <= q_wait6108;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6106;
                        end if;
                      when q_wait6112 =>
                        \$v6113\ := \$ram_ptr_take\;
                        if \$v6113\(0) = '1' then
                          state_var6675 <= q_wait6112;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(64 to 94),16) & eclat_sub(X"000" & X"4" & X"000" & X"1")) & X"000" & X"1")));
                          state_var6675 <= pause_getI6110;
                        end if;
                      when q_wait6116 =>
                        \$v6117\ := \$ram_ptr_take\;
                        if \$v6117\(0) = '1' then
                          state_var6675 <= q_wait6116;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6114;
                        end if;
                      when q_wait6120 =>
                        \$v6121\ := \$ram_ptr_take\;
                        if \$v6121\(0) = '1' then
                          state_var6675 <= q_wait6120;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$13539_loop_push598_arg\(0 to 15)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$13589\;
                          state_var6675 <= pause_setI6118;
                        end if;
                      when q_wait6124 =>
                        \$v6125\ := \$ram_ptr_take\;
                        if \$v6125\(0) = '1' then
                          state_var6675 <= q_wait6124;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$13539_loop_push598_arg\(24 to 54),16) & eclat_resize(eclat_add(\$13539_loop_push598_arg\(16 to 23) & "00000010"),16)) & X"000" & X"1")));
                          state_var6675 <= pause_getI6122;
                        end if;
                      when q_wait6129 =>
                        \$v6130\ := \$ram_ptr_take\;
                        if \$v6130\(0) = '1' then
                          state_var6675 <= q_wait6129;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(64 to 94),16) & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6127;
                        end if;
                      when q_wait6133 =>
                        \$v6134\ := \$ram_ptr_take\;
                        if \$v6134\(0) = '1' then
                          state_var6675 <= q_wait6133;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$12190\(64 to 94),16)));
                          state_var6675 <= pause_getI6131;
                        end if;
                      when q_wait6137 =>
                        \$v6138\ := \$ram_ptr_take\;
                        if \$v6138\(0) = '1' then
                          state_var6675 <= q_wait6137;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6135;
                        end if;
                      when q_wait6141 =>
                        \$v6142\ := \$ram_ptr_take\;
                        if \$v6142\(0) = '1' then
                          state_var6675 <= q_wait6141;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6139;
                        end if;
                      when q_wait6145 =>
                        \$v6146\ := \$ram_ptr_take\;
                        if \$v6146\(0) = '1' then
                          state_var6675 <= q_wait6145;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6143;
                        end if;
                      when q_wait6149 =>
                        \$v6150\ := \$ram_ptr_take\;
                        if \$v6150\(0) = '1' then
                          state_var6675 <= q_wait6149;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6147;
                        end if;
                      when q_wait6153 =>
                        \$v6154\ := \$ram_ptr_take\;
                        if \$v6154\(0) = '1' then
                          state_var6675 <= q_wait6153;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & X"000" & X"0") & X"000" & X"1")));
                          state_var6675 <= pause_getI6151;
                        end if;
                      when q_wait6157 =>
                        \$v6158\ := \$ram_ptr_take\;
                        if \$v6158\(0) = '1' then
                          state_var6675 <= q_wait6157;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6155;
                        end if;
                      when q_wait6161 =>
                        \$v6162\ := \$ram_ptr_take\;
                        if \$v6162\(0) = '1' then
                          state_var6675 <= q_wait6161;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & X"000" & X"2") & X"000" & X"1")));
                          state_var6675 <= pause_getI6159;
                        end if;
                      when q_wait6165 =>
                        \$v6166\ := \$ram_ptr_take\;
                        if \$v6166\(0) = '1' then
                          state_var6675 <= q_wait6165;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & X"000" & X"3") & X"000" & X"1")));
                          state_var6675 <= pause_getI6163;
                        end if;
                      when q_wait6169 =>
                        \$v6170\ := \$ram_ptr_take\;
                        if \$v6170\(0) = '1' then
                          state_var6675 <= q_wait6169;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & X"000" & X"0") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$13699_v\;
                          state_var6675 <= pause_setI6167;
                        end if;
                      when q_wait6173 =>
                        \$v6174\ := \$ram_ptr_take\;
                        if \$v6174\(0) = '1' then
                          state_var6675 <= q_wait6173;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12190\(48 to 63) & X"000" & X"1")));
                          state_var6675 <= pause_getI6171;
                        end if;
                      when q_wait6177 =>
                        \$v6178\ := \$ram_ptr_take\;
                        if \$v6178\(0) = '1' then
                          state_var6675 <= q_wait6177;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & X"000" & X"1") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$13712_v\;
                          state_var6675 <= pause_setI6175;
                        end if;
                      when q_wait6181 =>
                        \$v6182\ := \$ram_ptr_take\;
                        if \$v6182\(0) = '1' then
                          state_var6675 <= q_wait6181;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12190\(48 to 63) & X"000" & X"1")));
                          state_var6675 <= pause_getI6179;
                        end if;
                      when q_wait6185 =>
                        \$v6186\ := \$ram_ptr_take\;
                        if \$v6186\(0) = '1' then
                          state_var6675 <= q_wait6185;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & X"000" & X"2") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$13725_v\;
                          state_var6675 <= pause_setI6183;
                        end if;
                      when q_wait6189 =>
                        \$v6190\ := \$ram_ptr_take\;
                        if \$v6190\(0) = '1' then
                          state_var6675 <= q_wait6189;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12190\(48 to 63) & X"000" & X"1")));
                          state_var6675 <= pause_getI6187;
                        end if;
                      when q_wait6193 =>
                        \$v6194\ := \$ram_ptr_take\;
                        if \$v6194\(0) = '1' then
                          state_var6675 <= q_wait6193;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & X"000" & X"3") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$13738_v\;
                          state_var6675 <= pause_setI6191;
                        end if;
                      when q_wait6197 =>
                        \$v6198\ := \$ram_ptr_take\;
                        if \$v6198\(0) = '1' then
                          state_var6675 <= q_wait6197;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12190\(48 to 63) & X"000" & X"1")));
                          state_var6675 <= pause_getI6195;
                        end if;
                      when q_wait6201 =>
                        \$v6202\ := \$ram_ptr_take\;
                        if \$v6202\(0) = '1' then
                          state_var6675 <= q_wait6201;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$12190\(16 to 46),16)));
                          state_var6675 <= pause_getI6199;
                        end if;
                      when q_wait6205 =>
                        \$v6206\ := \$ram_ptr_take\;
                        if \$v6206\(0) = '1' then
                          state_var6675 <= q_wait6205;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & eclat_resize(\$13767_v\(0 to 30),16)) & X"000" & X"1")));
                          state_var6675 <= pause_getI6203;
                        end if;
                      when q_wait6209 =>
                        \$v6210\ := \$ram_ptr_take\;
                        if \$v6210\(0) = '1' then
                          state_var6675 <= q_wait6209;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12190\(48 to 63) & X"000" & X"1")));
                          state_var6675 <= pause_getI6207;
                        end if;
                      when q_wait6213 =>
                        \$v6214\ := \$ram_ptr_take\;
                        if \$v6214\(0) = '1' then
                          state_var6675 <= q_wait6213;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & eclat_resize(\$13784_v\(0 to 30),16)) & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$13785_v\;
                          state_var6675 <= pause_setI6211;
                        end if;
                      when q_wait6217 =>
                        \$v6218\ := \$ram_ptr_take\;
                        if \$v6218\(0) = '1' then
                          state_var6675 <= q_wait6217;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6215;
                        end if;
                      when q_wait6221 =>
                        \$v6222\ := \$ram_ptr_take\;
                        if \$v6222\(0) = '1' then
                          state_var6675 <= q_wait6221;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12190\(48 to 63) & X"000" & X"1")));
                          state_var6675 <= pause_getI6219;
                        end if;
                      when q_wait6225 =>
                        \$v6226\ := \$ram_ptr_take\;
                        if \$v6226\(0) = '1' then
                          state_var6675 <= q_wait6225;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & eclat_resize(\$13807_v\(0 to 30),16)) & X"000" & X"1")));
                          state_var6675 <= pause_getI6223;
                        end if;
                      when q_wait6229 =>
                        \$v6230\ := \$ram_ptr_take\;
                        if \$v6230\(0) = '1' then
                          state_var6675 <= q_wait6229;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12190\(48 to 63) & X"000" & X"1")));
                          state_var6675 <= pause_getI6227;
                        end if;
                      when q_wait6233 =>
                        \$v6234\ := \$ram_ptr_take\;
                        if \$v6234\(0) = '1' then
                          state_var6675 <= q_wait6233;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & eclat_resize(\$13824_v\(0 to 30),16)) & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$13825_v\;
                          state_var6675 <= pause_setI6231;
                        end if;
                      when q_wait6237 =>
                        \$v6238\ := \$ram_ptr_take\;
                        if \$v6238\(0) = '1' then
                          state_var6675 <= q_wait6237;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6235;
                        end if;
                      when q_wait6241 =>
                        \$v6242\ := \$ram_ptr_take\;
                        if \$v6242\(0) = '1' then
                          state_var6675 <= q_wait6241;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12190\(48 to 63) & X"000" & X"1")));
                          state_var6675 <= pause_getI6239;
                        end if;
                      when q_wait6245 =>
                        \$v6246\ := \$ram_ptr_take\;
                        if \$v6246\(0) = '1' then
                          state_var6675 <= q_wait6245;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6243;
                        end if;
                      when q_wait6249 =>
                        \$v6250\ := \$ram_ptr_take\;
                        if \$v6250\(0) = '1' then
                          state_var6675 <= q_wait6249;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_sub(eclat_sub(\$12190\(104 to 119) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6247;
                        end if;
                      when q_wait6253 =>
                        \$v6254\ := \$ram_ptr_take\;
                        if \$v6254\(0) = '1' then
                          state_var6675 <= q_wait6253;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_sub(\$12190\(104 to 119) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6251;
                        end if;
                      when q_wait6257 =>
                        \$v6258\ := \$ram_ptr_take\;
                        if \$v6258\(0) = '1' then
                          state_var6675 <= q_wait6257;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(104 to 119) & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6255;
                        end if;
                      when q_wait6261 =>
                        \$v6262\ := \$ram_ptr_take\;
                        if \$v6262\(0) = '1' then
                          state_var6675 <= q_wait6261;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12190\(104 to 119) & X"000" & X"1")));
                          state_var6675 <= pause_getI6259;
                        end if;
                      when q_wait6265 =>
                        \$v6266\ := \$ram_ptr_take\;
                        if \$v6266\(0) = '1' then
                          state_var6675 <= q_wait6265;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6263;
                        end if;
                      when q_wait6269 =>
                        \$v6270\ := \$ram_ptr_take\;
                        if \$v6270\(0) = '1' then
                          state_var6675 <= q_wait6269;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6267;
                        end if;
                      when q_wait6273 =>
                        \$v6274\ := \$ram_ptr_take\;
                        if \$v6274\(0) = '1' then
                          state_var6675 <= q_wait6273;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6271;
                        end if;
                      when q_wait6277 =>
                        \$v6278\ := \$ram_ptr_take\;
                        if \$v6278\(0) = '1' then
                          state_var6675 <= q_wait6277;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6275;
                        end if;
                      when q_wait6281 =>
                        \$v6282\ := \$ram_ptr_take\;
                        if \$v6282\(0) = '1' then
                          state_var6675 <= q_wait6281;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & eclat_resize(\$12246_argument1\,16)) & X"000" & X"1")));
                          state_var6675 <= pause_getI6279;
                        end if;
                      when q_wait6285 =>
                        \$v6286\ := \$ram_ptr_take\;
                        if \$v6286\(0) = '1' then
                          state_var6675 <= q_wait6285;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_add(\$12190\(48 to 63) & X"000" & X"1") & eclat_resize(\$12246_argument1\,16)) & X"000" & X"1")));
                          state_var6675 <= pause_getI6283;
                        end if;
                      when q_wait6289 =>
                        \$v6290\ := \$ram_ptr_take\;
                        if \$v6290\(0) = '1' then
                          state_var6675 <= q_wait6289;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6287;
                        end if;
                      when q_wait6293 =>
                        \$v6294\ := \$ram_ptr_take\;
                        if \$v6294\(0) = '1' then
                          state_var6675 <= q_wait6293;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & eclat_resize(\$12246_argument1\,16))));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6291;
                        end if;
                      when q_wait6297 =>
                        \$v6298\ := \$ram_ptr_take\;
                        if \$v6298\(0) = '1' then
                          state_var6675 <= q_wait6297;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(64 to 94),16) & eclat_sub(eclat_resize(\$12246_argument1\,16) & X"000" & X"1")) & X"000" & X"1")));
                          state_var6675 <= pause_getI6295;
                        end if;
                      when q_wait6301 =>
                        \$v6302\ := \$ram_ptr_take\;
                        if \$v6302\(0) = '1' then
                          state_var6675 <= q_wait6301;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(64 to 94),16) & eclat_sub(eclat_resize(\$12246_argument1\,16) & X"000" & X"1")) & X"000" & X"1")));
                          state_var6675 <= pause_getI6299;
                        end if;
                      when q_wait6305 =>
                        \$v6306\ := \$ram_ptr_take\;
                        if \$v6306\(0) = '1' then
                          state_var6675 <= q_wait6305;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6303;
                        end if;
                      when q_wait6309 =>
                        \$v6310\ := \$ram_ptr_take\;
                        if \$v6310\(0) = '1' then
                          state_var6675 <= q_wait6309;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= eclat_resize(eclat_add(eclat_add(\$12190\(0 to 15) & X"000" & X"1") & eclat_resize(\$12246_argument1\,16)),31) & eclat_true;
                          state_var6675 <= pause_setI6307;
                        end if;
                      when q_wait6313 =>
                        \$v6314\ := \$ram_ptr_take\;
                        if \$v6314\(0) = '1' then
                          state_var6675 <= q_wait6313;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(\$12190\(48 to 63) & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(64 to 95);
                          state_var6675 <= pause_setI6311;
                        end if;
                      when q_wait6317 =>
                        \$v6318\ := \$ram_ptr_take\;
                        if \$v6318\(0) = '1' then
                          state_var6675 <= q_wait6317;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= eclat_resize(\$12190\(96 to 103),31) & eclat_true;
                          state_var6675 <= pause_setI6315;
                        end if;
                      when q_wait6321 =>
                        \$v6322\ := \$ram_ptr_take\;
                        if \$v6322\(0) = '1' then
                          state_var6675 <= q_wait6321;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & X"000" & X"0") & X"000" & X"1")));
                          state_var6675 <= pause_getI6319;
                        end if;
                      when q_wait6325 =>
                        \$v6326\ := \$ram_ptr_take\;
                        if \$v6326\(0) = '1' then
                          state_var6675 <= q_wait6325;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & X"000" & X"0") & X"000" & X"1")));
                          state_var6675 <= pause_getI6323;
                        end if;
                      when q_wait6329 =>
                        \$v6330\ := \$ram_ptr_take\;
                        if \$v6330\(0) = '1' then
                          state_var6675 <= q_wait6329;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_sub(eclat_sub(\$12190\(48 to 63) & eclat_resize(\$12246_argument1\,16)) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6327;
                        end if;
                      when q_wait6333 =>
                        \$v6334\ := \$ram_ptr_take\;
                        if \$v6334\(0) = '1' then
                          state_var6675 <= q_wait6333;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_sub(\$12190\(48 to 63) & eclat_resize(\$12246_argument1\,16)) & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6331;
                        end if;
                      when q_wait6337 =>
                        \$v6338\ := \$ram_ptr_take\;
                        if \$v6338\(0) = '1' then
                          state_var6675 <= q_wait6337;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & eclat_resize(\$12246_argument1\,16)) & X"000" & X"1")));
                          state_var6675 <= pause_getI6335;
                        end if;
                      when q_wait6342 =>
                        \$v6343\ := \$ram_ptr_take\;
                        if \$v6343\(0) = '1' then
                          state_var6675 <= q_wait6342;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12782_w597_arg\(32 to 62),16) & eclat_resize(eclat_add(\$12782_w597_arg\(0 to 7) & "00000010"),16)) & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12820_v\;
                          state_var6675 <= pause_setI6340;
                        end if;
                      when q_wait6346 =>
                        \$v6347\ := \$ram_ptr_take\;
                        if \$v6347\(0) = '1' then
                          state_var6675 <= q_wait6346;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12782_w597_arg\(8 to 23) & X"000" & X"1")));
                          state_var6675 <= pause_getI6344;
                        end if;
                      when q_wait6351 =>
                        \$v6352\ := \$ram_ptr_take\;
                        if \$v6352\(0) = '1' then
                          state_var6675 <= q_wait6351;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_sub(\$12783_sp\ & X"000" & X"1") & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6349;
                        end if;
                      when q_wait6355 =>
                        \$v6356\ := \$ram_ptr_take\;
                        if \$v6356\(0) = '1' then
                          state_var6675 <= q_wait6355;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12783_sp\ & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6353;
                        end if;
                      when q_wait6359 =>
                        \$v6360\ := \$ram_ptr_take\;
                        if \$v6360\(0) = '1' then
                          state_var6675 <= q_wait6359;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12783_sp\ & X"000" & X"1")));
                          state_var6675 <= pause_getI6357;
                        end if;
                      when q_wait6363 =>
                        \$v6364\ := \$ram_ptr_take\;
                        if \$v6364\(0) = '1' then
                          state_var6675 <= q_wait6363;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12770\(64 to 94),16) & X"000" & X"1") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12770\(32 to 63);
                          state_var6675 <= pause_setI6361;
                        end if;
                      when q_wait6367 =>
                        \$v6368\ := \$ram_ptr_take\;
                        if \$v6368\(0) = '1' then
                          state_var6675 <= q_wait6367;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12770\(64 to 94),16) & X"000" & X"0") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= eclat_resize(eclat_sub(eclat_add(\$12190\(0 to 15) & X"000" & X"2") & X"000" & X"3"),31) & eclat_true;
                          state_var6675 <= pause_setI6365;
                        end if;
                      when q_wait6372 =>
                        \$v6373\ := \$ram_ptr_take\;
                        if \$v6373\(0) = '1' then
                          state_var6675 <= q_wait6372;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6370;
                        end if;
                      when q_wait6376 =>
                        \$v6377\ := \$ram_ptr_take\;
                        if \$v6377\(0) = '1' then
                          state_var6675 <= q_wait6376;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(X"3e80" & eclat_resize(\$12246_argument1\,16))));
                          state_var6675 <= pause_getI6374;
                        end if;
                      when q_wait6380 =>
                        \$v6381\ := \$ram_ptr_take\;
                        if \$v6381\(0) = '1' then
                          state_var6675 <= q_wait6380;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(X"3e80" & eclat_resize(\$12246_argument1\,16))));
                          state_var6675 <= pause_getI6378;
                        end if;
                      when q_wait6384 =>
                        \$v6385\ := \$ram_ptr_take\;
                        if \$v6385\(0) = '1' then
                          state_var6675 <= q_wait6384;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6382;
                        end if;
                      when q_wait6388 =>
                        \$v6389\ := \$ram_ptr_take\;
                        if \$v6389\(0) = '1' then
                          state_var6675 <= q_wait6388;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(X"3e80" & eclat_resize(\$12246_argument1\,16))));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6386;
                        end if;
                      when q_wait6392 =>
                        \$v6393\ := \$ram_ptr_take\;
                        if \$v6393\(0) = '1' then
                          state_var6675 <= q_wait6392;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6390;
                        end if;
                      when q_wait6396 =>
                        \$v6397\ := \$ram_ptr_take\;
                        if \$v6397\(0) = '1' then
                          state_var6675 <= q_wait6396;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & eclat_resize(\$12246_argument1\,16)) & X"000" & X"1")));
                          state_var6675 <= pause_getI6394;
                        end if;
                      when q_wait6400 =>
                        \$v6401\ := \$ram_ptr_take\;
                        if \$v6401\(0) = '1' then
                          state_var6675 <= q_wait6400;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & eclat_resize(\$12246_argument1\,16)) & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12929_v\;
                          state_var6675 <= pause_setI6398;
                        end if;
                      when q_wait6404 =>
                        \$v6405\ := \$ram_ptr_take\;
                        if \$v6405\(0) = '1' then
                          state_var6675 <= q_wait6404;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12190\(48 to 63) & X"000" & X"1")));
                          state_var6675 <= pause_getI6402;
                        end if;
                      when q_wait6408 =>
                        \$v6409\ := \$code_ptr_take\;
                        if \$v6409\(0) = '1' then
                          state_var6675 <= q_wait6408;
                        else
                          \$code_ptr_take\(0) := '1';
                          \$code_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(\$12190\(0 to 15) & X"000" & X"2") & \$12953_ofs\)));
                          state_var6675 <= pause_getI6406;
                        end if;
                      when q_wait6412 =>
                        \$v6413\ := \$ram_ptr_take\;
                        if \$v6413\(0) = '1' then
                          state_var6675 <= q_wait6412;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$12190\(16 to 46),16)));
                          state_var6675 <= pause_getI6410;
                        end if;
                      when q_wait6417 =>
                        \$v6418\ := \$ram_ptr_take\;
                        if \$v6418\(0) = '1' then
                          state_var6675 <= q_wait6417;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_add(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= eclat_resize(eclat_add(eclat_add(\$12190\(0 to 15) & X"000" & X"1") & eclat_resize(\$12246_argument1\,16)),31) & eclat_true;
                          state_var6675 <= pause_setI6415;
                        end if;
                      when q_wait6421 =>
                        \$v6422\ := \$ram_ptr_take\;
                        if \$v6422\(0) = '1' then
                          state_var6675 <= q_wait6421;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= eclat_resize(\$12190\(104 to 119),31) & eclat_true;
                          state_var6675 <= pause_setI6419;
                        end if;
                      when q_wait6425 =>
                        \$v6426\ := \$ram_ptr_take\;
                        if \$v6426\(0) = '1' then
                          state_var6675 <= q_wait6425;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(\$12190\(48 to 63) & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(64 to 95);
                          state_var6675 <= pause_setI6423;
                        end if;
                      when q_wait6429 =>
                        \$v6430\ := \$ram_ptr_take\;
                        if \$v6430\(0) = '1' then
                          state_var6675 <= q_wait6429;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= eclat_resize(\$12190\(96 to 103),31) & eclat_true;
                          state_var6675 <= pause_setI6427;
                        end if;
                      when q_wait6433 =>
                        \$v6434\ := \$ram_ptr_take\;
                        if \$v6434\(0) = '1' then
                          state_var6675 <= q_wait6433;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$13023\(80 to 95) & X"000" & X"1")));
                          state_var6675 <= pause_getI6431;
                        end if;
                      when q_wait6438 =>
                        \$v6439\ := \$ram_ptr_take\;
                        if \$v6439\(0) = '1' then
                          state_var6675 <= q_wait6438;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(64 to 95);
                          state_var6675 <= pause_setI6436;
                        end if;
                      when q_wait6442 =>
                        \$v6443\ := \$ram_ptr_take\;
                        if \$v6443\(0) = '1' then
                          state_var6675 <= q_wait6442;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$13052\(80 to 95) & X"000" & X"1")));
                          state_var6675 <= pause_getI6440;
                        end if;
                      when q_wait6447 =>
                        \$v6448\ := \$ram_ptr_take\;
                        if \$v6448\(0) = '1' then
                          state_var6675 <= q_wait6447;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_sub(\$12190\(48 to 63) & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(64 to 95);
                          state_var6675 <= pause_setI6445;
                        end if;
                      when q_wait6451 =>
                        \$v6452\ := \$ram_ptr_take\;
                        if \$v6452\(0) = '1' then
                          state_var6675 <= q_wait6451;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12190\(48 to 63) & X"000" & X"1")));
                          state_var6675 <= pause_getI6449;
                        end if;
                      when q_wait6455 =>
                        \$v6456\ := \$ram_ptr_take\;
                        if \$v6456\(0) = '1' then
                          state_var6675 <= q_wait6455;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$13088\(80 to 95) & X"000" & X"1")));
                          state_var6675 <= pause_getI6453;
                        end if;
                      when q_wait6460 =>
                        \$v6461\ := \$ram_ptr_take\;
                        if \$v6461\(0) = '1' then
                          state_var6675 <= q_wait6460;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(64 to 95);
                          state_var6675 <= pause_setI6458;
                        end if;
                      when q_wait6464 =>
                        \$v6465\ := \$ram_ptr_take\;
                        if \$v6465\(0) = '1' then
                          state_var6675 <= q_wait6464;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6462;
                        end if;
                      when q_wait6468 =>
                        \$v6469\ := \$ram_ptr_take\;
                        if \$v6469\(0) = '1' then
                          state_var6675 <= q_wait6468;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12190\(48 to 63) & X"000" & X"1")));
                          state_var6675 <= pause_getI6466;
                        end if;
                      when q_wait6472 =>
                        \$v6473\ := \$ram_ptr_take\;
                        if \$v6473\(0) = '1' then
                          state_var6675 <= q_wait6472;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$13134\(80 to 95) & X"000" & X"1")));
                          state_var6675 <= pause_getI6470;
                        end if;
                      when q_wait6477 =>
                        \$v6478\ := \$ram_ptr_take\;
                        if \$v6478\(0) = '1' then
                          state_var6675 <= q_wait6477;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(64 to 95);
                          state_var6675 <= pause_setI6475;
                        end if;
                      when q_wait6481 =>
                        \$v6482\ := \$ram_ptr_take\;
                        if \$v6482\(0) = '1' then
                          state_var6675 <= q_wait6481;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6479;
                        end if;
                      when q_wait6485 =>
                        \$v6486\ := \$ram_ptr_take\;
                        if \$v6486\(0) = '1' then
                          state_var6675 <= q_wait6485;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6483;
                        end if;
                      when q_wait6489 =>
                        \$v6490\ := \$ram_ptr_take\;
                        if \$v6490\(0) = '1' then
                          state_var6675 <= q_wait6489;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12190\(48 to 63) & X"000" & X"1")));
                          state_var6675 <= pause_getI6487;
                        end if;
                      when q_wait6493 =>
                        \$v6494\ := \$ram_ptr_take\;
                        if \$v6494\(0) = '1' then
                          state_var6675 <= q_wait6493;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$13192\(80 to 95) & X"000" & X"1")));
                          state_var6675 <= pause_getI6491;
                        end if;
                      when q_wait6498 =>
                        \$v6499\ := \$ram_ptr_take\;
                        if \$v6499\(0) = '1' then
                          state_var6675 <= q_wait6498;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(64 to 95);
                          state_var6675 <= pause_setI6496;
                        end if;
                      when q_wait6502 =>
                        \$v6503\ := \$ram_ptr_take\;
                        if \$v6503\(0) = '1' then
                          state_var6675 <= q_wait6502;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6500;
                        end if;
                      when q_wait6506 =>
                        \$v6507\ := \$ram_ptr_take\;
                        if \$v6507\(0) = '1' then
                          state_var6675 <= q_wait6506;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6504;
                        end if;
                      when q_wait6510 =>
                        \$v6511\ := \$ram_ptr_take\;
                        if \$v6511\(0) = '1' then
                          state_var6675 <= q_wait6510;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$12190\(48 to 63) & X"000" & X"1") & X"000" & X"1")));
                          state_var6675 <= pause_getI6508;
                        end if;
                      when q_wait6514 =>
                        \$v6515\ := \$ram_ptr_take\;
                        if \$v6515\(0) = '1' then
                          state_var6675 <= q_wait6514;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12190\(48 to 63) & X"000" & X"1")));
                          state_var6675 <= pause_getI6512;
                        end if;
                      when q_wait6518 =>
                        \$v6519\ := \$ram_ptr_take\;
                        if \$v6519\(0) = '1' then
                          state_var6675 <= q_wait6518;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6516;
                        end if;
                      when q_wait6522 =>
                        \$v6523\ := \$ram_ptr_take\;
                        if \$v6523\(0) = '1' then
                          state_var6675 <= q_wait6522;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & X"000" & X"0") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= eclat_add(\$13278_f0\(0 to 30) & \$12246_argument1\) & eclat_true;
                          state_var6675 <= pause_setI6520;
                        end if;
                      when q_wait6526 =>
                        \$v6527\ := \$ram_ptr_take\;
                        if \$v6527\(0) = '1' then
                          state_var6675 <= q_wait6526;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & X"000" & X"0") & X"000" & X"1")));
                          state_var6675 <= pause_getI6524;
                        end if;
                      when q_wait6530 =>
                        \$v6531\ := \$ram_ptr_take\;
                        if \$v6531\(0) = '1' then
                          state_var6675 <= q_wait6530;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(eclat_sub(\$12421_w594_arg\(16 to 31) & \$12421_w594_arg\(32 to 47)) & \$12421_w594_arg\(48 to 63)) & \$12421_w594_arg\(0 to 15))));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12455\;
                          state_var6675 <= pause_setI6528;
                        end if;
                      when q_wait6534 =>
                        \$v6535\ := \$ram_ptr_take\;
                        if \$v6535\(0) = '1' then
                          state_var6675 <= q_wait6534;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12421_w594_arg\(16 to 31) & \$12421_w594_arg\(0 to 15))));
                          state_var6675 <= pause_getI6532;
                        end if;
                      when q_wait6539 =>
                        \$v6540\ := \$ram_ptr_take\;
                        if \$v6540\(0) = '1' then
                          state_var6675 <= q_wait6539;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12190\(16 to 46),16) & X"000" & X"0") & X"000" & X"1")));
                          state_var6675 <= pause_getI6537;
                        end if;
                      when q_wait6543 =>
                        \$v6544\ := \$ram_ptr_take\;
                        if \$v6544\(0) = '1' then
                          state_var6675 <= q_wait6543;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12474_fill595_arg\(48 to 78),16) & \$12474_fill595_arg\(0 to 15)) & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12490_v\;
                          state_var6675 <= pause_setI6541;
                        end if;
                      when q_wait6547 =>
                        \$v6548\ := \$ram_ptr_take\;
                        if \$v6548\(0) = '1' then
                          state_var6675 <= q_wait6547;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12474_fill595_arg\(16 to 31) & X"000" & X"1")));
                          state_var6675 <= pause_getI6545;
                        end if;
                      when q_wait6552 =>
                        \$v6553\ := \$ram_ptr_take\;
                        if \$v6553\(0) = '1' then
                          state_var6675 <= q_wait6552;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12466\(64 to 94),16) & X"000" & X"0") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= eclat_resize(eclat_add(eclat_add(\$12190\(0 to 15) & X"000" & X"2") & eclat_resize(\$12248_argument2\,16)),31) & eclat_true;
                          state_var6675 <= pause_setI6550;
                        end if;
                      when q_wait6556 =>
                        \$v6557\ := \$ram_ptr_take\;
                        if \$v6557\(0) = '1' then
                          state_var6675 <= q_wait6556;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6554;
                        end if;
                      when q_wait6561 =>
                        \$v6562\ := \$ram_ptr_take\;
                        if \$v6562\(0) = '1' then
                          state_var6675 <= q_wait6561;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12524\(0 to 30),16) & eclat_resize(\$12248_argument2\,16)) & X"000" & X"1")));
                          state_var6675 <= pause_getI6559;
                        end if;
                      when q_wait6565 =>
                        \$v6566\ := \$ram_ptr_take\;
                        if \$v6566\(0) = '1' then
                          state_var6675 <= q_wait6565;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(X"3e80" & eclat_resize(\$12246_argument1\,16))));
                          state_var6675 <= pause_getI6563;
                        end if;
                      when q_wait6569 =>
                        \$v6570\ := \$ram_ptr_take\;
                        if \$v6570\(0) = '1' then
                          state_var6675 <= q_wait6569;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12540\(0 to 30),16) & eclat_resize(\$12248_argument2\,16)) & X"000" & X"1")));
                          state_var6675 <= pause_getI6567;
                        end if;
                      when q_wait6573 =>
                        \$v6574\ := \$ram_ptr_take\;
                        if \$v6574\(0) = '1' then
                          state_var6675 <= q_wait6573;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(X"3e80" & eclat_resize(\$12246_argument1\,16))));
                          state_var6675 <= pause_getI6571;
                        end if;
                      when q_wait6577 =>
                        \$v6578\ := \$ram_ptr_take\;
                        if \$v6578\(0) = '1' then
                          state_var6675 <= q_wait6577;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6575;
                        end if;
                      when q_wait6581 =>
                        \$v6582\ := \$ram_ptr_take\;
                        if \$v6582\(0) = '1' then
                          state_var6675 <= q_wait6581;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12564_fill596_arg\(48 to 78),16) & \$12564_fill596_arg\(0 to 15)) & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12580_v\;
                          state_var6675 <= pause_setI6579;
                        end if;
                      when q_wait6585 =>
                        \$v6586\ := \$ram_ptr_take\;
                        if \$v6586\(0) = '1' then
                          state_var6675 <= q_wait6585;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12564_fill596_arg\(16 to 31) & X"000" & X"1")));
                          state_var6675 <= pause_getI6583;
                        end if;
                      when q_wait6590 =>
                        \$v6591\ := \$ram_ptr_take\;
                        if \$v6591\(0) = '1' then
                          state_var6675 <= q_wait6590;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12556\(64 to 94),16) & X"000" & X"0") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12556\(0 to 31);
                          state_var6675 <= pause_setI6588;
                        end if;
                      when q_wait6594 =>
                        \$v6595\ := \$ram_ptr_take\;
                        if \$v6595\(0) = '1' then
                          state_var6675 <= q_wait6594;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12265_w0591_arg\(64 to 94),16) & eclat_sub(eclat_add(\$12265_w0591_arg\(0 to 15) & eclat_mult(X"000" & X"2" & \$12265_w0591_arg\(32 to 47))) & X"000" & X"1")) & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12376_v\;
                          state_var6675 <= pause_setI6592;
                        end if;
                      when q_wait6598 =>
                        \$v6599\ := \$ram_ptr_take\;
                        if \$v6599\(0) = '1' then
                          state_var6675 <= q_wait6598;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$12265_w0591_arg\(16 to 31) & X"000" & X"1")));
                          state_var6675 <= pause_getI6596;
                        end if;
                      when q_wait6603 =>
                        \$v6604\ := \$ram_ptr_take\;
                        if \$v6604\(0) = '1' then
                          state_var6675 <= q_wait6603;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12267_w1592_arg\(48 to 78),16) & eclat_mult(X"000" & X"2" & \$12267_w1592_arg\(0 to 15))) & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= eclat_resize(eclat_add(eclat_add(\$12267_w1592_arg\(16 to 31) & X"000" & X"2") & eclat_resize(\$12321\,16)),31) & eclat_true;
                          state_var6675 <= pause_setI6601;
                        end if;
                      when q_wait6607 =>
                        \$v6608\ := \$code_ptr_take\;
                        if \$v6608\(0) = '1' then
                          state_var6675 <= q_wait6607;
                        else
                          \$code_ptr_take\(0) := '1';
                          \$code_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(\$12267_w1592_arg\(16 to 31) & X"000" & X"3") & \$12267_w1592_arg\(0 to 15))));
                          state_var6675 <= pause_getI6605;
                        end if;
                      when q_wait6611 =>
                        \$v6612\ := \$ram_ptr_take\;
                        if \$v6612\(0) = '1' then
                          state_var6675 <= q_wait6611;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12267_w1592_arg\(48 to 78),16) & eclat_sub(eclat_mult(X"000" & X"2" & \$12267_w1592_arg\(0 to 15)) & X"000" & X"1")) & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= eclat_lor(eclat_lsl(eclat_resize("11111001",31) & "000"& X"00000" & X"18") & eclat_lsl(eclat_resize(eclat_mult(X"000" & X"2" & \$12267_w1592_arg\(0 to 15)),31) & "000"& X"000000" & X"2")) & eclat_true;
                          state_var6675 <= pause_setI6609;
                        end if;
                      when q_wait6616 =>
                        \$v6617\ := \$ram_ptr_take\;
                        if \$v6617\(0) = '1' then
                          state_var6675 <= q_wait6616;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12270_w3593_arg\(16 to 31)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= eclat_resize(eclat_add(eclat_resize(\$12270_w3593_arg\(48 to 78),16) & eclat_mult(X"000" & X"2" & \$12270_w3593_arg\(0 to 15))),31) & eclat_true;
                          state_var6675 <= pause_setI6614;
                        end if;
                      when q_wait6621 =>
                        \$v6622\ := \$ram_ptr_take\;
                        if \$v6622\(0) = '1' then
                          state_var6675 <= q_wait6621;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12266_sp\));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12257\(64 to 95);
                          state_var6675 <= pause_setI6619;
                        end if;
                      when q_wait6625 =>
                        \$v6626\ := \$ram_ptr_take\;
                        if \$v6626\(0) = '1' then
                          state_var6675 <= q_wait6625;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$12257\(64 to 94),16) & X"000" & X"0") & X"000" & X"1")));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= eclat_resize(eclat_add(eclat_add(\$12190\(0 to 15) & X"000" & X"3") & eclat_resize(\$12250_argument3\,16)),31) & eclat_true;
                          state_var6675 <= pause_setI6623;
                        end if;
                      when q_wait6629 =>
                        \$v6630\ := \$ram_ptr_take\;
                        if \$v6630\(0) = '1' then
                          state_var6675 <= q_wait6629;
                        else
                          \$ram_ptr_take\(0) := '1';
                          \$ram_ptr_write\ <= to_integer(unsigned(\$12190\(48 to 63)));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$12190\(16 to 47);
                          state_var6675 <= pause_setI6627;
                        end if;
                      when q_wait6634 =>
                        \$v6635\ := \$code_ptr_take\;
                        if \$v6635\(0) = '1' then
                          state_var6675 <= q_wait6634;
                        else
                          \$code_ptr_take\(0) := '1';
                          \$code_ptr\ <= to_integer(unsigned(\$12190\(0 to 15)));
                          state_var6675 <= pause_getI6632;
                        end if;
                      when q_wait6639 =>
                        \$v6640\ := \$code_ptr_take\;
                        if \$v6640\(0) = '1' then
                          state_var6675 <= q_wait6639;
                        else
                          \$code_ptr_take\(0) := '1';
                          \$code_ptr\ <= to_integer(unsigned(eclat_add(\$12190\(0 to 15) & X"000" & X"3")));
                          state_var6675 <= pause_getI6637;
                        end if;
                      when q_wait6644 =>
                        \$v6645\ := \$code_ptr_take\;
                        if \$v6645\(0) = '1' then
                          state_var6675 <= q_wait6644;
                        else
                          \$code_ptr_take\(0) := '1';
                          \$code_ptr\ <= to_integer(unsigned(eclat_add(\$12190\(0 to 15) & X"000" & X"2")));
                          state_var6675 <= pause_getI6642;
                        end if;
                      when q_wait6649 =>
                        \$v6650\ := \$code_ptr_take\;
                        if \$v6650\(0) = '1' then
                          state_var6675 <= q_wait6649;
                        else
                          \$code_ptr_take\(0) := '1';
                          \$code_ptr\ <= to_integer(unsigned(eclat_add(\$12190\(0 to 15) & X"000" & X"1")));
                          state_var6675 <= pause_getI6647;
                        end if;
                      when q_wait6654 =>
                        \$v6655\ := \$code_ptr_take\;
                        if \$v6655\(0) = '1' then
                          state_var6675 <= q_wait6654;
                        else
                          \$code_ptr_take\(0) := '1';
                          \$code_ptr\ <= to_integer(unsigned(\$12190\(0 to 15)));
                          state_var6675 <= pause_getI6652;
                        end if;
                      when compute5716 =>
                        rdy5715 := eclat_false;
                        eclat_print_string(of_string("pc:"));
                        
                        eclat_print_int(\$12190\(0 to 15));
                        
                        eclat_print_string(of_string("|acc:"));
                        
                        eclat_print_int(\$12190\(16 to 46));
                        
                        eclat_print_string(of_string("<"));
                        
                        \$v6657\ := ""&\$12190\(47);
                        if \$v6657\(0) = '1' then
                          eclat_print_string(of_string("int"));
                          
                          eclat_print_string(of_string(">"));
                          
                          eclat_print_string(of_string("|sp:"));
                          
                          eclat_print_int(\$12190\(48 to 63));
                          
                          eclat_print_string(of_string("|env:"));
                          
                          eclat_print_int(\$12190\(64 to 94));
                          
                          eclat_print_string(of_string("<"));
                          
                          \$v6656\ := ""&\$12190\(95);
                          if \$v6656\(0) = '1' then
                            eclat_print_string(of_string("int"));
                            
                            eclat_print_string(of_string(">"));
                            
                            eclat_print_newline(eclat_unit);
                            
                            assert eclat_lt(\$12190\(0 to 15) & std_logic_vector(to_unsigned(code'length,16))) = eclat_true report "assertion failed" severity error;
                            
                            \$v6655\ := \$code_ptr_take\;
                            if \$v6655\(0) = '1' then
                              state_var6675 <= q_wait6654;
                            else
                              \$code_ptr_take\(0) := '1';
                              \$code_ptr\ <= to_integer(unsigned(\$12190\(0 to 15)));
                              state_var6675 <= pause_getI6652;
                            end if;
                          else
                            eclat_print_string(of_string("ptr"));
                            
                            eclat_print_string(of_string(">"));
                            
                            eclat_print_newline(eclat_unit);
                            
                            assert eclat_lt(\$12190\(0 to 15) & std_logic_vector(to_unsigned(code'length,16))) = eclat_true report "assertion failed" severity error;
                            
                            \$v6655\ := \$code_ptr_take\;
                            if \$v6655\(0) = '1' then
                              state_var6675 <= q_wait6654;
                            else
                              \$code_ptr_take\(0) := '1';
                              \$code_ptr\ <= to_integer(unsigned(\$12190\(0 to 15)));
                              state_var6675 <= pause_getI6652;
                            end if;
                          end if;
                        else
                          eclat_print_string(of_string("ptr"));
                          
                          eclat_print_string(of_string(">"));
                          
                          eclat_print_string(of_string("|sp:"));
                          
                          eclat_print_int(\$12190\(48 to 63));
                          
                          eclat_print_string(of_string("|env:"));
                          
                          eclat_print_int(\$12190\(64 to 94));
                          
                          eclat_print_string(of_string("<"));
                          
                          \$v6656\ := ""&\$12190\(95);
                          if \$v6656\(0) = '1' then
                            eclat_print_string(of_string("int"));
                            
                            eclat_print_string(of_string(">"));
                            
                            eclat_print_newline(eclat_unit);
                            
                            assert eclat_lt(\$12190\(0 to 15) & std_logic_vector(to_unsigned(code'length,16))) = eclat_true report "assertion failed" severity error;
                            
                            \$v6655\ := \$code_ptr_take\;
                            if \$v6655\(0) = '1' then
                              state_var6675 <= q_wait6654;
                            else
                              \$code_ptr_take\(0) := '1';
                              \$code_ptr\ <= to_integer(unsigned(\$12190\(0 to 15)));
                              state_var6675 <= pause_getI6652;
                            end if;
                          else
                            eclat_print_string(of_string("ptr"));
                            
                            eclat_print_string(of_string(">"));
                            
                            eclat_print_newline(eclat_unit);
                            
                            assert eclat_lt(\$12190\(0 to 15) & std_logic_vector(to_unsigned(code'length,16))) = eclat_true report "assertion failed" severity error;
                            
                            \$v6655\ := \$code_ptr_take\;
                            if \$v6655\(0) = '1' then
                              state_var6675 <= q_wait6654;
                            else
                              \$code_ptr_take\(0) := '1';
                              \$code_ptr\ <= to_integer(unsigned(\$12190\(0 to 15)));
                              state_var6675 <= pause_getI6652;
                            end if;
                          end if;
                        end if;
                      end case;
                      \$v6659\ := eclat_not(rdy5715);
                      if \$v6659\(0) = '1' then
                        result5714 := \$12190\(0 to 121);
                      end if;
                      \$12196\ := result5714 & rdy5715;
                      \$12190\ := \$12196\(0 to 121) & ""&\$12196\(122);
                      rdy5712 := eclat_true;
                      state_var6674 <= compute5713;
                    end if;
                  end case;
                  \$12190\ := \$12190\;
                  \$12176\ := \$12190\;
                  \$12168\ := ""&\$12176\(120) & ""&\$12176\(122) & ""&\$12168\(2) & ""&\$12176\(121);
                  rdy5557 := eclat_true;
                  state_var6673 <= compute5558;
                end if;
              end case;
              \$12168\ := \$12168\;
              \$12143\ := \$12168\;
              \$v5556\ := ""&\$12143\(0);
              if \$v5556\(0) = '1' then
                eclat_print_string(of_string("(cy="));
                
                eclat_print_int(\$12142_cy\);
                
                eclat_print_string(of_string(")"));
                
                eclat_print_newline(eclat_unit);
                
                \$v5555\ := eclat_not(rdy5552);
                if \$v5555\(0) = '1' then
                  \$12160\ := X"0000000" & X"0";
                end if;
                case state_var6672 is
                when compute5553 =>
                  rdy5552 := eclat_false;
                  \$12160\ := eclat_if(eclat_eq(\$12160\ & eclat_add(X"00" & X"989680" & X"00" & X"989680")) & X"0000000" & X"0" & eclat_add(\$12160\ & X"0000000" & X"1"));
                  rdy5552 := eclat_true;
                  state_var6672 <= compute5553;
                end case;
                \$12160\ := \$12160\;
                \$12149\ := \$12160\;
                result5549 := ""&\$12143\(0) & eclat_not(""&\$12143\(1)) & eclat_gt(\$12149\ & X"00" & X"989680") & ""&\$12143\(3) & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & "00000011" & "00000011" & "00000011" & "00000011" & "00000011" & "00000011";
                rdy5550 := eclat_true;
                state <= compute5551;
              else
                \$v5555\ := eclat_not(rdy5552);
                if \$v5555\(0) = '1' then
                  \$12160\ := X"0000000" & X"0";
                end if;
                case state_var6672 is
                when compute5553 =>
                  rdy5552 := eclat_false;
                  \$12160\ := eclat_if(eclat_eq(\$12160\ & eclat_add(X"00" & X"989680" & X"00" & X"989680")) & X"0000000" & X"0" & eclat_add(\$12160\ & X"0000000" & X"1"));
                  rdy5552 := eclat_true;
                  state_var6672 <= compute5553;
                end case;
                \$12160\ := \$12160\;
                \$12149\ := \$12160\;
                result5549 := ""&\$12143\(0) & eclat_not(""&\$12143\(1)) & eclat_gt(\$12149\ & X"00" & X"989680") & ""&\$12143\(3) & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & "00000011" & "00000011" & "00000011" & "00000011" & "00000011" & "00000011";
                rdy5550 := eclat_true;
                state <= compute5551;
              end if;
            end if;
          end case;
          
          result <= result5549;
          rdy <= rdy5550;
          
        end if;
      end if;
    end if;
  end process;
end architecture;
